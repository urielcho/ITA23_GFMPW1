magic
tech gf180mcuD
magscale 1 10
timestamp 1699711871
<< metal1 >>
rect 40226 71150 40238 71202
rect 40290 71199 40302 71202
rect 43810 71199 43822 71202
rect 40290 71153 43822 71199
rect 40290 71150 40302 71153
rect 43810 71150 43822 71153
rect 43874 71150 43886 71202
rect 371186 70590 371198 70642
rect 371250 70639 371262 70642
rect 373538 70639 373550 70642
rect 371250 70593 373550 70639
rect 371250 70590 371262 70593
rect 373538 70590 373550 70593
rect 373602 70590 373614 70642
<< via1 >>
rect 40238 71150 40290 71202
rect 43822 71150 43874 71202
rect 371198 70590 371250 70642
rect 373550 70590 373602 70642
<< metal2 >>
rect 11032 595672 11256 597000
rect 11004 595560 11256 595672
rect 33096 595672 33320 597000
rect 33096 595560 33348 595672
rect 55160 595560 55384 597000
rect 77224 595560 77448 597000
rect 99288 595672 99512 597000
rect 99288 595560 99540 595672
rect 121352 595560 121576 597000
rect 143416 595672 143640 597000
rect 143388 595560 143640 595672
rect 165480 595672 165704 597000
rect 165480 595560 165732 595672
rect 187544 595560 187768 597000
rect 209608 595672 209832 597000
rect 231672 595672 231896 597000
rect 209580 595560 209832 595672
rect 231644 595560 231896 595672
rect 253736 595560 253960 597000
rect 275800 595672 276024 597000
rect 297864 595672 298088 597000
rect 275772 595560 276024 595672
rect 297836 595560 298088 595672
rect 319928 595560 320152 597000
rect 341992 595672 342216 597000
rect 364056 595672 364280 597000
rect 341964 595560 342216 595672
rect 364028 595560 364280 595672
rect 386120 595560 386344 597000
rect 408184 595560 408408 597000
rect 430248 595672 430472 597000
rect 430220 595560 430472 595672
rect 452312 595560 452536 597000
rect 474376 595672 474600 597000
rect 496440 595672 496664 597000
rect 474348 595560 474600 595672
rect 496412 595560 496664 595672
rect 518504 595560 518728 597000
rect 540568 595672 540792 597000
rect 562632 595672 562856 597000
rect 540540 595560 540792 595672
rect 562604 595560 562856 595672
rect 584696 595560 584920 597000
rect 11004 578788 11060 595560
rect 33292 590548 33348 595560
rect 33292 590482 33348 590492
rect 46172 590548 46228 590558
rect 46172 583828 46228 590492
rect 46172 583762 46228 583772
rect 11004 578722 11060 578732
rect 77308 573748 77364 595560
rect 99484 590548 99540 595560
rect 99484 590482 99540 590492
rect 143388 573972 143444 595560
rect 165676 590660 165732 595560
rect 165676 590594 165732 590604
rect 209580 582260 209636 595560
rect 209580 582194 209636 582204
rect 231644 577220 231700 595560
rect 231644 577154 231700 577164
rect 275772 574084 275828 595560
rect 284732 590660 284788 590670
rect 279244 582148 279300 582158
rect 275772 574018 275828 574028
rect 278124 575428 278180 575438
rect 143388 573906 143444 573916
rect 77308 573682 77364 573692
rect 76412 573076 76468 573086
rect 40236 571956 40292 571966
rect 38892 571396 38948 571406
rect 4284 570724 4340 570734
rect 4172 567252 4228 567262
rect 4172 559188 4228 567196
rect 4172 559122 4228 559132
rect 4172 523348 4228 523358
rect 4172 51156 4228 523292
rect 4284 220500 4340 570668
rect 36876 569604 36932 569614
rect 36876 569492 36932 569548
rect 36232 569436 36932 569492
rect 38892 569464 38948 571340
rect 40236 570724 40292 571900
rect 44268 571732 44324 571742
rect 41580 571508 41636 571518
rect 40236 570668 40404 570724
rect 40236 570500 40292 570510
rect 40012 570444 40236 570500
rect 40012 569492 40068 570444
rect 40236 570434 40292 570444
rect 40348 570276 40404 570668
rect 39592 569436 40068 569492
rect 40236 570220 40404 570276
rect 40236 569464 40292 570220
rect 41580 569464 41636 571452
rect 44268 569464 44324 571676
rect 62972 571732 63028 571742
rect 45612 571620 45668 571630
rect 45612 569464 45668 571564
rect 46956 571284 47012 571294
rect 46732 569716 46788 569726
rect 46732 569492 46788 569660
rect 46312 569436 46788 569492
rect 46956 569464 47012 571228
rect 4508 569380 4564 569390
rect 4396 567140 4452 567150
rect 4396 262836 4452 567084
rect 4508 474516 4564 569324
rect 15932 569156 15988 569166
rect 4508 474450 4564 474460
rect 7644 569044 7700 569054
rect 7532 403732 7588 403742
rect 4396 262770 4452 262780
rect 4508 296548 4564 296558
rect 4284 220434 4340 220444
rect 4396 234500 4452 234510
rect 4396 178052 4452 234444
rect 4396 177986 4452 177996
rect 4396 149716 4452 149726
rect 4172 51090 4228 51100
rect 4284 107380 4340 107390
rect 4284 31108 4340 107324
rect 4396 91588 4452 149660
rect 4508 135828 4564 296492
rect 4620 192052 4676 192062
rect 4620 150388 4676 191996
rect 4620 150322 4676 150332
rect 4508 135762 4564 135772
rect 4396 91522 4452 91532
rect 4396 65044 4452 65054
rect 4396 52948 4452 64988
rect 4396 52882 4452 52892
rect 4284 31042 4340 31052
rect 7532 29428 7588 403676
rect 7644 347508 7700 568988
rect 7644 347442 7700 347452
rect 12572 530740 12628 530750
rect 7532 29362 7588 29372
rect 10892 52948 10948 52958
rect 10892 26180 10948 52892
rect 12572 29652 12628 530684
rect 12572 29586 12628 29596
rect 14252 488404 14308 488414
rect 14252 29540 14308 488348
rect 15932 389620 15988 569100
rect 18396 554484 18452 554494
rect 18396 484036 18452 554428
rect 36204 525028 36260 527688
rect 36204 524962 36260 524972
rect 38220 511588 38276 527688
rect 38220 511522 38276 511532
rect 39564 503076 39620 527688
rect 40236 523460 40292 527688
rect 40236 523394 40292 523404
rect 40908 518532 40964 527688
rect 40908 518466 40964 518476
rect 62972 506548 63028 571676
rect 69692 571620 69748 571630
rect 63196 571284 63252 571294
rect 63196 528164 63252 571228
rect 63196 528098 63252 528108
rect 62972 506482 63028 506492
rect 69692 505876 69748 571564
rect 73052 571508 73108 571518
rect 73052 506660 73108 571452
rect 73052 506594 73108 506604
rect 69692 505810 69748 505820
rect 39564 503010 39620 503020
rect 36204 500948 36260 500958
rect 36204 498344 36260 500892
rect 62972 500948 63028 500958
rect 40908 500836 40964 500846
rect 36876 500724 36932 500734
rect 36876 498344 36932 500668
rect 37548 499044 37604 499054
rect 37548 498344 37604 498988
rect 40908 498344 40964 500780
rect 46956 499268 47012 499278
rect 46956 498344 47012 499212
rect 43596 497812 43652 497822
rect 43596 497746 43652 497756
rect 18396 483970 18452 483980
rect 38220 439348 38276 456456
rect 40236 452788 40292 456456
rect 40236 452722 40292 452732
rect 38220 439282 38276 439292
rect 42924 437780 42980 456456
rect 44940 439460 44996 456456
rect 62972 445396 63028 500892
rect 62972 445330 63028 445340
rect 74732 500836 74788 500846
rect 44940 439394 44996 439404
rect 74732 437892 74788 500780
rect 74732 437826 74788 437836
rect 42924 437714 42980 437724
rect 38892 430724 38948 430734
rect 38556 427588 38612 427598
rect 38556 427140 38612 427532
rect 38248 427084 38612 427140
rect 38892 427112 38948 430668
rect 39564 430276 39620 430286
rect 39564 427112 39620 430220
rect 69692 430276 69748 430286
rect 42924 428484 42980 428494
rect 42924 427112 42980 428428
rect 40236 426804 40292 426814
rect 40236 426738 40292 426748
rect 44268 426580 44324 426590
rect 44268 426514 44324 426524
rect 15932 389554 15988 389564
rect 18396 411796 18452 411806
rect 18396 409444 18452 411740
rect 18396 341684 18452 409388
rect 69692 385924 69748 430220
rect 69692 385858 69748 385868
rect 73052 426580 73108 426590
rect 42252 380660 42308 385336
rect 42252 380594 42308 380604
rect 42924 380548 42980 385336
rect 42924 380482 42980 380492
rect 73052 360836 73108 426524
rect 73052 360770 73108 360780
rect 45612 358260 45668 358270
rect 36204 358148 36260 358158
rect 35532 358036 35588 358046
rect 35532 355880 35588 357980
rect 36204 355880 36260 358092
rect 38892 357924 38948 357934
rect 38892 355880 38948 357868
rect 40908 356356 40964 356366
rect 40908 355880 40964 356300
rect 44268 356244 44324 356254
rect 44268 355880 44324 356188
rect 45612 355880 45668 358204
rect 62188 358260 62244 358270
rect 61292 358148 61348 358158
rect 34860 355572 34916 355582
rect 34860 355506 34916 355516
rect 40236 355348 40292 355358
rect 40236 355282 40292 355292
rect 61292 353668 61348 358092
rect 62188 353780 62244 358204
rect 62188 353714 62244 353724
rect 62972 358036 63028 358046
rect 61292 353602 61348 353612
rect 14252 29474 14308 29484
rect 15932 319060 15988 319070
rect 15932 28532 15988 319004
rect 18396 270452 18452 341628
rect 44268 314132 44324 314142
rect 36876 300916 36932 314104
rect 38892 305396 38948 314104
rect 38892 305330 38948 305340
rect 43596 302596 43652 314104
rect 55720 314076 56420 314132
rect 44268 314066 44324 314076
rect 56364 314020 56420 314076
rect 56364 313954 56420 313964
rect 43596 302530 43652 302540
rect 62972 301476 63028 357980
rect 62972 301410 63028 301420
rect 74732 357924 74788 357934
rect 36876 300850 36932 300860
rect 74732 300356 74788 357868
rect 74732 300290 74788 300300
rect 45052 288260 45108 288270
rect 40236 287476 40292 287486
rect 40236 284788 40292 287420
rect 41916 285796 41972 285806
rect 41356 285684 41412 285694
rect 41356 284788 41412 285628
rect 41916 284788 41972 285740
rect 45052 284788 45108 288204
rect 39592 284732 40292 284788
rect 40936 284732 41412 284788
rect 41608 284732 41972 284788
rect 44296 284732 45108 284788
rect 37548 284340 37604 284350
rect 37548 284274 37604 284284
rect 42252 284228 42308 284238
rect 42252 284162 42308 284172
rect 18396 198996 18452 270396
rect 18396 197876 18452 198940
rect 18396 127988 18452 197820
rect 18396 56868 18452 127932
rect 18396 56802 18452 56812
rect 19292 276724 19348 276734
rect 19292 29092 19348 276668
rect 26796 240212 26852 242872
rect 26796 240146 26852 240156
rect 37548 240100 37604 242872
rect 38220 241780 38276 242872
rect 38220 241714 38276 241724
rect 37548 240034 37604 240044
rect 40236 239540 40292 242872
rect 42924 239876 42980 242872
rect 44268 241892 44324 242872
rect 44268 241826 44324 241836
rect 46284 239988 46340 242872
rect 48636 241108 48692 241118
rect 48636 240212 48692 241052
rect 48636 240146 48692 240156
rect 46284 239922 46340 239932
rect 42924 239810 42980 239820
rect 40236 239474 40292 239484
rect 41580 216020 41636 216030
rect 40908 215460 40964 215470
rect 35532 215348 35588 215358
rect 35532 213528 35588 215292
rect 40908 213528 40964 215404
rect 41580 213528 41636 215964
rect 61292 215460 61348 215470
rect 44940 215124 44996 215134
rect 44940 213528 44996 215068
rect 46956 213668 47012 213678
rect 45612 213556 45668 213566
rect 46956 213556 47012 213612
rect 46312 213500 47012 213556
rect 45612 213490 45668 213500
rect 40236 213444 40292 213454
rect 40236 213378 40292 213388
rect 44268 212996 44324 213006
rect 44268 212930 44324 212940
rect 61292 210868 61348 215404
rect 61292 210802 61348 210812
rect 69692 213108 69748 213118
rect 62076 173908 62132 173918
rect 34888 171612 35252 171668
rect 38248 171612 38612 171668
rect 38920 171612 39620 171668
rect 40936 171612 41636 171668
rect 35196 169540 35252 171612
rect 35196 169474 35252 169484
rect 38556 168980 38612 171612
rect 39564 169428 39620 171612
rect 41580 171220 41636 171612
rect 41580 171154 41636 171164
rect 43484 171612 43624 171668
rect 44296 171612 44996 171668
rect 39564 169362 39620 169372
rect 43484 169316 43540 171612
rect 44940 171332 44996 171612
rect 44940 171266 44996 171276
rect 43484 169250 43540 169260
rect 62076 169316 62132 173852
rect 69692 171220 69748 213052
rect 69692 171154 69748 171164
rect 62076 169250 62132 169260
rect 38556 168914 38612 168924
rect 69692 155876 69748 155886
rect 42252 152516 42308 152526
rect 38220 145012 38276 145022
rect 38220 142296 38276 144956
rect 40908 142884 40964 142894
rect 40908 142296 40964 142828
rect 42252 142296 42308 152460
rect 62972 151956 63028 151966
rect 42924 144676 42980 144686
rect 42924 142296 42980 144620
rect 43596 101108 43652 101118
rect 43596 101042 43652 101052
rect 45612 101108 45668 101118
rect 45612 101042 45668 101052
rect 44268 100996 44324 101006
rect 44268 100930 44324 100940
rect 37548 100884 37604 100894
rect 37548 100818 37604 100828
rect 38220 98980 38276 100520
rect 38220 98914 38276 98924
rect 38892 98868 38948 100520
rect 42252 99092 42308 100520
rect 42252 99026 42308 99036
rect 38892 98802 38948 98812
rect 62972 98868 63028 151900
rect 69692 100884 69748 155820
rect 74732 155316 74788 155326
rect 69692 100818 69748 100828
rect 73052 152068 73108 152078
rect 73052 98980 73108 152012
rect 74732 101668 74788 155260
rect 74732 101602 74788 101612
rect 73052 98914 73108 98924
rect 62972 98802 63028 98812
rect 74732 95956 74788 95966
rect 62972 94836 63028 94846
rect 42252 90020 42308 90030
rect 41580 84980 41636 84990
rect 38892 79828 38948 79838
rect 35532 74228 35588 74238
rect 35532 71064 35588 74172
rect 38892 71064 38948 79772
rect 40236 71202 40292 71214
rect 40236 71150 40238 71202
rect 40290 71150 40292 71202
rect 40236 71092 40292 71150
rect 39592 71036 40292 71092
rect 41580 71064 41636 84924
rect 42252 71064 42308 89964
rect 50316 88228 50372 88238
rect 45612 74116 45668 74126
rect 45276 72436 45332 72446
rect 43820 71202 43876 71214
rect 43820 71150 43822 71202
rect 43874 71150 43876 71202
rect 43820 70532 43876 71150
rect 45276 71092 45332 72380
rect 44968 71036 45332 71092
rect 45612 71064 45668 74060
rect 50316 71064 50372 88172
rect 43820 70466 43876 70476
rect 61292 31220 61348 31230
rect 19292 29026 19348 29036
rect 15932 28466 15988 28476
rect 38892 26516 38948 29288
rect 39564 26628 39620 29288
rect 39564 26562 39620 26572
rect 38892 26450 38948 26460
rect 40236 26404 40292 29288
rect 42924 26740 42980 29288
rect 43596 28420 43652 29288
rect 43596 28354 43652 28364
rect 55692 26852 55748 29288
rect 55692 26786 55748 26796
rect 42924 26674 42980 26684
rect 40236 26338 40292 26348
rect 61292 26404 61348 31164
rect 62972 26516 63028 94780
rect 73052 93380 73108 93390
rect 63084 71316 63140 71326
rect 63084 28420 63140 71260
rect 63084 28354 63140 28364
rect 73052 26628 73108 93324
rect 74732 26852 74788 95900
rect 76412 29764 76468 573020
rect 266252 572404 266308 572414
rect 249452 572180 249508 572190
rect 160188 571844 160244 571854
rect 104860 571620 104916 571630
rect 100156 571508 100212 571518
rect 78092 571396 78148 571406
rect 78092 503188 78148 571340
rect 100156 569464 100212 571452
rect 104860 569464 104916 571564
rect 130172 571620 130228 571630
rect 107548 571396 107604 571406
rect 107548 569464 107604 571340
rect 125132 569716 125188 569726
rect 98812 525140 98868 527688
rect 98812 525074 98868 525084
rect 99484 512036 99540 527688
rect 100156 523572 100212 527688
rect 100156 523506 100212 523516
rect 99484 511970 99540 511980
rect 102172 510020 102228 527688
rect 102844 511476 102900 527688
rect 103516 516740 103572 527688
rect 106876 522004 106932 527688
rect 106876 521938 106932 521948
rect 107548 521892 107604 527688
rect 107548 521826 107604 521836
rect 103516 516674 103572 516684
rect 102844 511410 102900 511420
rect 102172 509954 102228 509964
rect 125132 503636 125188 569660
rect 130172 513268 130228 571564
rect 130172 513202 130228 513212
rect 136892 571508 136948 571518
rect 125132 503570 125188 503580
rect 78092 503122 78148 503132
rect 98812 501172 98868 501182
rect 98812 498344 98868 501116
rect 125132 501172 125188 501182
rect 100156 501060 100212 501070
rect 100156 498344 100212 501004
rect 100828 500948 100884 500958
rect 100828 498344 100884 500892
rect 104860 500836 104916 500846
rect 104188 499156 104244 499166
rect 103516 498372 103572 498382
rect 104188 498344 104244 499100
rect 104860 498344 104916 500780
rect 103516 498306 103572 498316
rect 125132 456596 125188 501116
rect 125132 456530 125188 456540
rect 130172 501060 130228 501070
rect 76412 29698 76468 29708
rect 78092 446068 78148 446078
rect 78092 28420 78148 446012
rect 100828 444388 100884 456456
rect 102844 447748 102900 456456
rect 103516 453236 103572 456456
rect 103516 453170 103572 453180
rect 104188 452116 104244 456456
rect 104188 452050 104244 452060
rect 102844 447682 102900 447692
rect 100828 444322 100884 444332
rect 130172 439684 130228 501004
rect 135212 500948 135268 500958
rect 135212 441252 135268 500892
rect 136892 496468 136948 571452
rect 160188 569464 160244 571788
rect 187292 571844 187348 571854
rect 170268 571732 170324 571742
rect 164220 571620 164276 571630
rect 160860 571508 160916 571518
rect 160860 569464 160916 571452
rect 162876 569940 162932 569950
rect 162876 569464 162932 569884
rect 164220 569464 164276 571564
rect 169596 570052 169652 570062
rect 168924 569828 168980 569838
rect 166460 569716 166516 569726
rect 166460 569492 166516 569660
rect 166264 569436 166516 569492
rect 168924 569464 168980 569772
rect 169596 569464 169652 569996
rect 170268 569464 170324 571676
rect 157052 518532 157108 518542
rect 157052 501396 157108 518476
rect 160188 513380 160244 527688
rect 162876 523796 162932 527688
rect 164220 525252 164276 527688
rect 164220 525186 164276 525196
rect 162876 523730 162932 523740
rect 160188 513314 160244 513324
rect 167580 508228 167636 527688
rect 168252 518756 168308 527688
rect 168924 523684 168980 527688
rect 168924 523618 168980 523628
rect 168252 518690 168308 518700
rect 167580 508162 167636 508172
rect 169596 504980 169652 527688
rect 170492 523572 170548 523582
rect 170492 510356 170548 523516
rect 170492 510290 170548 510300
rect 169596 504914 169652 504924
rect 157052 501330 157108 501340
rect 166236 501060 166292 501070
rect 164220 499492 164276 499502
rect 155484 499380 155540 499390
rect 155484 498344 155540 499324
rect 162876 498484 162932 498494
rect 162876 498372 162932 498428
rect 162232 498316 162932 498372
rect 164220 498344 164276 499436
rect 166236 498344 166292 501004
rect 170940 500948 170996 500958
rect 170940 498344 170996 500892
rect 166908 498260 166964 498270
rect 166908 498194 166964 498204
rect 187292 498148 187348 571788
rect 224812 571844 224868 571854
rect 224140 571284 224196 571294
rect 187404 570052 187460 570062
rect 187404 518196 187460 569996
rect 192332 569940 192388 569950
rect 187404 518130 187460 518140
rect 188076 522004 188132 522014
rect 188076 515396 188132 521948
rect 192332 519316 192388 569884
rect 199052 569828 199108 569838
rect 198156 523684 198212 523694
rect 192332 519250 192388 519260
rect 192444 521892 192500 521902
rect 188076 515330 188132 515340
rect 192444 509796 192500 521836
rect 198156 517076 198212 523628
rect 199052 517636 199108 569772
rect 224140 569464 224196 571228
rect 224812 569464 224868 571788
rect 247996 571732 248052 571742
rect 247772 571620 247828 571630
rect 231532 570052 231588 570062
rect 228172 569940 228228 569950
rect 226156 569828 226212 569838
rect 226156 569464 226212 569772
rect 228172 569464 228228 569884
rect 231532 569464 231588 569996
rect 230860 568932 230916 568942
rect 230860 568866 230916 568876
rect 227500 527940 227556 527950
rect 226856 527884 227500 527940
rect 227500 527874 227556 527884
rect 224028 527828 224084 527838
rect 223496 527772 224028 527828
rect 224028 527762 224084 527772
rect 224812 527716 224868 527726
rect 224168 527660 224756 527716
rect 224700 526036 224756 527660
rect 224812 527650 224868 527660
rect 224700 525970 224756 525980
rect 230188 525364 230244 527688
rect 230188 525298 230244 525308
rect 244412 525364 244468 525374
rect 199052 517570 199108 517580
rect 198156 517010 198212 517020
rect 192444 509730 192500 509740
rect 187292 498082 187348 498092
rect 187404 501060 187460 501070
rect 164892 498036 164948 498046
rect 164892 497970 164948 497980
rect 179004 497924 179060 497934
rect 179004 497858 179060 497868
rect 136892 496402 136948 496412
rect 160860 456932 160916 456942
rect 160860 456866 160916 456876
rect 162876 449540 162932 456456
rect 162876 449474 162932 449484
rect 166236 442708 166292 456456
rect 166236 442642 166292 442652
rect 135212 441186 135268 441196
rect 130172 439618 130228 439628
rect 166908 434196 166964 456456
rect 168924 435316 168980 456456
rect 168924 435250 168980 435260
rect 170492 449540 170548 449550
rect 166908 434130 166964 434140
rect 170492 432516 170548 449484
rect 170492 432450 170548 432460
rect 171388 430724 171444 430734
rect 162876 430612 162932 430622
rect 105532 430500 105588 430510
rect 103516 430388 103572 430398
rect 98140 430276 98196 430286
rect 98140 427112 98196 430220
rect 102844 428596 102900 428606
rect 102844 427112 102900 428540
rect 103516 427112 103572 430332
rect 105532 427112 105588 430444
rect 130172 430500 130228 430510
rect 99484 427028 99540 427038
rect 99484 426962 99540 426972
rect 102172 426916 102228 426926
rect 102172 426850 102228 426860
rect 88060 426468 88116 426478
rect 88060 426402 88116 426412
rect 100156 365876 100212 385336
rect 100828 367556 100884 385336
rect 103516 368676 103572 385336
rect 105532 384692 105588 385336
rect 105532 384626 105588 384636
rect 106204 384580 106260 385336
rect 106204 384514 106260 384524
rect 103516 368610 103572 368620
rect 100828 367490 100884 367500
rect 107548 366996 107604 385336
rect 130172 373828 130228 430444
rect 161532 430164 161588 430174
rect 161532 427112 161588 430108
rect 162876 427112 162932 430556
rect 168924 430500 168980 430510
rect 165564 428820 165620 428830
rect 164220 428708 164276 428718
rect 164220 427112 164276 428652
rect 165564 427112 165620 428764
rect 167580 427140 167636 427150
rect 168924 427112 168980 430444
rect 171388 427700 171444 430668
rect 187292 430612 187348 430622
rect 171388 427634 171444 427644
rect 174636 430388 174692 430398
rect 167580 427074 167636 427084
rect 166236 426692 166292 426702
rect 166236 426626 166292 426636
rect 174636 426692 174692 430332
rect 174636 426626 174692 426636
rect 160860 426468 160916 426478
rect 160860 426402 160916 426412
rect 170268 426468 170324 426478
rect 170268 426402 170324 426412
rect 168252 385364 168308 385374
rect 167580 376516 167636 385336
rect 168252 385298 168308 385308
rect 167580 376450 167636 376460
rect 130172 373762 130228 373772
rect 187292 370916 187348 430556
rect 187404 429716 187460 501004
rect 195692 500948 195748 500958
rect 187516 498260 187572 498270
rect 187516 431396 187572 498204
rect 187516 431330 187572 431340
rect 192332 498036 192388 498046
rect 192332 430836 192388 497980
rect 195692 447860 195748 500892
rect 230188 500948 230244 500958
rect 200732 500836 200788 500846
rect 197372 499268 197428 499278
rect 197372 449876 197428 499212
rect 197372 449810 197428 449820
rect 199052 497812 199108 497822
rect 195692 447794 195748 447804
rect 199052 447076 199108 497756
rect 199052 447010 199108 447020
rect 192332 430770 192388 430780
rect 197372 430500 197428 430510
rect 187404 429650 187460 429660
rect 195692 430164 195748 430174
rect 192332 428820 192388 428830
rect 188972 427140 189028 427150
rect 187404 426020 187460 426030
rect 187404 373156 187460 425964
rect 188972 373716 189028 427084
rect 189084 426132 189140 426142
rect 189084 375956 189140 426076
rect 189084 375890 189140 375900
rect 192332 374836 192388 428764
rect 192332 374770 192388 374780
rect 188972 373650 189028 373660
rect 187404 373090 187460 373100
rect 195692 372596 195748 430108
rect 197372 375396 197428 430444
rect 200732 424676 200788 500780
rect 226156 500836 226212 500846
rect 222796 499604 222852 499614
rect 205772 499044 205828 499054
rect 205772 443716 205828 498988
rect 222796 498344 222852 499548
rect 226156 498344 226212 500780
rect 230188 498344 230244 500892
rect 231532 499268 231588 499278
rect 231532 498344 231588 499212
rect 232204 499044 232260 499054
rect 232204 498344 232260 498988
rect 244412 498596 244468 525308
rect 244412 498530 244468 498540
rect 226828 497812 226884 497822
rect 226828 497746 226884 497756
rect 247772 489076 247828 571564
rect 247996 489636 248052 571676
rect 249452 523348 249508 572124
rect 257852 571956 257908 571966
rect 256172 571844 256228 571854
rect 249676 571284 249732 571294
rect 249676 525476 249732 571228
rect 249676 525410 249732 525420
rect 252812 569604 252868 569614
rect 249900 525028 249956 525038
rect 249452 523282 249508 523292
rect 249676 523460 249732 523470
rect 249564 513380 249620 513390
rect 247996 489570 248052 489580
rect 249452 498484 249508 498494
rect 247772 489010 247828 489020
rect 248108 472836 248164 472846
rect 247772 470596 247828 470606
rect 230860 456932 230916 456942
rect 230860 456866 230916 456876
rect 229516 456708 229572 456718
rect 229516 456642 229572 456652
rect 227500 456484 227556 456494
rect 222124 450324 222180 456456
rect 222796 453572 222852 456456
rect 226156 455252 226212 456456
rect 227500 456418 227556 456428
rect 226156 455186 226212 455196
rect 231532 455140 231588 456456
rect 231532 455074 231588 455084
rect 247772 455140 247828 470540
rect 248108 456708 248164 472780
rect 249452 464436 249508 498428
rect 249564 493556 249620 513324
rect 249564 493490 249620 493500
rect 249676 476756 249732 523404
rect 249900 479668 249956 524972
rect 249900 479602 249956 479612
rect 249676 476690 249732 476700
rect 252812 476196 252868 569548
rect 254492 568932 254548 568942
rect 253036 525252 253092 525262
rect 252812 476130 252868 476140
rect 252924 499604 252980 499614
rect 249452 464370 249508 464380
rect 249564 467236 249620 467246
rect 248108 456642 248164 456652
rect 249564 455252 249620 467180
rect 252028 465556 252084 465566
rect 252028 458052 252084 465500
rect 252028 457986 252084 457996
rect 249564 455186 249620 455196
rect 247772 455074 247828 455084
rect 222796 453506 222852 453516
rect 247772 452788 247828 452798
rect 222124 450258 222180 450268
rect 225932 450324 225988 450334
rect 205772 443650 205828 443660
rect 202412 442708 202468 442718
rect 202412 432068 202468 442652
rect 225932 438676 225988 450268
rect 225932 438610 225988 438620
rect 202412 432002 202468 432012
rect 230860 430612 230916 430622
rect 222124 430500 222180 430510
rect 211372 427140 211428 427150
rect 222124 427112 222180 430444
rect 226828 430388 226884 430398
rect 223356 430276 223412 430286
rect 223356 429268 223412 430220
rect 223356 429202 223412 429212
rect 224140 430164 224196 430174
rect 224140 427112 224196 430108
rect 226828 427112 226884 430332
rect 228172 430276 228228 430286
rect 228172 427112 228228 430220
rect 229628 427252 229684 427262
rect 229628 427140 229684 427196
rect 228872 427084 229684 427140
rect 230860 427112 230916 430556
rect 240268 428820 240324 428830
rect 240268 427112 240324 428764
rect 211372 427074 211428 427084
rect 222796 426468 222852 426478
rect 222796 426402 222852 426412
rect 232204 426468 232260 426478
rect 232204 426402 232260 426412
rect 200732 424610 200788 424620
rect 247772 421316 247828 452732
rect 249564 447748 249620 447758
rect 249452 428596 249508 428606
rect 247772 421250 247828 421260
rect 247884 427252 247940 427262
rect 247884 414596 247940 427196
rect 247884 414530 247940 414540
rect 247772 401156 247828 401166
rect 230860 385588 230916 385598
rect 230860 385522 230916 385532
rect 247772 385364 247828 401100
rect 249452 394436 249508 428540
rect 249564 422996 249620 447692
rect 252924 440356 252980 499548
rect 253036 491876 253092 525196
rect 253036 491810 253092 491820
rect 253148 499044 253204 499054
rect 253148 466676 253204 498988
rect 254492 495796 254548 568876
rect 254492 495730 254548 495740
rect 254604 510020 254660 510030
rect 254604 482916 254660 509964
rect 254716 504980 254772 504990
rect 254716 490196 254772 504924
rect 256172 494676 256228 571788
rect 256172 494610 256228 494620
rect 256284 497924 256340 497934
rect 254716 490130 254772 490140
rect 254604 482850 254660 482860
rect 253148 466610 253204 466620
rect 256172 471156 256228 471166
rect 256172 458164 256228 471100
rect 256284 461076 256340 497868
rect 257852 480452 257908 571900
rect 263004 571508 263060 571518
rect 261212 571396 261268 571406
rect 259756 570052 259812 570062
rect 257964 569940 258020 569950
rect 257964 494116 258020 569884
rect 259532 569716 259588 569726
rect 258188 525140 258244 525150
rect 257964 494050 258020 494060
rect 258076 498372 258132 498382
rect 257852 480386 257908 480396
rect 256284 461010 256340 461020
rect 257852 468692 257908 468702
rect 256172 458098 256228 458108
rect 257852 453572 257908 468636
rect 258076 454916 258132 498316
rect 258188 481236 258244 525084
rect 258188 481170 258244 481180
rect 258300 499268 258356 499278
rect 258300 468356 258356 499212
rect 259532 491316 259588 569660
rect 259756 527156 259812 569996
rect 259756 527090 259812 527100
rect 259756 516740 259812 516750
rect 259532 491250 259588 491260
rect 259644 499156 259700 499166
rect 258300 468290 258356 468300
rect 259532 468916 259588 468926
rect 259532 456484 259588 468860
rect 259532 456418 259588 456428
rect 258076 454850 258132 454860
rect 257852 453506 257908 453516
rect 252924 440290 252980 440300
rect 258076 444388 258132 444398
rect 253036 439348 253092 439358
rect 249788 430500 249844 430510
rect 249564 422930 249620 422940
rect 249676 426244 249732 426254
rect 249676 402276 249732 426188
rect 249788 409556 249844 430444
rect 252924 428708 252980 428718
rect 249788 409490 249844 409500
rect 252812 427028 252868 427038
rect 249676 402210 249732 402220
rect 252812 396116 252868 426972
rect 252924 405636 252980 428652
rect 253036 421876 253092 439292
rect 257852 430612 257908 430622
rect 256172 428484 256228 428494
rect 253036 421810 253092 421820
rect 253148 426020 253204 426030
rect 253148 412356 253204 425964
rect 253148 412290 253204 412300
rect 252924 405570 252980 405580
rect 252812 396050 252868 396060
rect 249452 394370 249508 394380
rect 222796 384468 222852 385336
rect 222796 384402 222852 384412
rect 229516 377636 229572 385336
rect 247772 385298 247828 385308
rect 249676 393876 249732 393886
rect 249676 384580 249732 393820
rect 256172 391636 256228 428428
rect 256284 427140 256340 427150
rect 256284 408436 256340 427084
rect 256284 408370 256340 408380
rect 256172 391570 256228 391580
rect 256284 393316 256340 393326
rect 256284 384692 256340 393260
rect 256284 384626 256340 384636
rect 249676 384514 249732 384524
rect 257852 383124 257908 430556
rect 257964 426356 258020 426366
rect 257964 392196 258020 426300
rect 258076 422436 258132 444332
rect 258300 439460 258356 439470
rect 258076 422370 258132 422380
rect 258188 426916 258244 426926
rect 257964 392130 258020 392140
rect 258076 411796 258132 411806
rect 258076 384468 258132 411740
rect 258188 399476 258244 426860
rect 258300 417396 258356 439404
rect 258300 417330 258356 417340
rect 259532 430388 259588 430398
rect 258188 399410 258244 399420
rect 258076 384402 258132 384412
rect 257852 383058 257908 383068
rect 229516 377570 229572 377580
rect 247772 380660 247828 380670
rect 197372 375330 197428 375340
rect 195692 372530 195748 372540
rect 187292 370850 187348 370860
rect 107548 366930 107604 366940
rect 100156 365810 100212 365820
rect 247772 359156 247828 380604
rect 259532 379316 259588 430332
rect 259644 427476 259700 499100
rect 259756 484036 259812 516684
rect 259756 483970 259812 483980
rect 259868 500948 259924 500958
rect 259868 469476 259924 500892
rect 261212 482356 261268 571340
rect 261660 511588 261716 511598
rect 261212 482290 261268 482300
rect 261324 500836 261380 500846
rect 259868 469410 259924 469420
rect 261324 435876 261380 500780
rect 261548 499380 261604 499390
rect 261436 497812 261492 497822
rect 261436 436996 261492 497756
rect 261548 458276 261604 499324
rect 261660 477316 261716 511532
rect 261772 508228 261828 508238
rect 261772 492436 261828 508172
rect 261772 492370 261828 492380
rect 262892 500724 262948 500734
rect 261660 477250 261716 477260
rect 261548 458210 261604 458220
rect 261436 436930 261492 436940
rect 261660 437780 261716 437790
rect 261324 435810 261380 435820
rect 261212 430276 261268 430286
rect 259644 427410 259700 427420
rect 259756 428820 259812 428830
rect 259756 410116 259812 428764
rect 259756 410050 259812 410060
rect 261212 379876 261268 430220
rect 261324 426804 261380 426814
rect 261324 388836 261380 426748
rect 261660 416836 261716 437724
rect 262892 417956 262948 500668
rect 263004 487956 263060 571452
rect 264572 570500 264628 570510
rect 263116 569828 263172 569838
rect 263116 496356 263172 569772
rect 263788 530516 263844 530526
rect 263788 527828 263844 530460
rect 263788 527762 263844 527772
rect 264572 506996 264628 570444
rect 265132 528164 265188 528174
rect 264572 506930 264628 506940
rect 264684 513268 264740 513278
rect 263116 496290 263172 496300
rect 263228 499492 263284 499502
rect 263004 487890 263060 487900
rect 263228 459396 263284 499436
rect 264572 498148 264628 498158
rect 264572 488516 264628 498092
rect 264572 488450 264628 488460
rect 264684 480676 264740 513212
rect 264684 480610 264740 480620
rect 264796 506660 264852 506670
rect 263900 480452 263956 480462
rect 263788 479668 263844 479678
rect 263788 478436 263844 479612
rect 263788 478370 263844 478380
rect 263900 474516 263956 480396
rect 263900 474450 263956 474460
rect 264796 473956 264852 506604
rect 265020 506548 265076 506558
rect 264908 503188 264964 503198
rect 264908 475636 264964 503132
rect 265020 480116 265076 506492
rect 265132 500836 265188 528108
rect 265132 500770 265188 500780
rect 265132 496468 265188 496478
rect 265132 485716 265188 496412
rect 265132 485650 265188 485660
rect 265020 480050 265076 480060
rect 264908 475570 264964 475580
rect 264796 473890 264852 473900
rect 263788 472276 263844 472286
rect 263788 468692 263844 472220
rect 263788 468626 263844 468636
rect 263228 459330 263284 459340
rect 264572 447860 264628 447870
rect 264572 430276 264628 447804
rect 265132 441252 265188 441262
rect 264572 430210 264628 430220
rect 265020 437892 265076 437902
rect 262892 417890 262948 417900
rect 263004 430164 263060 430174
rect 261660 416770 261716 416780
rect 261324 388770 261380 388780
rect 261436 411236 261492 411246
rect 261436 385588 261492 411180
rect 261436 385522 261492 385532
rect 263004 380996 263060 430108
rect 264684 429268 264740 429278
rect 264572 427700 264628 427710
rect 263116 426132 263172 426142
rect 263116 407876 263172 426076
rect 263116 407810 263172 407820
rect 264572 389396 264628 427644
rect 264684 398916 264740 429212
rect 264684 398850 264740 398860
rect 264796 427588 264852 427598
rect 264572 389330 264628 389340
rect 264796 388276 264852 427532
rect 264908 426692 264964 426702
rect 264908 397236 264964 426636
rect 265020 415716 265076 437836
rect 265132 426916 265188 441196
rect 265356 439684 265412 439694
rect 265356 428036 265412 439628
rect 265356 427970 265412 427980
rect 265132 426850 265188 426860
rect 265020 415650 265076 415660
rect 264908 397170 264964 397180
rect 264796 388210 264852 388220
rect 263004 380930 263060 380940
rect 263788 383124 263844 383134
rect 261212 379810 261268 379820
rect 261436 380548 261492 380558
rect 259532 379250 259588 379260
rect 247772 359090 247828 359100
rect 229516 358372 229572 358382
rect 158844 358260 158900 358270
rect 97468 358148 97524 358158
rect 81452 356356 81508 356366
rect 81452 303156 81508 356300
rect 97468 355880 97524 358092
rect 122668 358148 122724 358158
rect 100828 358036 100884 358046
rect 99484 356356 99540 356366
rect 99484 355880 99540 356300
rect 100828 355880 100884 357980
rect 104188 357924 104244 357934
rect 104188 355880 104244 357868
rect 108220 356468 108276 356478
rect 108220 355880 108276 356412
rect 107548 355684 107604 355694
rect 107548 355618 107604 355628
rect 104860 355460 104916 355470
rect 104860 355394 104916 355404
rect 122668 353892 122724 358092
rect 122668 353826 122724 353836
rect 138572 358036 138628 358046
rect 99484 306516 99540 314104
rect 100156 313908 100212 314104
rect 100156 313842 100212 313852
rect 101500 307076 101556 314104
rect 104188 308756 104244 314104
rect 104860 311668 104916 314104
rect 104860 311602 104916 311612
rect 104188 308690 104244 308700
rect 101500 307010 101556 307020
rect 99484 306450 99540 306460
rect 106204 305956 106260 314104
rect 138572 310996 138628 357980
rect 158172 356580 158228 356590
rect 158172 355880 158228 356524
rect 158844 355880 158900 358204
rect 186396 358260 186452 358270
rect 163548 358148 163604 358158
rect 163548 355880 163604 358092
rect 166236 358036 166292 358046
rect 166236 355880 166292 357980
rect 166908 356692 166964 356702
rect 166908 355880 166964 356636
rect 168924 355908 168980 355918
rect 168924 355842 168980 355852
rect 161532 355796 161588 355806
rect 161532 355730 161588 355740
rect 186396 354004 186452 358204
rect 225484 358260 225540 358270
rect 199052 358148 199108 358158
rect 186396 353938 186452 353948
rect 187292 356692 187348 356702
rect 187292 315476 187348 356636
rect 187292 315410 187348 315420
rect 187516 355796 187572 355806
rect 166236 314692 166292 314702
rect 166236 314626 166292 314636
rect 163548 314580 163604 314590
rect 163548 314514 163604 314524
rect 187516 314244 187572 355740
rect 187516 314178 187572 314188
rect 160188 313796 160244 314104
rect 160188 313730 160244 313740
rect 164220 312340 164276 314104
rect 167580 312452 167636 314104
rect 167580 312386 167636 312396
rect 164220 312274 164276 312284
rect 168924 312228 168980 314104
rect 199052 313236 199108 358092
rect 224812 358148 224868 358158
rect 223356 356020 223412 356030
rect 223356 355908 223412 355964
rect 222824 355852 223412 355908
rect 224812 355880 224868 358092
rect 225484 355880 225540 358204
rect 228172 356692 228228 356702
rect 228172 355880 228228 356636
rect 229516 355880 229572 358316
rect 249452 358372 249508 358382
rect 248556 358260 248612 358270
rect 247996 358036 248052 358046
rect 247772 356580 247828 356590
rect 232204 356132 232260 356142
rect 232204 355880 232260 356076
rect 247772 344596 247828 356524
rect 247996 348628 248052 357980
rect 248332 355908 248388 355918
rect 248332 349076 248388 355852
rect 248556 349636 248612 358204
rect 248556 349570 248612 349580
rect 248332 349010 248388 349020
rect 247996 348562 248052 348572
rect 247772 344530 247828 344540
rect 247772 319956 247828 319966
rect 225484 314468 225540 314478
rect 225484 314402 225540 314412
rect 199052 313170 199108 313180
rect 168924 312162 168980 312172
rect 221452 312004 221508 314104
rect 221452 311938 221508 311948
rect 224140 311892 224196 314104
rect 224140 311826 224196 311836
rect 247772 311892 247828 319900
rect 249452 319396 249508 358316
rect 257964 358148 258020 358158
rect 252924 356356 252980 356366
rect 249564 356132 249620 356142
rect 249564 324436 249620 356076
rect 252812 356020 252868 356030
rect 249788 355684 249844 355694
rect 249788 336196 249844 355628
rect 249788 336130 249844 336140
rect 249564 324370 249620 324380
rect 252812 321076 252868 355964
rect 252924 337316 252980 356300
rect 256284 355348 256340 355358
rect 252924 337250 252980 337260
rect 256172 340116 256228 340126
rect 252812 321010 252868 321020
rect 249452 319330 249508 319340
rect 249452 318836 249508 318846
rect 247996 318276 248052 318286
rect 247996 312228 248052 318220
rect 248556 317716 248612 317726
rect 248556 314580 248612 317660
rect 248556 314514 248612 314524
rect 249452 313796 249508 318780
rect 256172 313908 256228 340060
rect 256284 330036 256340 355292
rect 256284 329970 256340 329980
rect 257852 346836 257908 346846
rect 256172 313842 256228 313852
rect 249452 313730 249508 313740
rect 257852 312340 257908 346780
rect 257964 323316 258020 358092
rect 261436 358036 261492 380492
rect 263788 378196 263844 383068
rect 263788 378130 263844 378140
rect 263788 373828 263844 373838
rect 263788 369796 263844 373772
rect 263788 369730 263844 369740
rect 261436 357970 261492 357980
rect 261660 357924 261716 357934
rect 258076 356468 258132 356478
rect 258076 334516 258132 356412
rect 258076 334450 258132 334460
rect 259532 356356 259588 356366
rect 257964 323250 258020 323260
rect 258076 327236 258132 327246
rect 258076 314132 258132 327180
rect 259532 314468 259588 356300
rect 261324 356244 261380 356254
rect 259644 355460 259700 355470
rect 259644 338436 259700 355404
rect 259644 338370 259700 338380
rect 261212 351316 261268 351326
rect 259532 314402 259588 314412
rect 258076 314066 258132 314076
rect 257852 312274 257908 312284
rect 247996 312162 248052 312172
rect 261212 312004 261268 351260
rect 261324 329476 261380 356188
rect 261324 329410 261380 329420
rect 261436 342916 261492 342926
rect 261324 326116 261380 326126
rect 261324 314020 261380 326060
rect 261324 313954 261380 313964
rect 261436 312452 261492 342860
rect 261660 338996 261716 357868
rect 263788 356692 263844 356702
rect 263788 353556 263844 356636
rect 264572 355572 264628 355582
rect 263788 353490 263844 353500
rect 264460 354004 264516 354014
rect 263788 348628 263844 348638
rect 261660 338930 261716 338940
rect 262892 348516 262948 348526
rect 262892 314692 262948 348460
rect 263788 341796 263844 348572
rect 264460 343476 264516 353948
rect 264460 343410 264516 343420
rect 263788 341730 263844 341740
rect 264572 326676 264628 355516
rect 265356 353892 265412 353902
rect 264908 353780 264964 353790
rect 264684 353668 264740 353678
rect 264684 328356 264740 353612
rect 264908 332276 264964 353724
rect 265356 337876 265412 353836
rect 265356 337810 265412 337820
rect 264908 332210 264964 332220
rect 264684 328290 264740 328300
rect 264572 326610 264628 326620
rect 262892 314626 262948 314636
rect 261436 312386 261492 312396
rect 261212 311938 261268 311948
rect 247772 311826 247828 311836
rect 138572 310930 138628 310940
rect 166236 311668 166292 311678
rect 166236 309876 166292 311612
rect 166236 309810 166292 309820
rect 106204 305890 106260 305900
rect 81452 303090 81508 303100
rect 263900 298116 263956 298126
rect 263788 297556 263844 297566
rect 257852 296996 257908 297006
rect 225932 296660 225988 296670
rect 224812 295316 224868 295326
rect 224140 294196 224196 294206
rect 187292 289716 187348 289726
rect 166908 287924 166964 287934
rect 98812 287812 98868 287822
rect 98140 287588 98196 287598
rect 98140 284760 98196 287532
rect 98812 284760 98868 287756
rect 122668 287812 122724 287822
rect 105532 287700 105588 287710
rect 102172 285908 102228 285918
rect 102172 284760 102228 285852
rect 105532 284760 105588 287644
rect 106204 286020 106260 286030
rect 106204 284760 106260 285964
rect 102844 284564 102900 284574
rect 102844 284498 102900 284508
rect 101500 284452 101556 284462
rect 101500 284386 101556 284396
rect 122668 283108 122724 287756
rect 162876 287812 162932 287822
rect 143612 287476 143668 287486
rect 143612 283332 143668 287420
rect 160860 284788 160916 284798
rect 162876 284760 162932 287756
rect 164220 286132 164276 286142
rect 164220 284760 164276 286076
rect 166908 284760 166964 287868
rect 169596 287476 169652 287486
rect 168924 286356 168980 286366
rect 168924 284760 168980 286300
rect 169596 284760 169652 287420
rect 170940 286916 170996 286926
rect 170940 284788 170996 286860
rect 170296 284732 170996 284788
rect 160860 284722 160916 284732
rect 143612 283266 143668 283276
rect 122668 283042 122724 283052
rect 108892 243012 108948 243022
rect 108892 242946 108948 242956
rect 94108 242900 94164 242910
rect 94108 242834 94164 242844
rect 106204 241668 106260 242872
rect 106204 241602 106260 241612
rect 162204 239652 162260 242872
rect 163548 239764 163604 242872
rect 163548 239698 163604 239708
rect 162204 239586 162260 239596
rect 165564 239316 165620 242872
rect 166236 241444 166292 242872
rect 166236 241378 166292 241388
rect 167132 242788 167188 242798
rect 167132 239876 167188 242732
rect 170268 240212 170324 242872
rect 170268 240146 170324 240156
rect 187292 240212 187348 289660
rect 223468 287364 223524 287374
rect 197372 285236 197428 285246
rect 192332 284340 192388 284350
rect 192332 241556 192388 284284
rect 192332 241490 192388 241500
rect 187292 240146 187348 240156
rect 167132 239810 167188 239820
rect 197372 239652 197428 285180
rect 223468 284760 223524 287308
rect 224140 284760 224196 294140
rect 224812 284760 224868 295260
rect 225932 287364 225988 296604
rect 228844 296436 228900 296446
rect 225932 287298 225988 287308
rect 228172 287364 228228 287374
rect 228172 284760 228228 287308
rect 228844 284760 228900 296380
rect 230860 294868 230916 294878
rect 230860 284760 230916 294812
rect 232876 291956 232932 291966
rect 232876 284760 232932 291900
rect 249676 288596 249732 288606
rect 247772 287924 247828 287934
rect 247772 256116 247828 287868
rect 248108 287812 248164 287822
rect 248108 267988 248164 287756
rect 248108 267922 248164 267932
rect 249452 286020 249508 286030
rect 247772 256050 247828 256060
rect 248108 267316 248164 267326
rect 248108 243628 248164 267260
rect 249452 249956 249508 285964
rect 249564 284564 249620 284574
rect 249564 276276 249620 284508
rect 249564 276210 249620 276220
rect 249452 249890 249508 249900
rect 249564 265076 249620 265086
rect 248556 246596 248612 246606
rect 247884 243572 248164 243628
rect 248444 246148 248500 246158
rect 222124 243124 222180 243134
rect 222124 243058 222180 243068
rect 222796 240212 222852 242872
rect 222796 240146 222852 240156
rect 197372 239586 197428 239596
rect 230860 239652 230916 242872
rect 247884 240212 247940 243572
rect 247884 240146 247940 240156
rect 248444 239988 248500 246092
rect 248556 241780 248612 246540
rect 249564 243124 249620 265020
rect 249564 243058 249620 243068
rect 248556 241714 248612 241724
rect 248444 239922 248500 239932
rect 230860 239586 230916 239596
rect 165564 239250 165620 239260
rect 249452 239428 249508 239438
rect 225484 233156 225540 233166
rect 199052 232036 199108 232046
rect 195692 230916 195748 230926
rect 166236 229236 166292 229246
rect 163548 228676 163604 228686
rect 158844 226996 158900 227006
rect 133532 224196 133588 224206
rect 105532 219716 105588 219726
rect 102172 219156 102228 219166
rect 101500 215908 101556 215918
rect 83804 215348 83860 215358
rect 83804 210980 83860 215292
rect 98140 215236 98196 215246
rect 98140 213528 98196 215180
rect 99484 215124 99540 215134
rect 98812 213780 98868 213790
rect 98812 213528 98868 213724
rect 99484 213220 99540 215068
rect 101500 213528 101556 215852
rect 102172 213528 102228 219100
rect 104188 217476 104244 217486
rect 103516 215348 103572 215358
rect 103516 213528 103572 215292
rect 104188 213528 104244 217420
rect 105532 213528 105588 219660
rect 106204 218036 106260 218046
rect 106204 213528 106260 217980
rect 106876 215460 106932 215470
rect 106876 213528 106932 215404
rect 99484 213154 99540 213164
rect 102844 212884 102900 212894
rect 102844 212818 102900 212828
rect 83804 210914 83860 210924
rect 125132 211316 125188 211326
rect 102844 171668 102900 171678
rect 100156 171220 100212 171640
rect 102844 171602 102900 171612
rect 100156 171154 100212 171164
rect 125132 169428 125188 211260
rect 133532 171220 133588 224140
rect 141932 216916 141988 216926
rect 141932 171332 141988 216860
rect 158844 213528 158900 226940
rect 159516 215124 159572 215134
rect 159516 213528 159572 215068
rect 163548 213528 163604 228620
rect 164220 215684 164276 215694
rect 164220 213528 164276 215628
rect 166236 213528 166292 229180
rect 186396 215124 186452 215134
rect 166908 213892 166964 213902
rect 166908 213528 166964 213836
rect 160188 212884 160244 212894
rect 160188 212818 160244 212828
rect 186396 211204 186452 215068
rect 186396 211138 186452 211148
rect 186508 174356 186564 174366
rect 185612 173236 185668 173246
rect 164892 171780 164948 171790
rect 164892 171714 164948 171724
rect 141932 171266 141988 171276
rect 133532 171154 133588 171164
rect 125132 169362 125188 169372
rect 162204 169204 162260 171640
rect 162876 169428 162932 171640
rect 166908 171332 166964 171640
rect 166908 171266 166964 171276
rect 162876 169362 162932 169372
rect 167580 170548 167636 170558
rect 162204 169138 162260 169148
rect 125132 166516 125188 166526
rect 88060 159236 88116 159246
rect 81452 158116 81508 158126
rect 81452 101108 81508 158060
rect 88060 142296 88116 159180
rect 105532 150612 105588 150622
rect 102508 143668 102564 143678
rect 102396 143612 102508 143668
rect 102396 142324 102452 143612
rect 102508 143602 102564 143612
rect 102200 142268 102452 142324
rect 102844 143108 102900 143118
rect 102844 142296 102900 143052
rect 105532 142296 105588 150556
rect 106876 144900 106932 144910
rect 106876 142296 106932 144844
rect 99484 142100 99540 142110
rect 98840 142044 99484 142100
rect 99484 142034 99540 142044
rect 98588 141988 98644 141998
rect 98168 141932 98588 141988
rect 98588 141922 98644 141932
rect 125132 101668 125188 166460
rect 130172 165956 130228 165966
rect 125132 101602 125188 101612
rect 125244 160356 125300 160366
rect 81452 101042 81508 101052
rect 99484 100884 99540 100894
rect 99484 100818 99540 100828
rect 102844 100772 102900 100782
rect 102844 100706 102900 100716
rect 106876 100660 106932 100670
rect 106876 100594 106932 100604
rect 101500 100548 101556 100558
rect 101500 100482 101556 100492
rect 104188 98868 104244 100520
rect 104188 98802 104244 98812
rect 104860 98756 104916 100520
rect 105532 98980 105588 100520
rect 105532 98914 105588 98924
rect 104860 98690 104916 98700
rect 125244 98756 125300 160300
rect 130172 100660 130228 165900
rect 135212 162036 135268 162046
rect 133532 154196 133588 154206
rect 133532 100996 133588 154140
rect 133532 100930 133588 100940
rect 130172 100594 130228 100604
rect 135212 98868 135268 161980
rect 162876 150724 162932 150734
rect 161532 147140 161588 147150
rect 161532 142296 161588 147084
rect 162876 142296 162932 150668
rect 164220 147252 164276 147262
rect 164220 142296 164276 147196
rect 167580 142296 167636 170492
rect 168252 169316 168308 171640
rect 168252 169250 168308 169260
rect 168364 170660 168420 170670
rect 168364 142324 168420 170604
rect 185612 147252 185668 173180
rect 186508 170660 186564 174300
rect 195692 171332 195748 230860
rect 199052 171780 199108 231980
rect 222796 215796 222852 215806
rect 222796 213528 222852 215740
rect 223468 215572 223524 215582
rect 223468 213528 223524 215516
rect 225484 213528 225540 233100
rect 228508 215908 228564 215918
rect 228508 214340 228564 215852
rect 228508 214274 228564 214284
rect 228844 215124 228900 215134
rect 228844 213528 228900 215068
rect 247996 215124 248052 215134
rect 226828 212884 226884 212894
rect 226828 212818 226884 212828
rect 231532 212884 231588 212894
rect 231532 212818 231588 212828
rect 247884 212548 247940 212558
rect 247772 207956 247828 207966
rect 246428 172676 246484 172686
rect 199052 171714 199108 171724
rect 230860 171780 230916 171790
rect 230860 171714 230916 171724
rect 195692 171266 195748 171276
rect 223468 171332 223524 171640
rect 223468 171266 223524 171276
rect 186508 170594 186564 170604
rect 200732 170996 200788 171006
rect 185612 147186 185668 147196
rect 187292 170436 187348 170446
rect 168280 142268 168420 142324
rect 160860 100996 160916 101006
rect 160860 100930 160916 100940
rect 165564 100996 165620 101006
rect 165564 100930 165620 100940
rect 169596 100772 169652 100782
rect 169596 100706 169652 100716
rect 187292 100772 187348 170380
rect 192332 142436 192388 142446
rect 187404 141876 187460 141886
rect 187404 101780 187460 141820
rect 187404 101714 187460 101724
rect 187292 100706 187348 100716
rect 170268 100660 170324 100670
rect 170268 100594 170324 100604
rect 192332 100660 192388 142380
rect 192332 100594 192388 100604
rect 135212 98802 135268 98812
rect 125244 98690 125300 98700
rect 166236 98756 166292 100520
rect 168924 98868 168980 100520
rect 168924 98802 168980 98812
rect 166236 98690 166292 98700
rect 200732 98756 200788 170940
rect 225484 169092 225540 171640
rect 226156 169652 226212 171640
rect 228172 171108 228228 171640
rect 229516 171220 229572 171640
rect 229516 171154 229572 171164
rect 228172 171042 228228 171052
rect 226156 169586 226212 169596
rect 225484 169026 225540 169036
rect 204204 165508 204260 165518
rect 200844 140756 200900 140766
rect 200844 100996 200900 140700
rect 200844 100930 200900 100940
rect 204092 100996 204148 101006
rect 200732 98690 200788 98700
rect 135436 97636 135492 97646
rect 110012 96628 110068 96638
rect 106204 91812 106260 91822
rect 104188 86660 104244 86670
rect 98812 78148 98868 78158
rect 83916 74116 83972 74126
rect 83916 71876 83972 74060
rect 83916 71810 83972 71820
rect 98812 71064 98868 78092
rect 100828 74900 100884 74910
rect 100156 74788 100212 74798
rect 100156 71064 100212 74732
rect 100828 71064 100884 74844
rect 102844 73556 102900 73566
rect 102844 71064 102900 73500
rect 104188 71064 104244 86604
rect 105532 74676 105588 74686
rect 105532 71064 105588 74620
rect 106204 71064 106260 91756
rect 110012 74900 110068 96572
rect 135436 79828 135492 97580
rect 167356 95396 167412 95406
rect 165564 90132 165620 90142
rect 135436 79762 135492 79772
rect 160860 86772 160916 86782
rect 110012 74834 110068 74844
rect 125132 79156 125188 79166
rect 122668 31332 122724 31342
rect 78092 28354 78148 28364
rect 74732 26786 74788 26796
rect 73052 26562 73108 26572
rect 62972 26450 63028 26460
rect 89404 26516 89460 29288
rect 103516 26628 103572 29288
rect 103516 26562 103572 26572
rect 89404 26450 89460 26460
rect 61292 26338 61348 26348
rect 104188 26404 104244 29288
rect 107548 26852 107604 29288
rect 107548 26786 107604 26796
rect 104188 26338 104244 26348
rect 122668 26404 122724 31276
rect 125132 26852 125188 79100
rect 134428 76356 134484 76366
rect 134428 74788 134484 76300
rect 134428 74722 134484 74732
rect 160860 71064 160916 86716
rect 162876 79828 162932 79838
rect 162876 71064 162932 79772
rect 163548 74788 163604 74798
rect 163548 71064 163604 74732
rect 165564 71064 165620 90076
rect 167356 84980 167412 95340
rect 167356 84914 167412 84924
rect 168252 88452 168308 88462
rect 167132 84756 167188 84766
rect 167132 74788 167188 84700
rect 167132 74722 167188 74732
rect 168252 71064 168308 88396
rect 187292 81956 187348 81966
rect 160860 28308 160916 29288
rect 160860 28242 160916 28252
rect 125132 26786 125188 26796
rect 122668 26338 122724 26348
rect 167580 26292 167636 29288
rect 169596 26404 169652 29288
rect 187292 28308 187348 81900
rect 187292 28242 187348 28252
rect 204092 26516 204148 100940
rect 204204 98868 204260 165452
rect 230188 160468 230244 160478
rect 228172 158788 228228 158798
rect 204204 98802 204260 98812
rect 205772 150388 205828 150398
rect 204092 26450 204148 26460
rect 205772 26516 205828 150332
rect 226156 148596 226212 148606
rect 224812 145796 224868 145806
rect 224812 142296 224868 145740
rect 226156 142296 226212 148540
rect 228172 142296 228228 158732
rect 228844 157108 228900 157118
rect 228844 142296 228900 157052
rect 229516 147252 229572 147262
rect 229516 142296 229572 147196
rect 230188 142296 230244 160412
rect 246428 150724 246484 172620
rect 247772 171108 247828 207900
rect 247884 200116 247940 212492
rect 247996 207396 248052 215068
rect 248556 213668 248612 213678
rect 247996 207330 248052 207340
rect 248108 212436 248164 212446
rect 248108 204036 248164 212380
rect 248556 210196 248612 213612
rect 248556 210130 248612 210140
rect 248108 203970 248164 203980
rect 247884 200050 247940 200060
rect 247772 171042 247828 171052
rect 249452 169652 249508 239372
rect 249676 239316 249732 288540
rect 256172 287588 256228 287598
rect 252924 287364 252980 287374
rect 252812 284452 252868 284462
rect 249788 249396 249844 249406
rect 249788 243012 249844 249340
rect 252812 248276 252868 284396
rect 252924 263956 252980 287308
rect 252924 263890 252980 263900
rect 252812 248210 252868 248220
rect 252924 258916 252980 258926
rect 249788 242946 249844 242956
rect 252924 239764 252980 258860
rect 256172 252196 256228 287532
rect 256284 285908 256340 285918
rect 256284 277956 256340 285852
rect 256284 277890 256340 277900
rect 256172 252130 256228 252140
rect 256284 273812 256340 273822
rect 253036 247716 253092 247726
rect 253036 241668 253092 247660
rect 253036 241602 253092 241612
rect 256284 240100 256340 273756
rect 256284 240034 256340 240044
rect 252924 239698 252980 239708
rect 257852 239652 257908 296940
rect 263788 296660 263844 297500
rect 263788 296594 263844 296604
rect 263900 294868 263956 298060
rect 263900 294802 263956 294812
rect 259532 288260 259588 288270
rect 258636 287700 258692 287710
rect 258076 286132 258132 286142
rect 257964 278516 258020 278526
rect 257964 242900 258020 278460
rect 258076 254996 258132 286076
rect 258636 280196 258692 287644
rect 258636 280130 258692 280140
rect 258076 254930 258132 254940
rect 259532 246036 259588 288204
rect 259532 245970 259588 245980
rect 261212 286020 261268 286030
rect 261212 243796 261268 285964
rect 261436 285796 261492 285806
rect 261212 243730 261268 243740
rect 261324 273476 261380 273486
rect 257964 242834 258020 242844
rect 261324 241892 261380 273420
rect 261436 268996 261492 285740
rect 262892 284788 262948 284798
rect 262892 278908 262948 284732
rect 264908 284228 264964 284238
rect 264572 283108 264628 283118
rect 262892 278852 263060 278908
rect 261436 268930 261492 268940
rect 262892 274596 262948 274606
rect 261324 241826 261380 241836
rect 261548 260596 261604 260606
rect 261548 241444 261604 260540
rect 261548 241378 261604 241388
rect 257852 239586 257908 239596
rect 262892 239540 262948 274540
rect 263004 254436 263060 278852
rect 263004 254370 263060 254380
rect 264572 251636 264628 283052
rect 264572 251570 264628 251580
rect 264684 271236 264740 271246
rect 263788 247156 263844 247166
rect 263788 246148 263844 247100
rect 263788 246082 263844 246092
rect 264684 242788 264740 271180
rect 264684 242722 264740 242732
rect 264796 270116 264852 270126
rect 264796 241108 264852 270060
rect 264908 268436 264964 284172
rect 265020 283332 265076 283342
rect 265020 270676 265076 283276
rect 265020 270610 265076 270620
rect 264908 268370 264964 268380
rect 265132 267988 265188 267998
rect 265132 255556 265188 267932
rect 265132 255490 265188 255500
rect 264796 241042 264852 241052
rect 262892 239474 262948 239484
rect 263788 240436 263844 240446
rect 263788 239428 263844 240380
rect 263788 239362 263844 239372
rect 249676 239250 249732 239260
rect 262892 238196 262948 238206
rect 261212 237636 261268 237646
rect 259532 237076 259588 237086
rect 256284 216020 256340 216030
rect 249676 215796 249732 215806
rect 249564 213556 249620 213566
rect 249564 184436 249620 213500
rect 249676 202916 249732 215740
rect 253036 215684 253092 215694
rect 249676 202850 249732 202860
rect 249788 213780 249844 213790
rect 249788 195076 249844 213724
rect 252812 212660 252868 212670
rect 249900 212324 249956 212334
rect 249900 203476 249956 212268
rect 249900 203410 249956 203420
rect 249788 195010 249844 195020
rect 252812 193956 252868 212604
rect 252812 193890 252868 193900
rect 252924 208516 252980 208526
rect 249564 184370 249620 184380
rect 249676 192276 249732 192286
rect 249452 169586 249508 169596
rect 249564 175476 249620 175486
rect 246428 150658 246484 150668
rect 237692 149156 237748 149166
rect 237692 147252 237748 149100
rect 237692 147186 237748 147196
rect 247772 145012 247828 145022
rect 247772 126868 247828 144956
rect 248108 144900 248164 144910
rect 247996 142884 248052 142894
rect 247996 132020 248052 142828
rect 248108 137396 248164 144844
rect 248108 137330 248164 137340
rect 249452 144676 249508 144686
rect 247996 131964 248276 132020
rect 248108 126868 248164 126878
rect 247772 126812 248108 126868
rect 248108 126802 248164 126812
rect 248220 126196 248276 131964
rect 248332 126196 248388 126206
rect 248220 126140 248332 126196
rect 248332 126130 248388 126140
rect 249452 125636 249508 144620
rect 249452 125570 249508 125580
rect 247996 123508 248052 123518
rect 247884 113428 247940 113438
rect 247772 105028 247828 105038
rect 230188 100772 230244 100782
rect 230188 100706 230244 100716
rect 232876 100772 232932 100782
rect 232876 100706 232932 100716
rect 231532 100660 231588 100670
rect 231532 100594 231588 100604
rect 227500 98868 227556 100520
rect 227500 98802 227556 98812
rect 232204 98756 232260 100520
rect 232204 98690 232260 98700
rect 229516 95060 229572 95070
rect 228172 94948 228228 94958
rect 226716 93716 226772 93726
rect 226716 90020 226772 93660
rect 226716 89954 226772 89964
rect 227612 90356 227668 90366
rect 225484 89796 225540 89806
rect 224140 75012 224196 75022
rect 223468 74900 223524 74910
rect 223468 71064 223524 74844
rect 224140 71064 224196 74956
rect 224812 74788 224868 74798
rect 224812 71064 224868 74732
rect 225484 71064 225540 89740
rect 225932 88676 225988 88686
rect 225932 74900 225988 88620
rect 225932 74834 225988 74844
rect 227612 74788 227668 90300
rect 227612 74722 227668 74732
rect 228172 71064 228228 94892
rect 228844 74900 228900 74910
rect 228844 71064 228900 74844
rect 229516 71064 229572 95004
rect 232204 84980 232260 84990
rect 232204 71064 232260 84924
rect 226828 29876 226884 29886
rect 226828 29810 226884 29820
rect 230188 29316 230244 29326
rect 222124 28308 222180 29288
rect 222124 28242 222180 28252
rect 227500 26852 227556 29288
rect 230188 29250 230244 29260
rect 231532 28196 231588 29288
rect 231532 28130 231588 28140
rect 227500 26786 227556 26796
rect 247772 26852 247828 104972
rect 247884 74788 247940 113372
rect 247996 99092 248052 123452
rect 249452 122276 249508 122286
rect 247996 99026 248052 99036
rect 248108 108388 248164 108398
rect 248108 74900 248164 108332
rect 248108 74834 248164 74844
rect 247884 74722 247940 74732
rect 248332 74228 248388 74238
rect 248332 66836 248388 74172
rect 248332 66770 248388 66780
rect 249452 29876 249508 122220
rect 249564 100772 249620 175420
rect 249676 171668 249732 192220
rect 249676 171602 249732 171612
rect 252812 177156 252868 177166
rect 252700 139188 252756 139198
rect 252700 138964 252756 139132
rect 252700 138898 252756 138908
rect 249564 100706 249620 100716
rect 249676 115556 249732 115566
rect 249452 29810 249508 29820
rect 249564 90916 249620 90926
rect 249564 28196 249620 90860
rect 249676 86772 249732 115500
rect 252812 100660 252868 177100
rect 252924 169092 252980 208460
rect 253036 199556 253092 215628
rect 254492 213892 254548 213902
rect 254492 201236 254548 213836
rect 254492 201170 254548 201180
rect 256172 202356 256228 202366
rect 253036 199490 253092 199500
rect 256172 169204 256228 202300
rect 256284 187796 256340 215964
rect 256508 215572 256564 215582
rect 256508 204596 256564 215516
rect 256508 204530 256564 204540
rect 258188 215348 258244 215358
rect 258188 194516 258244 215292
rect 258188 194450 258244 194460
rect 256284 187730 256340 187740
rect 257852 180516 257908 180526
rect 256172 169138 256228 169148
rect 256284 174916 256340 174926
rect 252924 169026 252980 169036
rect 256284 160468 256340 174860
rect 256284 160402 256340 160412
rect 256172 143108 256228 143118
rect 256172 135716 256228 143052
rect 256172 135650 256228 135660
rect 254492 132916 254548 132926
rect 252812 100594 252868 100604
rect 252924 114996 252980 115006
rect 249676 86706 249732 86716
rect 249788 100436 249844 100446
rect 249564 28130 249620 28140
rect 247772 26786 247828 26796
rect 249788 26740 249844 100380
rect 252812 89236 252868 89246
rect 252700 70532 252756 70542
rect 252700 70084 252756 70476
rect 252700 70018 252756 70028
rect 252812 29204 252868 89180
rect 252924 88452 252980 114940
rect 253036 110516 253092 110526
rect 253036 90132 253092 110460
rect 254492 100548 254548 132860
rect 256284 117236 256340 117246
rect 254492 100482 254548 100492
rect 256172 112756 256228 112766
rect 253036 90066 253092 90076
rect 252924 88386 252980 88396
rect 252812 29138 252868 29148
rect 249788 26674 249844 26684
rect 205772 26450 205828 26460
rect 169596 26338 169652 26348
rect 167580 26226 167636 26236
rect 256172 26292 256228 112700
rect 256284 95060 256340 117180
rect 256284 94994 256340 95004
rect 256396 106596 256452 106606
rect 256396 86660 256452 106540
rect 257852 101780 257908 180460
rect 257964 176596 258020 176606
rect 257964 158788 258020 176540
rect 259532 171332 259588 237020
rect 259756 215460 259812 215470
rect 259532 171266 259588 171276
rect 259644 212436 259700 212446
rect 259644 169540 259700 212380
rect 259756 190596 259812 215404
rect 259756 190530 259812 190540
rect 259644 169474 259700 169484
rect 259756 181076 259812 181086
rect 257964 158722 258020 158732
rect 259756 157108 259812 181020
rect 261212 171780 261268 237580
rect 261548 215236 261604 215246
rect 261436 212996 261492 213006
rect 261212 171714 261268 171724
rect 261324 198436 261380 198446
rect 261324 169428 261380 198380
rect 261436 183316 261492 212940
rect 261548 195636 261604 215180
rect 261548 195570 261604 195580
rect 261436 183250 261492 183260
rect 261324 169362 261380 169372
rect 261436 172116 261492 172126
rect 259756 157042 259812 157052
rect 261436 147140 261492 172060
rect 262892 171220 262948 238140
rect 264572 234388 264628 234398
rect 263116 213444 263172 213454
rect 262892 171154 262948 171164
rect 263004 201796 263060 201806
rect 263004 169316 263060 201740
rect 263116 187236 263172 213388
rect 263788 211204 263844 211214
rect 263788 200676 263844 211148
rect 263788 200610 263844 200620
rect 263116 187170 263172 187180
rect 263228 188916 263284 188926
rect 263004 169250 263060 169260
rect 263228 168980 263284 188860
rect 263788 171556 263844 171566
rect 263788 170548 263844 171500
rect 263788 170482 263844 170492
rect 263228 168914 263284 168924
rect 263788 169316 263844 169326
rect 263788 165508 263844 169260
rect 263788 165442 263844 165452
rect 261548 165396 261604 165406
rect 261548 150612 261604 165340
rect 261548 150546 261604 150556
rect 263004 164836 263060 164846
rect 261436 147074 261492 147084
rect 259644 146132 259700 146142
rect 258076 127652 258132 127662
rect 257852 101714 257908 101724
rect 257964 107716 258020 107726
rect 257068 93156 257124 93166
rect 257068 88228 257124 93100
rect 257068 88162 257124 88172
rect 256396 86594 256452 86604
rect 257964 78148 258020 107660
rect 258076 98980 258132 127596
rect 259532 109284 259588 109294
rect 258076 98914 258132 98924
rect 258188 105476 258244 105486
rect 258188 91812 258244 105420
rect 258188 91746 258244 91756
rect 257964 78082 258020 78092
rect 259532 26404 259588 109228
rect 259644 98868 259700 146076
rect 261436 123396 261492 123406
rect 259644 98802 259700 98812
rect 261212 116676 261268 116686
rect 261212 28308 261268 116620
rect 261324 111076 261380 111086
rect 261324 79828 261380 111020
rect 261436 94948 261492 123340
rect 261436 94882 261492 94892
rect 262892 105364 262948 105374
rect 261324 79762 261380 79772
rect 261212 28242 261268 28252
rect 262892 26628 262948 105308
rect 263004 100884 263060 164780
rect 263788 153636 263844 153646
rect 263788 152068 263844 153580
rect 263788 152002 263844 152012
rect 263004 100818 263060 100828
rect 263116 147812 263172 147822
rect 263116 98756 263172 147756
rect 263788 131796 263844 131806
rect 263788 127652 263844 131740
rect 263788 127586 263844 127596
rect 263900 127316 263956 127326
rect 263788 126868 263844 126878
rect 263788 125076 263844 126812
rect 263788 125010 263844 125020
rect 263900 123508 263956 127260
rect 263900 123442 263956 123452
rect 263116 98690 263172 98700
rect 263228 117796 263284 117806
rect 262892 26562 262948 26572
rect 263116 91588 263172 91598
rect 263116 26628 263172 91532
rect 263228 84980 263284 117740
rect 263788 112196 263844 112206
rect 263788 109284 263844 112140
rect 263788 109218 263844 109228
rect 263788 102676 263844 102686
rect 263788 96628 263844 102620
rect 263788 96562 263844 96572
rect 263788 94276 263844 94286
rect 263788 93380 263844 94220
rect 263788 93314 263844 93324
rect 263228 84914 263284 84924
rect 264572 28308 264628 234332
rect 264684 215236 264740 215246
rect 264684 173908 264740 215180
rect 264908 214340 264964 214350
rect 264796 210868 264852 210878
rect 264796 182756 264852 210812
rect 264908 192836 264964 214284
rect 264908 192770 264964 192780
rect 265020 210980 265076 210990
rect 265020 186116 265076 210924
rect 265020 186050 265076 186060
rect 264796 182690 264852 182700
rect 264684 173842 264740 173852
rect 264684 143668 264740 143678
rect 264684 131236 264740 143612
rect 265132 141988 265188 141998
rect 264908 141764 264964 141774
rect 264908 132356 264964 141708
rect 265132 135156 265188 141932
rect 265356 141988 265412 141998
rect 265356 141652 265412 141932
rect 265356 141586 265412 141596
rect 265132 135090 265188 135100
rect 264908 132290 264964 132300
rect 264684 131170 264740 131180
rect 264684 123956 264740 123966
rect 264684 105028 264740 123900
rect 264908 119476 264964 119486
rect 264796 118916 264852 118926
rect 264796 108388 264852 118860
rect 264908 113428 264964 119420
rect 264908 113362 264964 113372
rect 264796 108322 264852 108332
rect 265020 108276 265076 108286
rect 265020 105364 265076 108220
rect 265020 105298 265076 105308
rect 264684 104962 264740 104972
rect 266252 93268 266308 572348
rect 277004 571956 277060 571966
rect 268156 571844 268212 571854
rect 267932 571732 267988 571742
rect 266476 571508 266532 571518
rect 266364 568708 266420 568718
rect 266364 431956 266420 568652
rect 266364 431890 266420 431900
rect 266252 93202 266308 93212
rect 266364 361284 266420 361294
rect 264684 78596 264740 78606
rect 264684 31332 264740 78540
rect 264684 31266 264740 31276
rect 264908 66276 264964 66286
rect 264908 31220 264964 66220
rect 264908 31154 264964 31164
rect 264572 28242 264628 28252
rect 265468 31108 265524 31118
rect 265468 26740 265524 31052
rect 266364 29204 266420 361228
rect 266476 234500 266532 571452
rect 266588 569492 266644 569502
rect 266588 304948 266644 569436
rect 266588 304882 266644 304892
rect 267932 296548 267988 571676
rect 268156 516628 268212 571788
rect 275884 571620 275940 571630
rect 273644 570612 273700 570622
rect 269164 570164 269220 570174
rect 269164 569464 269220 570108
rect 273644 569464 273700 570556
rect 274764 570276 274820 570286
rect 274764 569464 274820 570220
rect 275884 569464 275940 571564
rect 277004 569464 277060 571900
rect 278124 569464 278180 575372
rect 279244 569464 279300 582092
rect 280364 577108 280420 577118
rect 280364 569464 280420 577052
rect 283724 576212 283780 576222
rect 281484 575540 281540 575550
rect 281484 569464 281540 575484
rect 282604 574420 282660 574430
rect 282604 569464 282660 574364
rect 283724 569464 283780 576156
rect 284732 574532 284788 590604
rect 288092 590660 288148 590670
rect 287084 590548 287140 590558
rect 284732 574466 284788 574476
rect 284844 577220 284900 577230
rect 284844 569464 284900 577164
rect 285964 574532 286020 574542
rect 285964 569464 286020 574476
rect 287084 569464 287140 590492
rect 288092 574420 288148 590604
rect 289772 590548 289828 590558
rect 288092 574354 288148 574364
rect 288204 583828 288260 583838
rect 288204 569464 288260 583772
rect 289772 576212 289828 590492
rect 297836 590548 297892 595560
rect 297836 590482 297892 590492
rect 303212 590548 303268 590558
rect 289772 576146 289828 576156
rect 303212 575540 303268 590492
rect 303212 575474 303268 575484
rect 305004 588644 305060 588654
rect 299404 572292 299460 572302
rect 296492 572068 296548 572078
rect 296492 570724 296548 572012
rect 296492 570658 296548 570668
rect 298284 570724 298340 570734
rect 294924 570500 294980 570510
rect 292684 570388 292740 570398
rect 290444 569828 290500 569838
rect 290444 569464 290500 569772
rect 292684 569464 292740 570332
rect 293804 569828 293860 569838
rect 293804 569464 293860 569772
rect 294924 569464 294980 570444
rect 296044 569940 296100 569950
rect 296044 569464 296100 569884
rect 296940 569716 296996 569726
rect 291564 569268 291620 569278
rect 296940 569268 296996 569660
rect 298284 569464 298340 570668
rect 299404 569464 299460 572236
rect 303660 569604 303716 569614
rect 303660 569492 303716 569548
rect 303660 569436 303912 569492
rect 305004 569464 305060 588588
rect 307244 583828 307300 583838
rect 306124 573860 306180 573870
rect 306124 569464 306180 573804
rect 307244 569464 307300 583772
rect 311724 582260 311780 582270
rect 309484 578900 309540 578910
rect 308364 577220 308420 577230
rect 308364 569464 308420 577164
rect 309484 569464 309540 578844
rect 310604 574084 310660 574094
rect 310604 569464 310660 574028
rect 311724 569464 311780 582204
rect 341964 578900 342020 595560
rect 364028 590660 364084 595560
rect 364028 590594 364084 590604
rect 407372 591332 407428 591342
rect 341964 578834 342020 578844
rect 315084 578788 315140 578798
rect 312844 573972 312900 573982
rect 312844 569464 312900 573916
rect 313964 573748 314020 573758
rect 313964 569464 314020 573692
rect 315084 569464 315140 578732
rect 407372 577220 407428 591276
rect 408268 591332 408324 595560
rect 408268 591266 408324 591276
rect 430220 590548 430276 595560
rect 430220 590482 430276 590492
rect 432572 590548 432628 590558
rect 407372 577154 407428 577164
rect 432572 577108 432628 590492
rect 474348 583828 474404 595560
rect 496412 590548 496468 595560
rect 496412 590482 496468 590492
rect 499772 590548 499828 590558
rect 474348 583762 474404 583772
rect 499772 582148 499828 590492
rect 499772 582082 499828 582092
rect 432572 577042 432628 577052
rect 540540 573860 540596 595560
rect 562604 590548 562660 595560
rect 562604 590482 562660 590492
rect 540540 573794 540596 573804
rect 328524 572404 328580 572414
rect 325164 572068 325220 572078
rect 315756 571956 315812 571966
rect 315756 570052 315812 571900
rect 315756 569986 315812 569996
rect 317324 571844 317380 571854
rect 315868 569604 315924 569614
rect 315868 569492 315924 569548
rect 315868 569436 316232 569492
rect 317324 569464 317380 571788
rect 324044 571284 324100 571294
rect 322924 569492 322980 569502
rect 324044 569464 324100 571228
rect 325164 569464 325220 572012
rect 327404 571732 327460 571742
rect 326284 571508 326340 571518
rect 326284 569464 326340 571452
rect 327404 569464 327460 571676
rect 328524 569464 328580 572348
rect 335244 572292 335300 572302
rect 329644 572180 329700 572190
rect 329644 569464 329700 572124
rect 330764 571284 330820 571294
rect 330764 569464 330820 571228
rect 333676 570276 333732 570286
rect 333452 570164 333508 570174
rect 322924 569426 322980 569436
rect 317772 569380 317828 569390
rect 317828 569324 318472 569380
rect 317772 569314 317828 569324
rect 296940 569212 297192 569268
rect 291564 569202 291620 569212
rect 320684 569156 320740 569166
rect 320684 569090 320740 569100
rect 321804 569044 321860 569054
rect 321804 568978 321860 568988
rect 270284 568932 270340 568942
rect 270284 568866 270340 568876
rect 271404 568932 271460 568942
rect 271404 568866 271460 568876
rect 272524 568932 272580 568942
rect 272524 568866 272580 568876
rect 289324 568932 289380 568942
rect 289324 568866 289380 568876
rect 300524 568932 300580 568942
rect 300524 568866 300580 568876
rect 301644 568932 301700 568942
rect 301644 568866 301700 568876
rect 302764 568932 302820 568942
rect 302764 568866 302820 568876
rect 319564 568932 319620 568942
rect 319564 568866 319620 568876
rect 268156 516562 268212 516572
rect 267932 296482 267988 296492
rect 333452 245028 333508 570108
rect 333564 567812 333620 567822
rect 333564 284676 333620 567756
rect 333676 443268 333732 570220
rect 335132 568596 335188 568606
rect 334460 518420 334516 518430
rect 334460 514276 334516 518364
rect 334460 514210 334516 514220
rect 335132 509348 335188 568540
rect 335244 521668 335300 572236
rect 338716 571956 338772 571966
rect 336924 571844 336980 571854
rect 335468 571620 335524 571630
rect 335468 528388 335524 571564
rect 336812 570500 336868 570510
rect 335468 528322 335524 528332
rect 335916 530068 335972 530078
rect 335916 527156 335972 530012
rect 335916 527090 335972 527100
rect 335916 526708 335972 526718
rect 335916 524916 335972 526652
rect 335916 524850 335972 524860
rect 335244 521602 335300 521612
rect 335132 509282 335188 509292
rect 335244 514948 335300 514958
rect 335132 501620 335188 501630
rect 335132 482916 335188 501564
rect 335244 490756 335300 514892
rect 335244 490690 335300 490700
rect 335132 482850 335188 482860
rect 335580 484708 335636 484718
rect 335580 475636 335636 484652
rect 335580 475570 335636 475580
rect 335132 472836 335188 472846
rect 334460 472276 334516 472286
rect 334460 469588 334516 472220
rect 334460 469522 334516 469532
rect 335132 453572 335188 472780
rect 335132 453506 335188 453516
rect 333676 443202 333732 443212
rect 335804 444388 335860 444398
rect 334460 439348 334516 439358
rect 334460 435316 334516 439292
rect 334460 435250 334516 435260
rect 335132 437780 335188 437790
rect 334460 426580 334516 426590
rect 334460 422436 334516 426524
rect 334460 422370 334516 422380
rect 335132 415716 335188 437724
rect 335804 436996 335860 444332
rect 335804 436930 335860 436940
rect 335244 434308 335300 434318
rect 335244 417956 335300 434252
rect 335244 417890 335300 417900
rect 335468 432740 335524 432750
rect 335468 416836 335524 432684
rect 335468 416770 335524 416780
rect 335132 415650 335188 415660
rect 335132 414036 335188 414046
rect 335132 387604 335188 413980
rect 335132 387538 335188 387548
rect 335356 410676 335412 410686
rect 335356 387380 335412 410620
rect 335580 408436 335636 408446
rect 335580 387492 335636 408380
rect 335580 387426 335636 387436
rect 336028 388836 336084 388846
rect 335356 387314 335412 387324
rect 336028 385700 336084 388780
rect 336028 385634 336084 385644
rect 335916 384916 335972 384926
rect 335916 383908 335972 384860
rect 335916 383842 335972 383852
rect 335916 362180 335972 362190
rect 335916 359156 335972 362124
rect 335916 359090 335972 359100
rect 334348 356244 334404 356254
rect 334348 353556 334404 356188
rect 335132 355684 335188 355694
rect 334348 353490 334404 353500
rect 334460 353668 334516 353678
rect 334460 349636 334516 353612
rect 334460 349570 334516 349580
rect 335132 346276 335188 355628
rect 335132 346210 335188 346220
rect 335244 353892 335300 353902
rect 335132 338548 335188 338558
rect 334460 325556 334516 325566
rect 334460 314244 334516 325500
rect 334460 314178 334516 314188
rect 335132 300356 335188 338492
rect 335244 316036 335300 353836
rect 335468 353780 335524 353790
rect 335244 315970 335300 315980
rect 335356 350196 335412 350206
rect 335356 314692 335412 350140
rect 335468 348516 335524 353724
rect 335468 348450 335524 348460
rect 335356 314626 335412 314636
rect 335468 321076 335524 321086
rect 335468 313348 335524 321020
rect 335468 313282 335524 313292
rect 335692 318388 335748 318398
rect 335692 312676 335748 318332
rect 335692 312610 335748 312620
rect 335132 300290 335188 300300
rect 334460 298116 334516 298126
rect 334348 297556 334404 297566
rect 334348 294868 334404 297500
rect 334460 296548 334516 298060
rect 334460 296482 334516 296492
rect 334348 294802 334404 294812
rect 333564 284610 333620 284620
rect 335132 286468 335188 286478
rect 335132 257236 335188 286412
rect 336028 284228 336084 284238
rect 336028 279076 336084 284172
rect 336028 279010 336084 279020
rect 335132 257170 335188 257180
rect 335244 266756 335300 266766
rect 333452 244962 333508 244972
rect 335244 239652 335300 266700
rect 335468 265636 335524 265646
rect 335356 263396 335412 263406
rect 335356 246148 335412 263340
rect 335356 246082 335412 246092
rect 335468 240100 335524 265580
rect 335468 240034 335524 240044
rect 335244 239586 335300 239596
rect 266476 234434 266532 234444
rect 334348 239316 334404 239326
rect 334348 232708 334404 239260
rect 334460 238196 334516 238206
rect 334460 236068 334516 238140
rect 334460 236002 334516 236012
rect 334348 232642 334404 232652
rect 336812 231924 336868 570444
rect 336924 485156 336980 571788
rect 337148 571732 337204 571742
rect 336924 485090 336980 485100
rect 337036 498260 337092 498270
rect 337036 453236 337092 498204
rect 337148 486276 337204 571676
rect 338492 571508 338548 571518
rect 337596 531636 337652 531646
rect 337596 525812 337652 531580
rect 337596 525746 337652 525756
rect 337148 486210 337204 486220
rect 337260 503748 337316 503758
rect 337260 477876 337316 503692
rect 337708 503188 337764 503198
rect 337708 500836 337764 503132
rect 337708 500770 337764 500780
rect 337260 477810 337316 477820
rect 338492 476756 338548 571452
rect 338492 476690 338548 476700
rect 338604 500836 338660 500846
rect 338492 470036 338548 470046
rect 338492 453348 338548 469980
rect 338492 453282 338548 453292
rect 337036 453170 337092 453180
rect 336924 430388 336980 430398
rect 336924 407316 336980 430332
rect 336924 407250 336980 407260
rect 338492 426916 338548 426926
rect 338492 400036 338548 426860
rect 338604 418516 338660 500780
rect 338716 494676 338772 571900
rect 557564 571956 557620 571966
rect 433468 571844 433524 571854
rect 351932 571620 351988 571630
rect 341852 571396 341908 571406
rect 340172 570388 340228 570398
rect 339276 511812 339332 511822
rect 339276 508676 339332 511756
rect 339276 508610 339332 508620
rect 338716 494610 338772 494620
rect 338828 499380 338884 499390
rect 338828 443716 338884 499324
rect 338828 443650 338884 443660
rect 338604 418450 338660 418460
rect 338716 430276 338772 430286
rect 338716 406756 338772 430220
rect 338716 406690 338772 406700
rect 338492 399970 338548 399980
rect 339276 358708 339332 358718
rect 337148 357140 337204 357150
rect 336924 356804 336980 356814
rect 336924 304836 336980 356748
rect 337148 313796 337204 357084
rect 339276 356244 339332 358652
rect 339276 356178 339332 356188
rect 338604 355572 338660 355582
rect 337148 313730 337204 313740
rect 338492 351876 338548 351886
rect 338492 311668 338548 351820
rect 338604 344036 338660 355516
rect 338604 343970 338660 343980
rect 338492 311602 338548 311612
rect 336924 304770 336980 304780
rect 338604 287364 338660 287374
rect 338492 271796 338548 271806
rect 336924 260484 336980 260494
rect 336924 239764 336980 260428
rect 338492 243348 338548 271740
rect 338604 265076 338660 287308
rect 338716 285684 338772 285694
rect 338716 267876 338772 285628
rect 338716 267810 338772 267820
rect 338604 265010 338660 265020
rect 338492 243282 338548 243292
rect 336924 239698 336980 239708
rect 336812 231858 336868 231868
rect 338492 237636 338548 237646
rect 338492 227668 338548 237580
rect 338492 227602 338548 227612
rect 336812 215796 336868 215806
rect 335244 215684 335300 215694
rect 335132 208516 335188 208526
rect 335132 178052 335188 208460
rect 335244 207396 335300 215628
rect 335244 207330 335300 207340
rect 335356 211092 335412 211102
rect 335132 177986 335188 177996
rect 335244 202916 335300 202926
rect 335244 174020 335300 202860
rect 335356 198436 335412 211036
rect 335916 210868 335972 210878
rect 335916 205716 335972 210812
rect 335916 205650 335972 205660
rect 335356 198370 335412 198380
rect 335244 173954 335300 173964
rect 335356 179396 335412 179406
rect 335356 172228 335412 179340
rect 335356 172162 335412 172172
rect 336812 171220 336868 215740
rect 338492 215572 338548 215582
rect 338492 195636 338548 215516
rect 339276 213668 339332 213678
rect 339276 209636 339332 213612
rect 339276 209570 339332 209580
rect 338492 195570 338548 195580
rect 336812 171154 336868 171164
rect 338492 188356 338548 188366
rect 338492 169428 338548 188300
rect 338716 178052 338772 178062
rect 338716 169540 338772 177996
rect 338716 169474 338772 169484
rect 338492 169362 338548 169372
rect 334460 168756 334516 168766
rect 334460 167188 334516 168700
rect 334460 167122 334516 167132
rect 336924 168196 336980 168206
rect 336028 154196 336084 154206
rect 336028 150388 336084 154140
rect 336028 150322 336084 150332
rect 334460 148036 334516 148046
rect 334460 147028 334516 147980
rect 334460 146962 334516 146972
rect 335244 143780 335300 143790
rect 335132 140756 335188 140766
rect 334460 140532 334516 140542
rect 334460 139076 334516 140476
rect 334460 139010 334516 139020
rect 334348 113876 334404 113886
rect 334348 107492 334404 113820
rect 335132 110068 335188 140700
rect 335244 137396 335300 143724
rect 336812 142100 336868 142110
rect 335244 137330 335300 137340
rect 335804 140756 335860 140766
rect 335804 135156 335860 140700
rect 335804 135090 335860 135100
rect 335356 134036 335412 134046
rect 335356 113428 335412 133980
rect 336812 129556 336868 142044
rect 336812 129490 336868 129500
rect 335356 113362 335412 113372
rect 335692 116116 335748 116126
rect 335692 112868 335748 116060
rect 335692 112802 335748 112812
rect 335132 110002 335188 110012
rect 334348 107426 334404 107436
rect 336812 107492 336868 107502
rect 267708 101668 267764 101678
rect 267708 101220 267764 101612
rect 267708 101154 267764 101164
rect 335916 79156 335972 79166
rect 335916 78372 335972 79100
rect 335916 78306 335972 78316
rect 335132 77476 335188 77486
rect 334460 68628 334516 68638
rect 334460 67844 334516 68572
rect 334460 67778 334516 67788
rect 335132 31108 335188 77420
rect 335356 72436 335412 72446
rect 335356 59668 335412 72380
rect 335356 59602 335412 59612
rect 335132 31042 335188 31052
rect 270060 29988 270116 29998
rect 270060 29922 270116 29932
rect 274316 29764 274372 29774
rect 274316 29698 274372 29708
rect 278572 29652 278628 29662
rect 278572 29586 278628 29596
rect 282828 29540 282884 29550
rect 282828 29474 282884 29484
rect 291340 29428 291396 29438
rect 291340 29362 291396 29372
rect 295596 29316 295652 29326
rect 266364 29138 266420 29148
rect 287084 28420 287140 29288
rect 295596 29250 295652 29260
rect 299852 28532 299908 29288
rect 304108 29092 304164 29288
rect 304108 29026 304164 29036
rect 299852 28466 299908 28476
rect 287084 28354 287140 28364
rect 308364 28308 308420 29288
rect 308364 28242 308420 28252
rect 265468 26674 265524 26684
rect 263116 26562 263172 26572
rect 312620 26516 312676 29288
rect 316876 26628 316932 29288
rect 321132 26740 321188 29288
rect 321132 26674 321188 26684
rect 316876 26562 316932 26572
rect 312620 26450 312676 26460
rect 259532 26338 259588 26348
rect 256172 26226 256228 26236
rect 10892 26114 10948 26124
rect 325388 26180 325444 29288
rect 325388 26114 325444 26124
rect 4172 24388 4228 24398
rect 4172 22932 4228 24332
rect 329644 24388 329700 29288
rect 336812 26852 336868 107436
rect 336924 100996 336980 168140
rect 339276 153076 339332 153086
rect 339276 152180 339332 153020
rect 340172 152516 340228 570332
rect 341852 531076 341908 571340
rect 350252 571284 350308 571294
rect 341852 531010 341908 531020
rect 345212 570164 345268 570174
rect 340284 521892 340340 521902
rect 340284 480676 340340 521836
rect 342636 516852 342692 516862
rect 342636 511476 342692 516796
rect 342636 511410 342692 511420
rect 342076 507108 342132 507118
rect 340284 480610 340340 480620
rect 340396 500724 340452 500734
rect 340284 469476 340340 469486
rect 340284 453236 340340 469420
rect 340396 468356 340452 500668
rect 340396 468290 340452 468300
rect 341852 499268 341908 499278
rect 340284 453170 340340 453180
rect 341852 448756 341908 499212
rect 341964 497812 342020 497822
rect 341964 467236 342020 497756
rect 342076 478996 342132 507052
rect 345212 502516 345268 570108
rect 345324 568932 345380 568942
rect 345324 506996 345380 568876
rect 345324 506930 345380 506940
rect 349356 555268 349412 555278
rect 346892 503412 346948 503422
rect 345212 502450 345268 502460
rect 345548 503300 345604 503310
rect 342076 478930 342132 478940
rect 345212 501060 345268 501070
rect 341964 467170 342020 467180
rect 342076 469588 342132 469598
rect 342076 453460 342132 469532
rect 342636 466116 342692 466126
rect 342636 457828 342692 466060
rect 342636 457762 342692 457772
rect 342076 453394 342132 453404
rect 341852 448690 341908 448700
rect 345212 432740 345268 501004
rect 345324 499492 345380 499502
rect 345324 445396 345380 499436
rect 345436 498148 345492 498158
rect 345436 465556 345492 498092
rect 345548 482356 345604 503244
rect 346892 486836 346948 503356
rect 346892 486770 346948 486780
rect 348572 499604 348628 499614
rect 345548 482290 345604 482300
rect 348572 467796 348628 499548
rect 348572 467730 348628 467740
rect 349356 483364 349412 555212
rect 350252 484708 350308 571228
rect 350364 569604 350420 569614
rect 350364 506436 350420 569548
rect 350364 506370 350420 506380
rect 350588 508228 350644 508238
rect 350252 484642 350308 484652
rect 350364 500948 350420 500958
rect 345436 465490 345492 465500
rect 345436 464996 345492 465006
rect 345436 453124 345492 464940
rect 345436 453058 345492 453068
rect 345324 445330 345380 445340
rect 345212 432674 345268 432684
rect 345436 444948 345492 444958
rect 345212 430164 345268 430174
rect 340284 428484 340340 428494
rect 340284 404516 340340 428428
rect 342076 426804 342132 426814
rect 340284 404450 340340 404460
rect 341852 426244 341908 426254
rect 341852 393316 341908 426188
rect 342076 406196 342132 426748
rect 342076 406130 342132 406140
rect 341852 393250 341908 393260
rect 341852 389956 341908 389966
rect 341852 384244 341908 389900
rect 341852 384178 341908 384188
rect 345212 361396 345268 430108
rect 345324 428708 345380 428718
rect 345324 394996 345380 428652
rect 345436 421876 345492 444892
rect 345436 421810 345492 421820
rect 349356 411460 349412 483308
rect 350252 463876 350308 463886
rect 350252 455140 350308 463820
rect 350252 455074 350308 455084
rect 350252 446068 350308 446078
rect 350252 417396 350308 446012
rect 350364 422996 350420 500892
rect 350476 499044 350532 499054
rect 350476 446516 350532 498988
rect 350588 492436 350644 508172
rect 350588 492370 350644 492380
rect 351932 489076 351988 571564
rect 374220 571508 374276 571518
rect 370860 571284 370916 571294
rect 370860 569464 370916 571228
rect 374220 569464 374276 571452
rect 407372 571508 407428 571518
rect 380268 570164 380324 570174
rect 374892 569604 374948 569614
rect 374892 569492 374948 569548
rect 374892 569436 375592 569492
rect 380268 569464 380324 570108
rect 352044 569044 352100 569054
rect 352044 504196 352100 568988
rect 372204 569044 372260 569054
rect 372204 568978 372260 568988
rect 377580 568932 377636 568942
rect 377580 568866 377636 568876
rect 400652 567700 400708 567710
rect 393932 567588 393988 567598
rect 357868 527828 357924 527838
rect 357868 527492 357924 527772
rect 357868 527426 357924 527436
rect 368732 523460 368788 523470
rect 356188 521780 356244 521790
rect 356188 516516 356244 521724
rect 356188 516450 356244 516460
rect 368732 505316 368788 523404
rect 370188 507108 370244 527688
rect 370188 507042 370244 507052
rect 372092 523572 372148 523582
rect 372092 505876 372148 523516
rect 372092 505810 372148 505820
rect 368732 505250 368788 505260
rect 352044 504130 352100 504140
rect 372204 503748 372260 527688
rect 372204 503682 372260 503692
rect 376236 503188 376292 527688
rect 376908 523572 376964 527688
rect 376908 523506 376964 523516
rect 377580 523460 377636 527688
rect 377580 523394 377636 523404
rect 379708 523460 379764 523470
rect 379708 520436 379764 523404
rect 379708 520370 379764 520380
rect 381388 516964 381444 516974
rect 381388 515396 381444 516908
rect 381388 515330 381444 515340
rect 376236 503122 376292 503132
rect 370188 501060 370244 501070
rect 368172 499492 368228 499502
rect 352156 499156 352212 499166
rect 351932 489010 351988 489020
rect 352044 497924 352100 497934
rect 351036 462756 351092 462766
rect 351036 457940 351092 462700
rect 351036 457874 351092 457884
rect 351932 462196 351988 462206
rect 351932 455252 351988 462140
rect 351932 455186 351988 455196
rect 352044 448196 352100 497868
rect 352156 466676 352212 499100
rect 368172 498344 368228 499436
rect 369516 499380 369572 499390
rect 368844 499044 368900 499054
rect 368844 498344 368900 498988
rect 369516 498344 369572 499324
rect 370188 498344 370244 501004
rect 372876 500836 372932 500846
rect 372876 498344 372932 500780
rect 374220 499268 374276 499278
rect 374220 498344 374276 499212
rect 376236 497924 376292 497934
rect 376236 497858 376292 497868
rect 352156 466610 352212 466620
rect 352492 463316 352548 463326
rect 352492 456484 352548 463260
rect 352604 461636 352660 461646
rect 352604 456596 352660 461580
rect 352604 456530 352660 456540
rect 352492 456418 352548 456428
rect 352044 448130 352100 448140
rect 350476 446450 350532 446460
rect 369516 437780 369572 456456
rect 369628 451668 369684 451678
rect 369628 445956 369684 451612
rect 370188 446068 370244 456456
rect 370188 446002 370244 446012
rect 372092 452004 372148 452014
rect 369628 445890 369684 445900
rect 371308 444500 371364 444510
rect 371308 442036 371364 444444
rect 371308 441970 371364 441980
rect 369516 437714 369572 437724
rect 372092 434308 372148 451948
rect 373548 452004 373604 456456
rect 373548 451938 373604 451948
rect 374220 451668 374276 456456
rect 374220 451602 374276 451612
rect 375452 451108 375508 451118
rect 375452 436436 375508 451052
rect 377580 444948 377636 456456
rect 377580 444882 377636 444892
rect 375452 436370 375508 436380
rect 372092 434242 372148 434252
rect 350364 422930 350420 422940
rect 351932 430500 351988 430510
rect 350252 417330 350308 417340
rect 348572 408996 348628 409006
rect 345324 394930 345380 394940
rect 345436 400596 345492 400606
rect 345436 385364 345492 400540
rect 347788 391076 347844 391086
rect 347788 385812 347844 391020
rect 347788 385746 347844 385756
rect 345436 385298 345492 385308
rect 348572 384020 348628 408940
rect 348572 383954 348628 383964
rect 345212 361330 345268 361340
rect 342636 360388 342692 360398
rect 342636 358596 342692 360332
rect 342636 358530 342692 358540
rect 340284 358372 340340 358382
rect 340284 301476 340340 358316
rect 341852 358036 341908 358046
rect 340396 333956 340452 333966
rect 340396 313796 340452 333900
rect 341852 324996 341908 357980
rect 348684 357924 348740 357934
rect 341964 356692 342020 356702
rect 341964 330596 342020 356636
rect 345436 356468 345492 356478
rect 345324 355348 345380 355358
rect 341964 330530 342020 330540
rect 345212 347396 345268 347406
rect 341852 324930 341908 324940
rect 340396 313730 340452 313740
rect 341852 318276 341908 318286
rect 341852 313572 341908 318220
rect 345212 314468 345268 347340
rect 345324 331156 345380 355292
rect 345436 344596 345492 356412
rect 345436 344530 345492 344540
rect 345324 331090 345380 331100
rect 348572 339556 348628 339566
rect 345212 314402 345268 314412
rect 345324 323316 345380 323326
rect 341852 313506 341908 313516
rect 345324 312340 345380 323260
rect 348572 313684 348628 339500
rect 348684 338548 348740 357868
rect 349244 355908 349300 355918
rect 349244 355236 349300 355852
rect 349244 355170 349300 355180
rect 348684 338482 348740 338492
rect 349356 341684 349412 411404
rect 350252 403396 350308 403406
rect 350252 385476 350308 403340
rect 350252 385410 350308 385420
rect 350364 397796 350420 397806
rect 350364 384468 350420 397740
rect 350364 384402 350420 384412
rect 350588 390516 350644 390526
rect 350588 384356 350644 390460
rect 350588 384290 350644 384300
rect 351148 387156 351204 387166
rect 351148 384132 351204 387100
rect 351148 384066 351204 384076
rect 351932 362180 351988 430444
rect 374892 430500 374948 430510
rect 374892 427112 374948 430444
rect 376908 430164 376964 430174
rect 376908 427112 376964 430108
rect 352044 426356 352100 426366
rect 352044 405076 352100 426300
rect 352044 405010 352100 405020
rect 352044 402052 352100 402062
rect 352044 384580 352100 401996
rect 352492 391636 352548 391646
rect 352492 385252 352548 391580
rect 352492 385186 352548 385196
rect 352604 389396 352660 389406
rect 352604 385140 352660 389340
rect 370860 385924 370916 385934
rect 370188 385700 370244 385710
rect 370188 385634 370244 385644
rect 352604 385074 352660 385084
rect 352044 384514 352100 384524
rect 368844 384244 368900 385336
rect 369068 385308 369544 385364
rect 369068 385140 369124 385308
rect 369068 385074 369124 385084
rect 370860 384692 370916 385868
rect 374220 385812 374276 385822
rect 374220 385746 374276 385756
rect 372876 385364 372932 385374
rect 370860 384626 370916 384636
rect 368844 384178 368900 384188
rect 352716 383908 352772 383918
rect 352716 383012 352772 383852
rect 352716 382946 352772 382956
rect 351932 362114 351988 362124
rect 372204 359716 372260 385336
rect 372876 385298 372932 385308
rect 373548 383012 373604 385336
rect 374892 384132 374948 385336
rect 375564 384356 375620 385336
rect 376908 384692 376964 385336
rect 376908 384626 376964 384636
rect 375564 384290 375620 384300
rect 374892 384066 374948 384076
rect 373548 382946 373604 382956
rect 377580 360388 377636 385336
rect 393932 363972 393988 567532
rect 395164 504868 395220 504878
rect 395164 496356 395220 504812
rect 395164 496290 395220 496300
rect 398972 501060 399028 501070
rect 394044 451220 394100 451230
rect 394044 434196 394100 451164
rect 394044 434130 394100 434140
rect 398972 426580 399028 501004
rect 400652 430164 400708 567644
rect 407372 495236 407428 571452
rect 412412 571284 412468 571294
rect 412412 501620 412468 571228
rect 430780 571284 430836 571294
rect 412524 570164 412580 570174
rect 412524 510916 412580 570108
rect 412524 510850 412580 510860
rect 414092 569604 414148 569614
rect 414092 509236 414148 569548
rect 430780 569464 430836 571228
rect 433468 569464 433524 571788
rect 474684 571844 474740 571854
rect 438172 571732 438228 571742
rect 435484 570164 435540 570174
rect 435484 569464 435540 570108
rect 435708 569604 435764 569614
rect 435708 569492 435764 569548
rect 435708 569436 436184 569492
rect 438172 569464 438228 571676
rect 464492 571732 464548 571742
rect 428092 516852 428148 527688
rect 428092 516786 428148 516796
rect 414092 509170 414148 509180
rect 430108 503412 430164 527688
rect 430108 503346 430164 503356
rect 434812 503300 434868 527688
rect 435484 521892 435540 527688
rect 435484 521826 435540 521836
rect 436828 516964 436884 527688
rect 440188 518420 440244 527688
rect 440188 518354 440244 518364
rect 436828 516898 436884 516908
rect 442204 511812 442260 527688
rect 464492 514948 464548 571676
rect 471212 570052 471268 570062
rect 471212 523236 471268 569996
rect 471212 523170 471268 523180
rect 474572 569716 474628 569726
rect 464492 514882 464548 514892
rect 442204 511746 442260 511756
rect 434812 503234 434868 503244
rect 412412 501554 412468 501564
rect 436156 501060 436212 501070
rect 407372 495170 407428 495180
rect 407484 500836 407540 500846
rect 407484 438676 407540 500780
rect 412412 499268 412468 499278
rect 412412 457716 412468 499212
rect 432796 499268 432852 499278
rect 432796 498344 432852 499212
rect 436156 498344 436212 501004
rect 438844 500948 438900 500958
rect 438844 498344 438900 500892
rect 464492 499268 464548 499278
rect 434812 498260 434868 498270
rect 434812 498194 434868 498204
rect 412412 457650 412468 457660
rect 430780 456036 430836 456456
rect 430780 455970 430836 455980
rect 407484 438610 407540 438620
rect 412412 447972 412468 447982
rect 412412 434756 412468 447916
rect 412412 434690 412468 434700
rect 464492 431396 464548 499212
rect 464492 431330 464548 431340
rect 400652 430098 400708 430108
rect 412412 430500 412468 430510
rect 407372 426692 407428 426702
rect 398972 426514 399028 426524
rect 399196 426580 399252 426590
rect 399196 382116 399252 426524
rect 399196 382050 399252 382060
rect 404012 426132 404068 426142
rect 404012 368116 404068 426076
rect 407372 370916 407428 426636
rect 407372 370850 407428 370860
rect 404012 368050 404068 368060
rect 412412 365876 412468 430444
rect 436156 430500 436212 430510
rect 435484 428708 435540 428718
rect 435484 427112 435540 428652
rect 436156 427112 436212 430444
rect 467852 430500 467908 430510
rect 462812 428596 462868 428606
rect 436828 427028 436884 427038
rect 436828 426962 436884 426972
rect 438172 427028 438228 427038
rect 438172 426962 438228 426972
rect 430780 384468 430836 385336
rect 430780 384402 430836 384412
rect 462812 378196 462868 428540
rect 467852 382676 467908 430444
rect 467852 382610 467908 382620
rect 462812 378130 462868 378140
rect 412412 365810 412468 365820
rect 393932 363906 393988 363916
rect 377580 360322 377636 360332
rect 372204 359650 372260 359660
rect 402332 358484 402388 358494
rect 370860 358372 370916 358382
rect 348572 313618 348628 313628
rect 348684 322196 348740 322206
rect 345324 312274 345380 312284
rect 348684 312004 348740 322140
rect 348684 311938 348740 311948
rect 340284 301410 340340 301420
rect 340284 288596 340340 288606
rect 340284 241780 340340 288540
rect 341852 287812 341908 287822
rect 340284 241714 340340 241724
rect 340396 262276 340452 262286
rect 340396 239988 340452 262220
rect 341852 243236 341908 287756
rect 342076 287588 342132 287598
rect 342076 249956 342132 287532
rect 348684 285908 348740 285918
rect 345324 284340 345380 284350
rect 345212 281316 345268 281326
rect 342076 249890 342132 249900
rect 342188 277396 342244 277406
rect 341852 243170 341908 243180
rect 342188 243012 342244 277340
rect 342188 242946 342244 242956
rect 345212 241668 345268 281260
rect 345324 276276 345380 284284
rect 345324 276210 345380 276220
rect 348572 280196 348628 280206
rect 345212 241602 345268 241612
rect 347788 246148 347844 246158
rect 340396 239922 340452 239932
rect 347788 239876 347844 246092
rect 348572 243124 348628 280140
rect 348684 277956 348740 285852
rect 348684 277890 348740 277900
rect 348572 243058 348628 243068
rect 349356 268436 349412 341628
rect 350252 358260 350308 358270
rect 350252 318388 350308 358204
rect 352716 358148 352772 358158
rect 352716 356916 352772 358092
rect 352716 356850 352772 356860
rect 369516 357924 369572 357934
rect 352380 356580 352436 356590
rect 352156 356244 352212 356254
rect 351932 356020 351988 356030
rect 351932 349076 351988 355964
rect 351932 349010 351988 349020
rect 350252 318322 350308 318332
rect 350364 347956 350420 347966
rect 350364 314020 350420 347900
rect 351932 346836 351988 346846
rect 350588 328356 350644 328366
rect 350364 313954 350420 313964
rect 350476 319396 350532 319406
rect 350476 312228 350532 319340
rect 350588 314132 350644 328300
rect 351932 314580 351988 346780
rect 351932 314514 351988 314524
rect 352044 342916 352100 342926
rect 350588 314066 350644 314076
rect 352044 313908 352100 342860
rect 352156 332276 352212 356188
rect 352380 341796 352436 356524
rect 369516 355880 369572 357868
rect 370860 355880 370916 358316
rect 393148 358372 393204 358382
rect 372876 356804 372932 356814
rect 372876 355880 372932 356748
rect 378252 356692 378308 356702
rect 374220 356244 374276 356254
rect 374220 355880 374276 356188
rect 378252 355880 378308 356636
rect 374892 355348 374948 355358
rect 374892 355282 374948 355292
rect 393148 353892 393204 358316
rect 393148 353826 393204 353836
rect 398972 356804 399028 356814
rect 352380 341730 352436 341740
rect 352156 332210 352212 332220
rect 352268 332836 352324 332846
rect 352044 313842 352100 313852
rect 352156 317716 352212 317726
rect 350476 312162 350532 312172
rect 352156 311780 352212 317660
rect 352268 313460 352324 332780
rect 359436 314132 359492 314142
rect 359436 314066 359492 314076
rect 352268 313394 352324 313404
rect 352156 311714 352212 311724
rect 370188 303156 370244 314104
rect 370188 303090 370244 303100
rect 372204 302036 372260 314104
rect 373548 303716 373604 314104
rect 374220 313460 374276 314104
rect 374220 313394 374276 313404
rect 376236 304276 376292 314104
rect 398972 310996 399028 356748
rect 398972 310930 399028 310940
rect 400652 356692 400708 356702
rect 400652 310436 400708 356636
rect 400652 310370 400708 310380
rect 402332 309876 402388 358428
rect 439516 358484 439572 358494
rect 410732 357924 410788 357934
rect 404796 314244 404852 314254
rect 404796 311892 404852 314188
rect 404796 311826 404852 311836
rect 402332 309810 402388 309820
rect 410732 308196 410788 357868
rect 435484 357924 435540 357934
rect 432124 356804 432180 356814
rect 410732 308130 410788 308140
rect 412412 356244 412468 356254
rect 412412 307076 412468 356188
rect 430780 356244 430836 356254
rect 430780 355880 430836 356188
rect 432124 355880 432180 356748
rect 435484 355880 435540 357868
rect 436156 356692 436212 356702
rect 436156 355880 436212 356636
rect 439516 355880 439572 358428
rect 430108 309316 430164 314104
rect 430108 309250 430164 309260
rect 412412 307010 412468 307020
rect 430780 306516 430836 314104
rect 433468 308756 433524 314104
rect 434812 313684 434868 314104
rect 434812 313618 434868 313628
rect 436156 312116 436212 314104
rect 436156 312050 436212 312060
rect 437500 311556 437556 314104
rect 444220 313796 444276 314104
rect 444220 313730 444276 313740
rect 437500 311490 437556 311500
rect 474572 311108 474628 569660
rect 474684 521556 474740 571788
rect 501564 571844 501620 571854
rect 498204 571732 498260 571742
rect 496188 571620 496244 571630
rect 476252 569716 476308 569726
rect 474684 521490 474740 521500
rect 474796 569604 474852 569614
rect 474796 517636 474852 569548
rect 476252 525868 476308 569660
rect 492268 569716 492324 569726
rect 492268 569492 492324 569660
rect 494844 569604 494900 569614
rect 494844 569492 494900 569548
rect 492268 569436 492856 569492
rect 494844 569436 495544 569492
rect 496188 569464 496244 571564
rect 498204 569464 498260 571676
rect 500892 570052 500948 570062
rect 500892 569464 500948 569996
rect 501564 569464 501620 571788
rect 533372 571620 533428 571630
rect 533372 530068 533428 571564
rect 555548 571396 555604 571406
rect 533372 530002 533428 530012
rect 536732 571284 536788 571294
rect 476140 525812 476308 525868
rect 475468 523348 475524 523358
rect 475468 519876 475524 523292
rect 476140 520996 476196 525812
rect 476140 520930 476196 520940
rect 475468 519810 475524 519820
rect 474796 517570 474852 517580
rect 493500 508228 493556 527688
rect 494844 521780 494900 527688
rect 498204 523460 498260 527688
rect 498204 523394 498260 523404
rect 499548 523348 499604 527688
rect 536732 526708 536788 571228
rect 554204 571284 554260 571294
rect 554204 569464 554260 571228
rect 555548 569464 555604 571340
rect 557564 569464 557620 571900
rect 558236 571620 558292 571630
rect 558236 569464 558292 571564
rect 558908 571508 558964 571518
rect 558908 569464 558964 571452
rect 590492 570724 590548 570734
rect 580636 570612 580692 570622
rect 580412 569828 580468 569838
rect 539196 529396 539252 529406
rect 539196 527828 539252 529340
rect 539196 527762 539252 527772
rect 556892 527828 556948 527838
rect 556892 527762 556948 527772
rect 559580 527716 559636 527726
rect 536732 526642 536788 526652
rect 554876 525812 554932 527688
rect 557564 527492 557620 527688
rect 559580 527650 559636 527660
rect 557564 527426 557620 527436
rect 554876 525746 554932 525756
rect 562268 525476 562324 527688
rect 562268 525410 562324 525420
rect 499548 523282 499604 523292
rect 494844 521714 494900 521724
rect 493500 508162 493556 508172
rect 563612 504868 563668 527688
rect 564284 524356 564340 527688
rect 564284 524290 564340 524300
rect 563612 504802 563668 504812
rect 536732 501060 536788 501070
rect 476252 500948 476308 500958
rect 474684 497924 474740 497934
rect 474684 458276 474740 497868
rect 474684 458210 474740 458220
rect 476252 439348 476308 500892
rect 498876 500948 498932 500958
rect 493500 499268 493556 499278
rect 493500 498344 493556 499212
rect 498876 498344 498932 500892
rect 530012 500948 530068 500958
rect 492828 498148 492884 498158
rect 492828 498082 492884 498092
rect 494172 497924 494228 497934
rect 494172 497858 494228 497868
rect 496860 457156 496916 457166
rect 496860 457090 496916 457100
rect 494844 456596 494900 456606
rect 494844 456530 494900 456540
rect 496188 456484 496244 456494
rect 493500 455140 493556 456456
rect 493500 455074 493556 455084
rect 494172 451220 494228 456456
rect 496188 456418 496244 456428
rect 498876 453124 498932 456456
rect 498876 453058 498932 453068
rect 494172 451154 494228 451164
rect 499548 447972 499604 456456
rect 501564 455252 501620 456456
rect 501564 455186 501620 455196
rect 499548 447906 499604 447916
rect 530012 440916 530068 500892
rect 530012 440850 530068 440860
rect 533372 497924 533428 497934
rect 476252 439282 476308 439292
rect 533372 437556 533428 497868
rect 536732 444388 536788 501004
rect 558908 501060 558964 501070
rect 558236 500836 558292 500846
rect 554876 500724 554932 500734
rect 554876 498344 554932 500668
rect 556220 499156 556276 499166
rect 556220 498344 556276 499100
rect 558236 498344 558292 500780
rect 558908 498344 558964 501004
rect 562268 500948 562324 500958
rect 562268 498344 562324 500892
rect 562940 499604 562996 499614
rect 562940 498344 562996 499548
rect 555548 497924 555604 497934
rect 555548 497858 555604 497868
rect 564284 497812 564340 497822
rect 564284 497746 564340 497756
rect 558908 457044 558964 457054
rect 558908 456978 558964 456988
rect 555548 453348 555604 456456
rect 555548 453282 555604 453292
rect 556220 453236 556276 456456
rect 556220 453170 556276 453180
rect 559580 444500 559636 456456
rect 561596 451108 561652 456456
rect 562268 453572 562324 456456
rect 562268 453506 562324 453516
rect 562940 453460 562996 456456
rect 562940 453394 562996 453404
rect 561596 451042 561652 451052
rect 559580 444434 559636 444444
rect 536732 444322 536788 444332
rect 533372 437490 533428 437500
rect 561596 430500 561652 430510
rect 494172 430388 494228 430398
rect 494172 427112 494228 430332
rect 503580 430276 503636 430286
rect 500892 428484 500948 428494
rect 500892 427112 500948 428428
rect 503580 427112 503636 430220
rect 560252 428596 560308 428606
rect 560252 427112 560308 428540
rect 561596 427112 561652 430444
rect 474684 427028 474740 427038
rect 474684 380436 474740 426972
rect 556220 427028 556276 427038
rect 556220 426962 556276 426972
rect 493500 426916 493556 426926
rect 493500 426850 493556 426860
rect 500220 426804 500276 426814
rect 500220 426738 500276 426748
rect 497532 426692 497588 426702
rect 497532 426626 497588 426636
rect 557564 426580 557620 426590
rect 557564 426514 557620 426524
rect 502908 426468 502964 426478
rect 502908 426402 502964 426412
rect 535836 408772 535892 408782
rect 495516 385476 495572 385486
rect 495516 385410 495572 385420
rect 499548 385364 499604 385374
rect 474684 380370 474740 380380
rect 493500 374276 493556 385336
rect 493500 374210 493556 374220
rect 498204 373156 498260 385336
rect 498876 384580 498932 385336
rect 499548 385298 499604 385308
rect 498876 384514 498932 384524
rect 498204 373090 498260 373100
rect 498204 358372 498260 358382
rect 493500 358260 493556 358270
rect 475468 357924 475524 357934
rect 475468 353780 475524 357868
rect 493500 355880 493556 358204
rect 494844 357924 494900 357934
rect 494844 355880 494900 357868
rect 497532 356468 497588 356478
rect 495628 356020 495684 356030
rect 495628 355908 495684 355964
rect 495628 355852 496216 355908
rect 497532 355880 497588 356412
rect 498204 355880 498260 358316
rect 500220 357140 500276 357150
rect 500220 355880 500276 357084
rect 500892 356580 500948 356590
rect 500892 355880 500948 356524
rect 501116 355684 501172 355694
rect 501172 355628 501592 355684
rect 501116 355618 501172 355628
rect 499548 355572 499604 355582
rect 499548 355506 499604 355516
rect 475468 353714 475524 353724
rect 535836 341684 535892 408716
rect 535948 387604 536004 387614
rect 535948 382900 536004 387548
rect 537740 387492 537796 387502
rect 537628 387380 537684 387390
rect 537628 383012 537684 387324
rect 537628 382946 537684 382956
rect 535948 382834 536004 382844
rect 537740 382788 537796 387436
rect 537740 382722 537796 382732
rect 553532 382788 553588 385336
rect 554204 382900 554260 385336
rect 558908 383012 558964 385336
rect 559580 384020 559636 385336
rect 559580 383954 559636 383964
rect 558908 382946 558964 382956
rect 554204 382834 554260 382844
rect 553532 382722 553588 382732
rect 560252 378756 560308 385336
rect 560252 378690 560308 378700
rect 558908 358708 558964 358718
rect 539196 358260 539252 358270
rect 539196 353668 539252 358204
rect 557564 358036 557620 358046
rect 557564 355880 557620 357980
rect 558908 355880 558964 358652
rect 566972 358260 567028 358270
rect 562940 358148 562996 358158
rect 562940 355880 562996 358092
rect 566972 355880 567028 358204
rect 539196 353602 539252 353612
rect 535836 341618 535892 341628
rect 561036 314692 561092 314702
rect 561092 314636 561624 314692
rect 561036 314626 561092 314636
rect 500892 314580 500948 314590
rect 500892 314514 500948 314524
rect 493500 314468 493556 314478
rect 493500 314402 493556 314412
rect 562940 314132 562996 314142
rect 496188 313908 496244 314104
rect 496188 313842 496244 313852
rect 496860 311780 496916 314104
rect 499548 313572 499604 314104
rect 499772 314076 500248 314132
rect 499772 314020 499828 314076
rect 499772 313954 499828 313964
rect 499548 313506 499604 313516
rect 553532 312004 553588 314104
rect 553532 311938 553588 311948
rect 554876 311892 554932 314104
rect 557788 314076 558264 314132
rect 558348 314076 558936 314132
rect 557788 312340 557844 314076
rect 558124 313348 558180 313358
rect 558348 313348 558404 314076
rect 558180 313292 558404 313348
rect 558124 313282 558180 313292
rect 557788 312274 557844 312284
rect 554876 311826 554932 311836
rect 496860 311714 496916 311724
rect 560924 311668 560980 314104
rect 562268 312228 562324 314104
rect 562940 314066 562996 314076
rect 562268 312162 562324 312172
rect 560924 311602 560980 311612
rect 474572 311042 474628 311052
rect 433468 308690 433524 308700
rect 430780 306450 430836 306460
rect 376236 304210 376292 304220
rect 373548 303650 373604 303660
rect 372204 301970 372260 301980
rect 400652 298676 400708 298686
rect 351932 288148 351988 288158
rect 347788 239810 347844 239820
rect 348572 215348 348628 215358
rect 340284 215236 340340 215246
rect 340284 206836 340340 215180
rect 345548 213556 345604 213566
rect 342076 212996 342132 213006
rect 340284 206770 340340 206780
rect 341852 212436 341908 212446
rect 340284 205156 340340 205166
rect 340284 169652 340340 205100
rect 341852 186116 341908 212380
rect 342076 204036 342132 212940
rect 342076 203970 342132 203980
rect 345212 199556 345268 199566
rect 341852 186050 341908 186060
rect 341964 191044 342020 191054
rect 340284 169586 340340 169596
rect 340396 182196 340452 182206
rect 340396 160468 340452 182140
rect 341852 178276 341908 178286
rect 341852 162148 341908 178220
rect 341964 169204 342020 190988
rect 345212 171332 345268 199500
rect 345212 171266 345268 171276
rect 345324 192836 345380 192846
rect 345324 169316 345380 192780
rect 345548 191716 345604 213500
rect 348572 200116 348628 215292
rect 348572 200050 348628 200060
rect 345548 191650 345604 191660
rect 349356 198548 349412 268380
rect 350252 287700 350308 287710
rect 350252 249396 350308 287644
rect 350476 287476 350532 287486
rect 350476 259476 350532 287420
rect 350476 259410 350532 259420
rect 350252 249330 350308 249340
rect 350364 253316 350420 253326
rect 349468 245476 349524 245486
rect 349468 241892 349524 245420
rect 349468 241826 349524 241836
rect 350364 241444 350420 253260
rect 351932 242900 351988 288092
rect 376236 287812 376292 287822
rect 352268 286020 352324 286030
rect 352156 284452 352212 284462
rect 351932 242834 351988 242844
rect 352044 271236 352100 271246
rect 350364 241378 350420 241388
rect 352044 241332 352100 271180
rect 352156 269556 352212 284396
rect 352268 270676 352324 285964
rect 375564 286020 375620 286030
rect 368844 285684 368900 285694
rect 368844 284760 368900 285628
rect 375564 284760 375620 285964
rect 376236 284760 376292 287756
rect 376908 284452 376964 284462
rect 376908 284386 376964 284396
rect 352268 270610 352324 270620
rect 352156 269490 352212 269500
rect 352156 252196 352212 252206
rect 352156 243236 352212 252140
rect 374892 243348 374948 243358
rect 374892 243282 374948 243292
rect 352156 243170 352212 243180
rect 352044 241266 352100 241276
rect 359548 242116 359604 242126
rect 359548 240212 359604 242060
rect 370188 241892 370244 242872
rect 370188 241826 370244 241836
rect 359548 240146 359604 240156
rect 372876 240212 372932 242872
rect 375564 241332 375620 242872
rect 400652 241892 400708 298620
rect 563724 296996 563780 297006
rect 504812 296548 504868 296558
rect 499772 294868 499828 294878
rect 499772 288148 499828 294812
rect 504812 288260 504868 296492
rect 518252 296436 518308 296446
rect 518252 289828 518308 296380
rect 560364 295876 560420 295886
rect 518252 289762 518308 289772
rect 559468 289828 559524 289838
rect 504812 288194 504868 288204
rect 556108 288260 556164 288270
rect 499772 288082 499828 288092
rect 498876 288036 498932 288046
rect 436828 287700 436884 287710
rect 436884 287644 436996 287700
rect 436828 287634 436884 287644
rect 433468 285908 433524 285918
rect 433468 284788 433524 285852
rect 436940 284788 436996 287644
rect 433468 284732 434168 284788
rect 436856 284732 436996 284788
rect 438732 287588 438788 287598
rect 438732 284788 438788 287532
rect 477148 287588 477204 287598
rect 477148 286468 477204 287532
rect 477148 286402 477204 286412
rect 498204 287476 498260 287486
rect 475468 285796 475524 285806
rect 438732 284732 439544 284788
rect 434812 284340 434868 284350
rect 434812 284274 434868 284284
rect 432796 284228 432852 284238
rect 432796 284162 432852 284172
rect 475468 283556 475524 285740
rect 498204 284760 498260 287420
rect 498876 284760 498932 287980
rect 501564 287588 501620 287598
rect 500220 286356 500276 286366
rect 499548 285684 499604 285694
rect 499548 284760 499604 285628
rect 500220 284760 500276 286300
rect 500892 285796 500948 285806
rect 500892 284760 500948 285740
rect 501564 284760 501620 287532
rect 554428 287364 554484 287374
rect 554428 284788 554484 287308
rect 556108 284788 556164 288204
rect 559468 284788 559524 289772
rect 560364 284788 560420 295820
rect 554428 284732 554904 284788
rect 556108 284732 556920 284788
rect 559468 284732 559608 284788
rect 560280 284732 560420 284788
rect 561708 288148 561764 288158
rect 561708 284788 561764 288092
rect 563724 284788 563780 296940
rect 561708 284732 562296 284788
rect 563640 284732 563780 284788
rect 475468 283490 475524 283500
rect 438844 243236 438900 243246
rect 438844 243170 438900 243180
rect 436828 243124 436884 243134
rect 436828 243058 436884 243068
rect 448924 243012 448980 243022
rect 448924 242946 448980 242956
rect 493500 242900 493556 242910
rect 400652 241826 400708 241836
rect 432124 241668 432180 242872
rect 432124 241602 432180 241612
rect 434812 241444 434868 242872
rect 493500 242834 493556 242844
rect 494172 241780 494228 242872
rect 494172 241714 494228 241724
rect 434812 241378 434868 241388
rect 375564 241266 375620 241276
rect 372876 240146 372932 240156
rect 496188 239764 496244 242872
rect 496188 239698 496244 239708
rect 503132 240436 503188 240446
rect 350252 233156 350308 233166
rect 350252 222628 350308 233100
rect 437612 232596 437668 232606
rect 427532 224756 427588 224766
rect 414092 224196 414148 224206
rect 350252 222562 350308 222572
rect 406588 223076 406644 223086
rect 398972 220276 399028 220286
rect 372876 216916 372932 216926
rect 352156 215460 352212 215470
rect 350364 215124 350420 215134
rect 345324 169250 345380 169260
rect 348572 181636 348628 181646
rect 341964 169138 342020 169148
rect 341852 162082 341908 162092
rect 341964 167076 342020 167086
rect 340396 160402 340452 160412
rect 341964 158900 342020 167020
rect 341964 158834 342020 158844
rect 340172 152450 340228 152460
rect 340284 153636 340340 153646
rect 339276 152114 339332 152124
rect 338492 151956 338548 151966
rect 338492 101780 338548 151900
rect 338604 144564 338660 144574
rect 338604 136836 338660 144508
rect 338604 136770 338660 136780
rect 338492 101714 338548 101724
rect 340172 112868 340228 112878
rect 336924 100930 336980 100940
rect 338604 100436 338660 100446
rect 338492 94276 338548 94286
rect 336812 26786 336868 26796
rect 337036 69636 337092 69646
rect 337036 26516 337092 69580
rect 338492 29428 338548 94220
rect 338604 90020 338660 100380
rect 338604 89954 338660 89964
rect 338716 93156 338772 93166
rect 338716 29652 338772 93100
rect 338716 29586 338772 29596
rect 338492 29362 338548 29372
rect 340172 26740 340228 112812
rect 340284 101892 340340 153580
rect 340284 101826 340340 101836
rect 340396 143556 340452 143566
rect 340396 98868 340452 143500
rect 342076 142884 342132 142894
rect 341964 130676 342020 130686
rect 340396 98802 340452 98812
rect 340508 111076 340564 111086
rect 340508 94948 340564 111020
rect 340508 94882 340564 94892
rect 341852 108276 341908 108286
rect 341852 29316 341908 108220
rect 341964 100660 342020 130620
rect 342076 128996 342132 142828
rect 342076 128930 342132 128940
rect 345212 142212 345268 142222
rect 345212 125076 345268 142156
rect 345212 125010 345268 125020
rect 345324 123956 345380 123966
rect 342188 117796 342244 117806
rect 341964 100594 342020 100604
rect 342076 114996 342132 115006
rect 342076 86548 342132 114940
rect 342188 96740 342244 117740
rect 345212 115556 345268 115566
rect 343532 110068 343588 110078
rect 343532 98756 343588 110012
rect 343532 98690 343588 98700
rect 342188 96674 342244 96684
rect 342076 86482 342132 86492
rect 341852 29250 341908 29260
rect 345212 28532 345268 115500
rect 345324 93268 345380 123900
rect 346892 113428 346948 113438
rect 346892 98644 346948 113372
rect 348572 98980 348628 181580
rect 348684 144788 348740 144798
rect 348684 136276 348740 144732
rect 348684 136210 348740 136220
rect 349356 127988 349412 198492
rect 350252 212548 350308 212558
rect 350252 183876 350308 212492
rect 350364 188916 350420 215068
rect 351932 213780 351988 213790
rect 350476 213444 350532 213454
rect 350476 196756 350532 213388
rect 350476 196690 350532 196700
rect 351932 196588 351988 213724
rect 350364 188850 350420 188860
rect 351820 196532 351988 196588
rect 352044 213332 352100 213342
rect 350252 183810 350308 183820
rect 350588 187236 350644 187246
rect 348572 98914 348628 98924
rect 348684 119476 348740 119486
rect 346892 98578 346948 98588
rect 345324 93202 345380 93212
rect 348684 78148 348740 119420
rect 348684 78082 348740 78092
rect 348572 74228 348628 74238
rect 348572 66836 348628 74172
rect 348572 66770 348628 66780
rect 345212 28466 345268 28476
rect 348572 59668 348628 59678
rect 340172 26674 340228 26684
rect 337036 26450 337092 26460
rect 348572 26404 348628 59612
rect 349356 57092 349412 127932
rect 350252 180516 350308 180526
rect 350252 99092 350308 180460
rect 350588 171668 350644 187180
rect 351820 184996 351876 196532
rect 351932 195412 351988 195422
rect 352044 195412 352100 213276
rect 352156 201236 352212 215404
rect 368172 215124 368228 215134
rect 366716 213668 366772 213678
rect 366716 213556 366772 213612
rect 366716 213500 367528 213556
rect 368172 213528 368228 215068
rect 372876 213528 372932 216860
rect 376236 213780 376292 213790
rect 376236 213528 376292 213724
rect 370860 212884 370916 212894
rect 370860 212818 370916 212828
rect 378252 212884 378308 212894
rect 378252 212818 378308 212828
rect 352156 201170 352212 201180
rect 351988 195356 352100 195412
rect 351932 195346 351988 195356
rect 351820 184930 351876 184940
rect 352044 187796 352100 187806
rect 350588 171602 350644 171612
rect 351932 178836 351988 178846
rect 351932 152068 351988 178780
rect 352044 169092 352100 187740
rect 352156 182756 352212 182766
rect 352156 171780 352212 182700
rect 393932 174020 393988 174030
rect 352156 171714 352212 171724
rect 368844 171780 368900 171790
rect 368844 171714 368900 171724
rect 375564 171668 375620 171678
rect 373548 169428 373604 171640
rect 375564 171602 375620 171612
rect 376908 171220 376964 171640
rect 376908 171154 376964 171164
rect 373548 169362 373604 169372
rect 352044 169026 352100 169036
rect 377580 169092 377636 171640
rect 393932 169428 393988 173964
rect 398972 171220 399028 220220
rect 406588 219380 406644 223020
rect 406588 219314 406644 219324
rect 398972 171154 399028 171164
rect 412412 218596 412468 218606
rect 412412 171108 412468 218540
rect 414092 171668 414148 224140
rect 427532 218148 427588 224700
rect 427532 218082 427588 218092
rect 429212 221956 429268 221966
rect 429212 217812 429268 221900
rect 434140 219380 434196 219390
rect 429212 217746 429268 217756
rect 433468 218148 433524 218158
rect 430780 213556 430836 213566
rect 433468 213528 433524 218092
rect 434140 213528 434196 219324
rect 437612 217700 437668 232540
rect 473116 230916 473172 230926
rect 440972 230356 441028 230366
rect 437612 217634 437668 217644
rect 439516 217812 439572 217822
rect 436156 217476 436212 217486
rect 436156 213528 436212 217420
rect 437500 215572 437556 215582
rect 437500 213528 437556 215516
rect 439516 213528 439572 217756
rect 440972 217812 441028 230300
rect 464492 226436 464548 226446
rect 440972 217746 441028 217756
rect 461132 225876 461188 225886
rect 430780 213490 430836 213500
rect 436828 213332 436884 213342
rect 436828 213266 436884 213276
rect 414092 171602 414148 171612
rect 432124 171668 432180 171678
rect 432124 171602 432180 171612
rect 432348 171612 432824 171668
rect 438508 171612 438872 171668
rect 439068 171612 439544 171668
rect 440216 171612 440356 171668
rect 412412 171042 412468 171052
rect 393932 169362 393988 169372
rect 432348 169204 432404 171612
rect 438508 171220 438564 171612
rect 438508 171154 438564 171164
rect 439068 169316 439124 171612
rect 440300 171108 440356 171612
rect 461132 171220 461188 225820
rect 461132 171154 461188 171164
rect 440300 171042 440356 171052
rect 464492 171108 464548 226380
rect 464492 171042 464548 171052
rect 473116 170996 473172 230860
rect 474684 227556 474740 227566
rect 473116 170930 473172 170940
rect 474572 174356 474628 174366
rect 439068 169250 439124 169260
rect 472892 169876 472948 169886
rect 432348 169138 432404 169148
rect 377580 169026 377636 169036
rect 414092 165956 414148 165966
rect 398972 164276 399028 164286
rect 351932 152002 351988 152012
rect 372652 152404 372708 152414
rect 372652 147140 372708 152348
rect 376908 152180 376964 152190
rect 372652 147074 372708 147084
rect 372876 150388 372932 150398
rect 352716 144900 352772 144910
rect 352716 143780 352772 144844
rect 352716 143714 352772 143724
rect 350588 143220 350644 143230
rect 350364 137956 350420 137966
rect 350364 100548 350420 137900
rect 350588 126196 350644 143164
rect 369516 143220 369572 143230
rect 351932 143108 351988 143118
rect 351036 141764 351092 141774
rect 351036 138516 351092 141708
rect 351036 138450 351092 138460
rect 350588 126130 350644 126140
rect 351932 124516 351988 143052
rect 352156 142996 352212 143006
rect 352044 142324 352100 142334
rect 352044 128660 352100 142268
rect 352156 135716 352212 142940
rect 368172 142324 368228 142334
rect 369516 142296 369572 143164
rect 372204 142884 372260 142894
rect 372204 142296 372260 142828
rect 372876 142296 372932 150332
rect 374220 147140 374276 147150
rect 373548 143108 373604 143118
rect 373548 142296 373604 143052
rect 374220 142296 374276 147084
rect 376908 142296 376964 152124
rect 393148 142884 393204 142894
rect 368172 142258 368228 142268
rect 375564 142212 375620 142222
rect 375564 142146 375620 142156
rect 376236 142100 376292 142110
rect 376236 142034 376292 142044
rect 393148 139636 393204 142828
rect 393148 139570 393204 139580
rect 352156 135650 352212 135660
rect 352044 128594 352100 128604
rect 351932 124450 351988 124460
rect 352044 114436 352100 114446
rect 350364 100482 350420 100492
rect 350476 107716 350532 107726
rect 350252 99026 350308 99036
rect 350476 96964 350532 107660
rect 350476 96898 350532 96908
rect 351932 102676 351988 102686
rect 349356 57026 349412 57036
rect 350252 96516 350308 96526
rect 350252 29764 350308 96460
rect 350252 29698 350308 29708
rect 351932 29540 351988 102620
rect 352044 88228 352100 114380
rect 352044 88162 352100 88172
rect 352492 107156 352548 107166
rect 351932 29474 351988 29484
rect 352044 78596 352100 78606
rect 352044 26628 352100 78540
rect 352492 78484 352548 107100
rect 398972 101780 399028 164220
rect 410732 163716 410788 163726
rect 398972 101714 399028 101724
rect 407372 160916 407428 160926
rect 407372 100884 407428 160860
rect 407372 100818 407428 100828
rect 368172 100772 368228 100782
rect 368172 100706 368228 100716
rect 368844 100772 368900 100782
rect 368844 100706 368900 100716
rect 376908 100660 376964 100670
rect 376908 100594 376964 100604
rect 410732 100660 410788 163660
rect 412412 161476 412468 161486
rect 410844 159236 410900 159246
rect 410844 102004 410900 159180
rect 410844 101938 410900 101948
rect 412412 101892 412468 161420
rect 413980 145012 414036 145022
rect 413980 140756 414036 144956
rect 413980 140690 414036 140700
rect 412412 101826 412468 101836
rect 414092 101668 414148 165900
rect 414092 101602 414148 101612
rect 414204 159796 414260 159806
rect 410732 100594 410788 100604
rect 414204 100324 414260 159740
rect 437612 147028 437668 147038
rect 437612 145348 437668 146972
rect 437612 145282 437668 145292
rect 435484 145012 435540 145022
rect 434812 144900 434868 144910
rect 432796 144788 432852 144798
rect 432796 142296 432852 144732
rect 434812 142296 434868 144844
rect 435036 143108 435092 143118
rect 435036 142436 435092 143052
rect 435036 142370 435092 142380
rect 435484 142296 435540 144956
rect 437500 144564 437556 144574
rect 437500 142296 437556 144508
rect 438172 142996 438228 143006
rect 438172 142296 438228 142940
rect 444220 100884 444276 100894
rect 444220 100818 444276 100828
rect 472892 100884 472948 169820
rect 472892 100818 472948 100828
rect 422044 100772 422100 100782
rect 422044 100706 422100 100716
rect 429436 100772 429492 100782
rect 429436 100706 429492 100716
rect 434140 100772 434196 100782
rect 434140 100706 434196 100716
rect 438844 100772 438900 100782
rect 438844 100706 438900 100716
rect 435484 100660 435540 100670
rect 435484 100594 435540 100604
rect 474572 100660 474628 174300
rect 474684 170884 474740 227500
rect 501564 217812 501620 217822
rect 500892 217700 500948 217710
rect 475468 215572 475524 215582
rect 475468 211092 475524 215516
rect 496860 215572 496916 215582
rect 495516 215460 495572 215470
rect 492156 215348 492212 215358
rect 492156 213528 492212 215292
rect 495516 213528 495572 215404
rect 496860 213528 496916 215516
rect 500892 213528 500948 217644
rect 501564 213528 501620 217756
rect 503132 217588 503188 240380
rect 553532 239876 553588 242872
rect 555548 240100 555604 242872
rect 555548 240034 555604 240044
rect 553532 239810 553588 239820
rect 557564 239652 557620 242872
rect 560252 239988 560308 242872
rect 562268 241892 562324 242872
rect 562268 241826 562324 241836
rect 560252 239922 560308 239932
rect 557564 239586 557620 239596
rect 536732 236068 536788 236078
rect 503132 217522 503188 217532
rect 523292 234836 523348 234846
rect 496188 213444 496244 213454
rect 496188 213378 496244 213388
rect 475468 211026 475524 211036
rect 493500 171332 493556 171640
rect 493500 171266 493556 171276
rect 494172 170996 494228 171640
rect 494172 170930 494228 170940
rect 474684 170818 474740 170828
rect 494844 170884 494900 171640
rect 495516 171108 495572 171640
rect 496188 171220 496244 171640
rect 523292 171332 523348 234780
rect 533484 232708 533540 232718
rect 523292 171266 523348 171276
rect 533372 172228 533428 172238
rect 496188 171154 496244 171164
rect 495516 171042 495572 171052
rect 494844 170818 494900 170828
rect 493500 167188 493556 167198
rect 475468 144564 475524 144574
rect 475468 140532 475524 144508
rect 493500 142296 493556 167132
rect 494172 158900 494228 158910
rect 494172 142296 494228 158844
rect 497532 144564 497588 144574
rect 497532 142296 497588 144508
rect 500892 143108 500948 143118
rect 498204 142884 498260 142894
rect 498204 142296 498260 142828
rect 500892 142296 500948 143052
rect 492828 141764 492884 141774
rect 492828 141698 492884 141708
rect 475468 140466 475524 140476
rect 498876 100996 498932 101006
rect 498876 100930 498932 100940
rect 499548 100884 499604 100894
rect 499548 100818 499604 100828
rect 474572 100594 474628 100604
rect 495516 100660 495572 100670
rect 495516 100594 495572 100604
rect 420028 100548 420084 100558
rect 420476 100548 420532 100558
rect 420084 100492 420476 100548
rect 500892 100548 500948 100558
rect 420028 100482 420084 100492
rect 420476 100482 420532 100492
rect 414204 100258 414260 100268
rect 428764 100324 428820 100520
rect 428764 100258 428820 100268
rect 430108 98644 430164 100520
rect 492828 98868 492884 100520
rect 492828 98802 492884 98812
rect 494172 98756 494228 100520
rect 500892 100482 500948 100492
rect 533372 98868 533428 172172
rect 533484 169316 533540 232652
rect 533484 169250 533540 169260
rect 536732 169204 536788 236012
rect 560364 235956 560420 235966
rect 560252 227668 560308 227678
rect 555548 217588 555604 217598
rect 539196 215348 539252 215358
rect 539196 210868 539252 215292
rect 555548 213528 555604 217532
rect 558908 215348 558964 215358
rect 558908 213528 558964 215292
rect 560252 213528 560308 227612
rect 560364 216692 560420 235900
rect 564284 222628 564340 222638
rect 560364 216626 560420 216636
rect 562268 216692 562324 216702
rect 562268 213528 562324 216636
rect 562940 215684 562996 215694
rect 562940 213528 562996 215628
rect 563612 215236 563668 215246
rect 563612 213528 563668 215180
rect 564284 213528 564340 222572
rect 557564 212996 557620 213006
rect 557564 212930 557620 212940
rect 539196 210802 539252 210812
rect 580412 192164 580468 569772
rect 580636 403620 580692 570556
rect 580636 403554 580692 403564
rect 582092 569940 582148 569950
rect 582092 271460 582148 569884
rect 587132 569268 587188 569278
rect 582204 567476 582260 567486
rect 582204 548996 582260 567420
rect 582204 548930 582260 548940
rect 585452 567364 585508 567374
rect 585452 469924 585508 567308
rect 585452 469858 585508 469868
rect 582092 271394 582148 271404
rect 580412 192098 580468 192108
rect 536732 169138 536788 169148
rect 554876 171612 555576 171668
rect 556108 171612 556248 171668
rect 558236 171612 558936 171668
rect 559580 171612 560280 171668
rect 562828 171612 562968 171668
rect 571676 171612 572376 171668
rect 554876 169204 554932 171612
rect 556108 169540 556164 171612
rect 556108 169474 556164 169484
rect 558236 169316 558292 171612
rect 559580 169428 559636 171612
rect 562828 169652 562884 171612
rect 571676 171332 571732 171612
rect 571676 171266 571732 171276
rect 562828 169586 562884 169596
rect 559580 169362 559636 169372
rect 558236 169250 558292 169260
rect 554876 169138 554932 169148
rect 556892 162148 556948 162158
rect 556220 152068 556276 152078
rect 536732 150836 536788 150846
rect 536732 101108 536788 150780
rect 556220 142296 556276 152012
rect 556892 142296 556948 162092
rect 557564 160468 557620 160478
rect 557564 142296 557620 160412
rect 561596 145796 561652 145806
rect 560252 145348 560308 145358
rect 560252 142296 560308 145292
rect 561596 142296 561652 145740
rect 587132 113092 587188 569212
rect 587244 567028 587300 567038
rect 587244 324548 587300 566972
rect 590492 350980 590548 570668
rect 590604 569380 590660 569390
rect 590604 535892 590660 569324
rect 590604 535826 590660 535836
rect 590716 528164 590772 528174
rect 590604 521668 590660 521678
rect 590604 390628 590660 521612
rect 590716 496356 590772 528108
rect 590716 496290 590772 496300
rect 590604 390562 590660 390572
rect 590492 350914 590548 350924
rect 587244 324482 587300 324492
rect 587132 113026 587188 113036
rect 536732 101042 536788 101052
rect 556892 101108 556948 101118
rect 556892 101042 556948 101052
rect 533372 98802 533428 98812
rect 556220 98868 556276 100520
rect 558908 98980 558964 100520
rect 564284 99092 564340 100520
rect 564284 99026 564340 99036
rect 558908 98914 558964 98924
rect 556220 98802 556276 98812
rect 494172 98690 494228 98700
rect 430108 98578 430164 98588
rect 438172 96964 438228 96974
rect 355292 94836 355348 94846
rect 355292 80052 355348 94780
rect 355292 79986 355348 79996
rect 372204 90020 372260 90030
rect 352492 78418 352548 78428
rect 371308 78372 371364 78382
rect 371308 75124 371364 78316
rect 371308 75058 371364 75068
rect 352716 74116 352772 74126
rect 352268 70644 352324 70654
rect 352268 66948 352324 70588
rect 352716 68516 352772 74060
rect 359548 74004 359604 74014
rect 359548 70756 359604 73948
rect 368844 74004 368900 74014
rect 368844 71064 368900 73948
rect 372204 71064 372260 89964
rect 432572 89236 432628 89246
rect 403228 87556 403284 87566
rect 393932 85876 393988 85886
rect 375452 84756 375508 84766
rect 375452 74900 375508 84700
rect 375452 74834 375508 74844
rect 379596 80052 379652 80062
rect 376908 74228 376964 74238
rect 372876 74116 372932 74126
rect 372876 71064 372932 74060
rect 376908 71064 376964 74172
rect 379596 71064 379652 79996
rect 393932 75012 393988 85820
rect 403228 81508 403284 87500
rect 403228 81442 403284 81452
rect 407372 81956 407428 81966
rect 404796 80836 404852 80846
rect 404796 78372 404852 80780
rect 404796 78306 404852 78316
rect 404012 78036 404068 78046
rect 393932 74946 393988 74956
rect 402332 76356 402388 76366
rect 402332 74788 402388 76300
rect 402332 74722 402388 74732
rect 359548 70690 359604 70700
rect 371196 70756 371252 70766
rect 371196 70642 371252 70700
rect 371196 70590 371198 70642
rect 371250 70590 371252 70642
rect 371196 70578 371252 70590
rect 373548 70644 373604 70654
rect 377580 70644 377636 70654
rect 373548 70642 374248 70644
rect 373548 70590 373550 70642
rect 373602 70590 374248 70642
rect 373548 70588 374248 70590
rect 373548 70578 373604 70588
rect 377580 70578 377636 70588
rect 352716 68450 352772 68460
rect 352268 66882 352324 66892
rect 372204 29764 372260 29774
rect 372204 29698 372260 29708
rect 370860 29652 370916 29662
rect 370860 29586 370916 29596
rect 404012 29652 404068 77980
rect 404012 29586 404068 29596
rect 377580 29428 377636 29438
rect 377580 29362 377636 29372
rect 407372 29428 407428 81900
rect 432124 74788 432180 74798
rect 432124 71064 432180 74732
rect 432572 74788 432628 89180
rect 436156 78484 436212 78494
rect 432572 74722 432628 74732
rect 433468 75124 433524 75134
rect 433468 71064 433524 75068
rect 436156 71064 436212 78428
rect 438172 71064 438228 96908
rect 556892 96740 556948 96750
rect 504252 94948 504308 94958
rect 461916 91476 461972 91486
rect 461916 84980 461972 91420
rect 461916 84914 461972 84924
rect 464492 90356 464548 90366
rect 461132 83636 461188 83646
rect 407372 29362 407428 29372
rect 414092 31108 414148 31118
rect 352044 26562 352100 26572
rect 348572 26338 348628 26348
rect 374892 26404 374948 29288
rect 376908 26516 376964 29288
rect 376908 26450 376964 26460
rect 414092 26516 414148 31052
rect 434812 29652 434868 29662
rect 434812 29586 434868 29596
rect 434140 29540 434196 29550
rect 434140 29474 434196 29484
rect 436828 29316 436884 29326
rect 432796 26628 432852 29288
rect 461132 29316 461188 83580
rect 436828 29250 436884 29260
rect 432796 26562 432852 26572
rect 414092 26450 414148 26460
rect 438844 26516 438900 29288
rect 461132 29250 461188 29260
rect 464492 26628 464548 90300
rect 494844 88228 494900 88238
rect 492156 81396 492212 81406
rect 492156 75684 492212 81340
rect 494172 78372 494228 78382
rect 492156 75628 492324 75684
rect 492268 71092 492324 75628
rect 492268 71036 492856 71092
rect 494172 71064 494228 78316
rect 494844 71064 494900 88172
rect 498204 86548 498260 86558
rect 497532 75012 497588 75022
rect 497532 71064 497588 74956
rect 498204 71064 498260 86492
rect 499772 85316 499828 85326
rect 499772 74676 499828 85260
rect 501564 74900 501620 74910
rect 499772 74610 499828 74620
rect 500892 74676 500948 74686
rect 500892 71064 500948 74620
rect 501564 71064 501620 74844
rect 504252 71064 504308 94892
rect 554204 93268 554260 93278
rect 554204 71064 554260 93212
rect 556892 71064 556948 96684
rect 560252 84980 560308 84990
rect 557564 78148 557620 78158
rect 557564 71064 557620 78092
rect 560252 71064 560308 84924
rect 560924 81508 560980 81518
rect 560924 71064 560980 81452
rect 562268 74788 562324 74798
rect 562268 71064 562324 74732
rect 498204 29428 498260 29438
rect 498204 29362 498260 29372
rect 499548 29316 499604 29326
rect 492156 26740 492212 29288
rect 494172 26852 494228 29288
rect 495516 28532 495572 29288
rect 499548 29250 499604 29260
rect 495516 28466 495572 28476
rect 494172 26786 494228 26796
rect 492156 26674 492212 26684
rect 464492 26562 464548 26572
rect 562268 26628 562324 29288
rect 562268 26562 562324 26572
rect 438844 26450 438900 26460
rect 374892 26338 374948 26348
rect 329644 24322 329700 24332
rect 4172 22866 4228 22876
rect 11564 5124 11620 5134
rect 11564 480 11620 5068
rect 11368 392 11620 480
rect 11368 -960 11592 392
rect 13272 -960 13496 480
rect 15176 -960 15400 480
rect 17080 -960 17304 480
rect 18984 -960 19208 480
rect 20888 -960 21112 480
rect 22792 -960 23016 480
rect 24696 -960 24920 480
rect 26600 -960 26824 480
rect 28504 -960 28728 480
rect 30408 -960 30632 480
rect 32312 -960 32536 480
rect 34216 -960 34440 480
rect 36120 -960 36344 480
rect 38024 -960 38248 480
rect 39928 -960 40152 480
rect 41832 -960 42056 480
rect 43736 -960 43960 480
rect 45640 -960 45864 480
rect 47544 -960 47768 480
rect 49448 -960 49672 480
rect 51352 -960 51576 480
rect 53256 -960 53480 480
rect 55160 -960 55384 480
rect 57064 -960 57288 480
rect 58968 -960 59192 480
rect 60872 -960 61096 480
rect 62776 -960 63000 480
rect 64680 -960 64904 480
rect 66584 -960 66808 480
rect 68488 -960 68712 480
rect 70392 -960 70616 480
rect 72296 -960 72520 480
rect 74200 -960 74424 480
rect 76104 -960 76328 480
rect 78008 -960 78232 480
rect 79912 -960 80136 480
rect 81816 -960 82040 480
rect 83720 -960 83944 480
rect 85624 -960 85848 480
rect 87528 -960 87752 480
rect 89432 -960 89656 480
rect 91336 -960 91560 480
rect 93240 -960 93464 480
rect 95144 -960 95368 480
rect 97048 -960 97272 480
rect 98952 -960 99176 480
rect 100856 -960 101080 480
rect 102760 -960 102984 480
rect 104664 -960 104888 480
rect 106568 -960 106792 480
rect 108472 -960 108696 480
rect 110376 -960 110600 480
rect 112280 -960 112504 480
rect 114184 -960 114408 480
rect 116088 -960 116312 480
rect 117992 -960 118216 480
rect 119896 -960 120120 480
rect 121800 -960 122024 480
rect 123704 -960 123928 480
rect 125608 -960 125832 480
rect 127512 -960 127736 480
rect 129416 -960 129640 480
rect 131320 -960 131544 480
rect 133224 -960 133448 480
rect 135128 -960 135352 480
rect 137032 -960 137256 480
rect 138936 -960 139160 480
rect 140840 -960 141064 480
rect 142744 -960 142968 480
rect 144648 -960 144872 480
rect 146552 -960 146776 480
rect 148456 -960 148680 480
rect 150360 -960 150584 480
rect 152264 -960 152488 480
rect 154168 -960 154392 480
rect 156072 -960 156296 480
rect 157976 -960 158200 480
rect 159880 -960 160104 480
rect 161784 -960 162008 480
rect 163688 -960 163912 480
rect 165592 -960 165816 480
rect 167496 -960 167720 480
rect 169400 -960 169624 480
rect 171304 -960 171528 480
rect 173208 -960 173432 480
rect 175112 -960 175336 480
rect 177016 -960 177240 480
rect 178920 -960 179144 480
rect 180824 -960 181048 480
rect 182728 -960 182952 480
rect 184632 -960 184856 480
rect 186536 -960 186760 480
rect 188440 -960 188664 480
rect 190344 -960 190568 480
rect 192248 -960 192472 480
rect 194152 -960 194376 480
rect 196056 -960 196280 480
rect 197960 -960 198184 480
rect 199864 -960 200088 480
rect 201768 -960 201992 480
rect 203672 -960 203896 480
rect 205576 -960 205800 480
rect 207480 -960 207704 480
rect 209384 -960 209608 480
rect 211288 -960 211512 480
rect 213192 -960 213416 480
rect 215096 -960 215320 480
rect 217000 -960 217224 480
rect 218904 -960 219128 480
rect 220808 -960 221032 480
rect 222712 -960 222936 480
rect 224616 -960 224840 480
rect 226520 -960 226744 480
rect 228424 -960 228648 480
rect 230328 -960 230552 480
rect 232232 -960 232456 480
rect 234136 -960 234360 480
rect 236040 -960 236264 480
rect 237944 -960 238168 480
rect 239848 -960 240072 480
rect 241752 -960 241976 480
rect 243656 -960 243880 480
rect 245560 -960 245784 480
rect 247464 -960 247688 480
rect 249368 -960 249592 480
rect 251272 -960 251496 480
rect 253176 -960 253400 480
rect 255080 -960 255304 480
rect 256984 -960 257208 480
rect 258888 -960 259112 480
rect 260792 -960 261016 480
rect 262696 -960 262920 480
rect 264600 -960 264824 480
rect 266504 -960 266728 480
rect 268408 -960 268632 480
rect 270312 -960 270536 480
rect 272216 -960 272440 480
rect 274120 -960 274344 480
rect 276024 -960 276248 480
rect 277928 -960 278152 480
rect 279832 -960 280056 480
rect 281736 -960 281960 480
rect 283640 -960 283864 480
rect 285544 -960 285768 480
rect 287448 -960 287672 480
rect 289352 -960 289576 480
rect 291256 -960 291480 480
rect 293160 -960 293384 480
rect 295064 -960 295288 480
rect 296968 -960 297192 480
rect 298872 -960 299096 480
rect 300776 -960 301000 480
rect 302680 -960 302904 480
rect 304584 -960 304808 480
rect 306488 -960 306712 480
rect 308392 -960 308616 480
rect 310296 -960 310520 480
rect 312200 -960 312424 480
rect 314104 -960 314328 480
rect 316008 -960 316232 480
rect 317912 -960 318136 480
rect 319816 -960 320040 480
rect 321720 -960 321944 480
rect 323624 -960 323848 480
rect 325528 -960 325752 480
rect 327432 -960 327656 480
rect 329336 -960 329560 480
rect 331240 -960 331464 480
rect 333144 -960 333368 480
rect 335048 -960 335272 480
rect 336952 -960 337176 480
rect 338856 -960 339080 480
rect 340760 -960 340984 480
rect 342664 -960 342888 480
rect 344568 -960 344792 480
rect 346472 -960 346696 480
rect 348376 -960 348600 480
rect 350280 -960 350504 480
rect 352184 -960 352408 480
rect 354088 -960 354312 480
rect 355992 -960 356216 480
rect 357896 -960 358120 480
rect 359800 -960 360024 480
rect 361704 -960 361928 480
rect 363608 -960 363832 480
rect 365512 -960 365736 480
rect 367416 -960 367640 480
rect 369320 -960 369544 480
rect 371224 -960 371448 480
rect 373128 -960 373352 480
rect 375032 -960 375256 480
rect 376936 -960 377160 480
rect 378840 -960 379064 480
rect 380744 -960 380968 480
rect 382648 -960 382872 480
rect 384552 -960 384776 480
rect 386456 -960 386680 480
rect 388360 -960 388584 480
rect 390264 -960 390488 480
rect 392168 -960 392392 480
rect 394072 -960 394296 480
rect 395976 -960 396200 480
rect 397880 -960 398104 480
rect 399784 -960 400008 480
rect 401688 -960 401912 480
rect 403592 -960 403816 480
rect 405496 -960 405720 480
rect 407400 -960 407624 480
rect 409304 -960 409528 480
rect 411208 -960 411432 480
rect 413112 -960 413336 480
rect 415016 -960 415240 480
rect 416920 -960 417144 480
rect 418824 -960 419048 480
rect 420728 -960 420952 480
rect 422632 -960 422856 480
rect 424536 -960 424760 480
rect 426440 -960 426664 480
rect 428344 -960 428568 480
rect 430248 -960 430472 480
rect 432152 -960 432376 480
rect 434056 -960 434280 480
rect 435960 -960 436184 480
rect 437864 -960 438088 480
rect 439768 -960 439992 480
rect 441672 -960 441896 480
rect 443576 -960 443800 480
rect 445480 -960 445704 480
rect 447384 -960 447608 480
rect 449288 -960 449512 480
rect 451192 -960 451416 480
rect 453096 -960 453320 480
rect 455000 -960 455224 480
rect 456904 -960 457128 480
rect 458808 -960 459032 480
rect 460712 -960 460936 480
rect 462616 -960 462840 480
rect 464520 -960 464744 480
rect 466424 -960 466648 480
rect 468328 -960 468552 480
rect 470232 -960 470456 480
rect 472136 -960 472360 480
rect 474040 -960 474264 480
rect 475944 -960 476168 480
rect 477848 -960 478072 480
rect 479752 -960 479976 480
rect 481656 -960 481880 480
rect 483560 -960 483784 480
rect 485464 -960 485688 480
rect 487368 -960 487592 480
rect 489272 -960 489496 480
rect 491176 -960 491400 480
rect 493080 -960 493304 480
rect 494984 -960 495208 480
rect 496888 -960 497112 480
rect 498792 -960 499016 480
rect 500696 -960 500920 480
rect 502600 -960 502824 480
rect 504504 -960 504728 480
rect 506408 -960 506632 480
rect 508312 -960 508536 480
rect 510216 -960 510440 480
rect 512120 -960 512344 480
rect 514024 -960 514248 480
rect 515928 -960 516152 480
rect 517832 -960 518056 480
rect 519736 -960 519960 480
rect 521640 -960 521864 480
rect 523544 -960 523768 480
rect 525448 -960 525672 480
rect 527352 -960 527576 480
rect 529256 -960 529480 480
rect 531160 -960 531384 480
rect 533064 -960 533288 480
rect 534968 -960 535192 480
rect 536872 -960 537096 480
rect 538776 -960 539000 480
rect 540680 -960 540904 480
rect 542584 -960 542808 480
rect 544488 -960 544712 480
rect 546392 -960 546616 480
rect 548296 -960 548520 480
rect 550200 -960 550424 480
rect 552104 -960 552328 480
rect 554008 -960 554232 480
rect 555912 -960 556136 480
rect 557816 -960 558040 480
rect 559720 -960 559944 480
rect 561624 -960 561848 480
rect 563528 -960 563752 480
rect 565432 -960 565656 480
rect 567336 -960 567560 480
rect 569240 -960 569464 480
rect 571144 -960 571368 480
rect 573048 -960 573272 480
rect 574952 -960 575176 480
rect 576856 -960 577080 480
rect 578760 -960 578984 480
rect 580664 -960 580888 480
rect 582568 -960 582792 480
rect 584472 -960 584696 480
<< via2 >>
rect 33292 590492 33348 590548
rect 46172 590492 46228 590548
rect 46172 583772 46228 583828
rect 11004 578732 11060 578788
rect 99484 590492 99540 590548
rect 165676 590604 165732 590660
rect 209580 582204 209636 582260
rect 231644 577164 231700 577220
rect 284732 590604 284788 590660
rect 279244 582092 279300 582148
rect 275772 574028 275828 574084
rect 278124 575372 278180 575428
rect 143388 573916 143444 573972
rect 77308 573692 77364 573748
rect 76412 573020 76468 573076
rect 40236 571900 40292 571956
rect 38892 571340 38948 571396
rect 4284 570668 4340 570724
rect 4172 567196 4228 567252
rect 4172 559132 4228 559188
rect 4172 523292 4228 523348
rect 36876 569548 36932 569604
rect 44268 571676 44324 571732
rect 41580 571452 41636 571508
rect 40236 570444 40292 570500
rect 62972 571676 63028 571732
rect 45612 571564 45668 571620
rect 46956 571228 47012 571284
rect 46732 569660 46788 569716
rect 4508 569324 4564 569380
rect 4396 567084 4452 567140
rect 15932 569100 15988 569156
rect 4508 474460 4564 474516
rect 7644 568988 7700 569044
rect 7532 403676 7588 403732
rect 4396 262780 4452 262836
rect 4508 296492 4564 296548
rect 4284 220444 4340 220500
rect 4396 234444 4452 234500
rect 4396 177996 4452 178052
rect 4396 149660 4452 149716
rect 4172 51100 4228 51156
rect 4284 107324 4340 107380
rect 4620 191996 4676 192052
rect 4620 150332 4676 150388
rect 4508 135772 4564 135828
rect 4396 91532 4452 91588
rect 4396 64988 4452 65044
rect 4396 52892 4452 52948
rect 4284 31052 4340 31108
rect 7644 347452 7700 347508
rect 12572 530684 12628 530740
rect 7532 29372 7588 29428
rect 10892 52892 10948 52948
rect 12572 29596 12628 29652
rect 14252 488348 14308 488404
rect 18396 554428 18452 554484
rect 36204 524972 36260 525028
rect 38220 511532 38276 511588
rect 40236 523404 40292 523460
rect 40908 518476 40964 518532
rect 69692 571564 69748 571620
rect 63196 571228 63252 571284
rect 63196 528108 63252 528164
rect 62972 506492 63028 506548
rect 73052 571452 73108 571508
rect 73052 506604 73108 506660
rect 69692 505820 69748 505876
rect 39564 503020 39620 503076
rect 36204 500892 36260 500948
rect 62972 500892 63028 500948
rect 40908 500780 40964 500836
rect 36876 500668 36932 500724
rect 37548 498988 37604 499044
rect 46956 499212 47012 499268
rect 43596 497756 43652 497812
rect 18396 483980 18452 484036
rect 40236 452732 40292 452788
rect 38220 439292 38276 439348
rect 62972 445340 63028 445396
rect 74732 500780 74788 500836
rect 44940 439404 44996 439460
rect 74732 437836 74788 437892
rect 42924 437724 42980 437780
rect 38892 430668 38948 430724
rect 38556 427532 38612 427588
rect 39564 430220 39620 430276
rect 69692 430220 69748 430276
rect 42924 428428 42980 428484
rect 40236 426748 40292 426804
rect 44268 426524 44324 426580
rect 15932 389564 15988 389620
rect 18396 411740 18452 411796
rect 18396 409388 18452 409444
rect 69692 385868 69748 385924
rect 73052 426524 73108 426580
rect 42252 380604 42308 380660
rect 42924 380492 42980 380548
rect 73052 360780 73108 360836
rect 45612 358204 45668 358260
rect 36204 358092 36260 358148
rect 35532 357980 35588 358036
rect 38892 357868 38948 357924
rect 40908 356300 40964 356356
rect 44268 356188 44324 356244
rect 62188 358204 62244 358260
rect 61292 358092 61348 358148
rect 34860 355516 34916 355572
rect 40236 355292 40292 355348
rect 62188 353724 62244 353780
rect 62972 357980 63028 358036
rect 61292 353612 61348 353668
rect 18396 341628 18452 341684
rect 14252 29484 14308 29540
rect 15932 319004 15988 319060
rect 38892 305340 38948 305396
rect 44268 314076 44324 314132
rect 56364 313964 56420 314020
rect 43596 302540 43652 302596
rect 62972 301420 63028 301476
rect 74732 357868 74788 357924
rect 36876 300860 36932 300916
rect 74732 300300 74788 300356
rect 45052 288204 45108 288260
rect 40236 287420 40292 287476
rect 41916 285740 41972 285796
rect 41356 285628 41412 285684
rect 37548 284284 37604 284340
rect 42252 284172 42308 284228
rect 18396 270396 18452 270452
rect 18396 198940 18452 198996
rect 18396 197820 18452 197876
rect 18396 127932 18452 127988
rect 18396 56812 18452 56868
rect 19292 276668 19348 276724
rect 26796 240156 26852 240212
rect 38220 241724 38276 241780
rect 37548 240044 37604 240100
rect 44268 241836 44324 241892
rect 48636 241052 48692 241108
rect 48636 240156 48692 240212
rect 46284 239932 46340 239988
rect 42924 239820 42980 239876
rect 40236 239484 40292 239540
rect 41580 215964 41636 216020
rect 40908 215404 40964 215460
rect 35532 215292 35588 215348
rect 61292 215404 61348 215460
rect 44940 215068 44996 215124
rect 46956 213612 47012 213668
rect 45612 213500 45668 213556
rect 40236 213388 40292 213444
rect 44268 212940 44324 212996
rect 61292 210812 61348 210868
rect 69692 213052 69748 213108
rect 62076 173852 62132 173908
rect 35196 169484 35252 169540
rect 41580 171164 41636 171220
rect 39564 169372 39620 169428
rect 44940 171276 44996 171332
rect 43484 169260 43540 169316
rect 69692 171164 69748 171220
rect 62076 169260 62132 169316
rect 38556 168924 38612 168980
rect 69692 155820 69748 155876
rect 42252 152460 42308 152516
rect 38220 144956 38276 145012
rect 40908 142828 40964 142884
rect 62972 151900 63028 151956
rect 42924 144620 42980 144676
rect 43596 101052 43652 101108
rect 45612 101052 45668 101108
rect 44268 100940 44324 100996
rect 37548 100828 37604 100884
rect 38220 98924 38276 98980
rect 42252 99036 42308 99092
rect 38892 98812 38948 98868
rect 74732 155260 74788 155316
rect 69692 100828 69748 100884
rect 73052 152012 73108 152068
rect 74732 101612 74788 101668
rect 73052 98924 73108 98980
rect 62972 98812 63028 98868
rect 74732 95900 74788 95956
rect 62972 94780 63028 94836
rect 42252 89964 42308 90020
rect 41580 84924 41636 84980
rect 38892 79772 38948 79828
rect 35532 74172 35588 74228
rect 50316 88172 50372 88228
rect 45612 74060 45668 74116
rect 45276 72380 45332 72436
rect 43820 70476 43876 70532
rect 61292 31164 61348 31220
rect 19292 29036 19348 29092
rect 15932 28476 15988 28532
rect 39564 26572 39620 26628
rect 38892 26460 38948 26516
rect 43596 28364 43652 28420
rect 55692 26796 55748 26852
rect 42924 26684 42980 26740
rect 40236 26348 40292 26404
rect 73052 93324 73108 93380
rect 63084 71260 63140 71316
rect 63084 28364 63140 28420
rect 266252 572348 266308 572404
rect 249452 572124 249508 572180
rect 160188 571788 160244 571844
rect 104860 571564 104916 571620
rect 100156 571452 100212 571508
rect 78092 571340 78148 571396
rect 130172 571564 130228 571620
rect 107548 571340 107604 571396
rect 125132 569660 125188 569716
rect 98812 525084 98868 525140
rect 100156 523516 100212 523572
rect 99484 511980 99540 512036
rect 106876 521948 106932 522004
rect 107548 521836 107604 521892
rect 103516 516684 103572 516740
rect 102844 511420 102900 511476
rect 102172 509964 102228 510020
rect 130172 513212 130228 513268
rect 136892 571452 136948 571508
rect 125132 503580 125188 503636
rect 78092 503132 78148 503188
rect 98812 501116 98868 501172
rect 125132 501116 125188 501172
rect 100156 501004 100212 501060
rect 100828 500892 100884 500948
rect 104860 500780 104916 500836
rect 104188 499100 104244 499156
rect 103516 498316 103572 498372
rect 125132 456540 125188 456596
rect 130172 501004 130228 501060
rect 76412 29708 76468 29764
rect 78092 446012 78148 446068
rect 103516 453180 103572 453236
rect 104188 452060 104244 452116
rect 102844 447692 102900 447748
rect 100828 444332 100884 444388
rect 135212 500892 135268 500948
rect 187292 571788 187348 571844
rect 170268 571676 170324 571732
rect 164220 571564 164276 571620
rect 160860 571452 160916 571508
rect 162876 569884 162932 569940
rect 169596 569996 169652 570052
rect 168924 569772 168980 569828
rect 166460 569660 166516 569716
rect 157052 518476 157108 518532
rect 164220 525196 164276 525252
rect 162876 523740 162932 523796
rect 160188 513324 160244 513380
rect 168924 523628 168980 523684
rect 168252 518700 168308 518756
rect 167580 508172 167636 508228
rect 170492 523516 170548 523572
rect 170492 510300 170548 510356
rect 169596 504924 169652 504980
rect 157052 501340 157108 501396
rect 166236 501004 166292 501060
rect 164220 499436 164276 499492
rect 155484 499324 155540 499380
rect 162876 498428 162932 498484
rect 170940 500892 170996 500948
rect 166908 498204 166964 498260
rect 224812 571788 224868 571844
rect 224140 571228 224196 571284
rect 187404 569996 187460 570052
rect 192332 569884 192388 569940
rect 187404 518140 187460 518196
rect 188076 521948 188132 522004
rect 199052 569772 199108 569828
rect 198156 523628 198212 523684
rect 192332 519260 192388 519316
rect 192444 521836 192500 521892
rect 188076 515340 188132 515396
rect 247996 571676 248052 571732
rect 247772 571564 247828 571620
rect 231532 569996 231588 570052
rect 228172 569884 228228 569940
rect 226156 569772 226212 569828
rect 230860 568876 230916 568932
rect 227500 527884 227556 527940
rect 224028 527772 224084 527828
rect 224812 527660 224868 527716
rect 224700 525980 224756 526036
rect 230188 525308 230244 525364
rect 244412 525308 244468 525364
rect 199052 517580 199108 517636
rect 198156 517020 198212 517076
rect 192444 509740 192500 509796
rect 187292 498092 187348 498148
rect 187404 501004 187460 501060
rect 164892 497980 164948 498036
rect 179004 497868 179060 497924
rect 136892 496412 136948 496468
rect 160860 456876 160916 456932
rect 162876 449484 162932 449540
rect 166236 442652 166292 442708
rect 135212 441196 135268 441252
rect 130172 439628 130228 439684
rect 168924 435260 168980 435316
rect 170492 449484 170548 449540
rect 166908 434140 166964 434196
rect 170492 432460 170548 432516
rect 171388 430668 171444 430724
rect 162876 430556 162932 430612
rect 105532 430444 105588 430500
rect 103516 430332 103572 430388
rect 98140 430220 98196 430276
rect 102844 428540 102900 428596
rect 130172 430444 130228 430500
rect 99484 426972 99540 427028
rect 102172 426860 102228 426916
rect 88060 426412 88116 426468
rect 105532 384636 105588 384692
rect 106204 384524 106260 384580
rect 103516 368620 103572 368676
rect 100828 367500 100884 367556
rect 161532 430108 161588 430164
rect 168924 430444 168980 430500
rect 165564 428764 165620 428820
rect 164220 428652 164276 428708
rect 167580 427084 167636 427140
rect 187292 430556 187348 430612
rect 171388 427644 171444 427700
rect 174636 430332 174692 430388
rect 166236 426636 166292 426692
rect 174636 426636 174692 426692
rect 160860 426412 160916 426468
rect 170268 426412 170324 426468
rect 168252 385308 168308 385364
rect 167580 376460 167636 376516
rect 130172 373772 130228 373828
rect 195692 500892 195748 500948
rect 187516 498204 187572 498260
rect 187516 431340 187572 431396
rect 192332 497980 192388 498036
rect 230188 500892 230244 500948
rect 200732 500780 200788 500836
rect 197372 499212 197428 499268
rect 197372 449820 197428 449876
rect 199052 497756 199108 497812
rect 195692 447804 195748 447860
rect 199052 447020 199108 447076
rect 192332 430780 192388 430836
rect 197372 430444 197428 430500
rect 187404 429660 187460 429716
rect 195692 430108 195748 430164
rect 192332 428764 192388 428820
rect 188972 427084 189028 427140
rect 187404 425964 187460 426020
rect 189084 426076 189140 426132
rect 189084 375900 189140 375956
rect 192332 374780 192388 374836
rect 188972 373660 189028 373716
rect 187404 373100 187460 373156
rect 226156 500780 226212 500836
rect 222796 499548 222852 499604
rect 205772 498988 205828 499044
rect 231532 499212 231588 499268
rect 232204 498988 232260 499044
rect 244412 498540 244468 498596
rect 226828 497756 226884 497812
rect 257852 571900 257908 571956
rect 256172 571788 256228 571844
rect 249676 571228 249732 571284
rect 249676 525420 249732 525476
rect 252812 569548 252868 569604
rect 249900 524972 249956 525028
rect 249452 523292 249508 523348
rect 249676 523404 249732 523460
rect 249564 513324 249620 513380
rect 247996 489580 248052 489636
rect 249452 498428 249508 498484
rect 247772 489020 247828 489076
rect 248108 472780 248164 472836
rect 247772 470540 247828 470596
rect 230860 456876 230916 456932
rect 229516 456652 229572 456708
rect 227500 456428 227556 456484
rect 226156 455196 226212 455252
rect 231532 455084 231588 455140
rect 249564 493500 249620 493556
rect 249900 479612 249956 479668
rect 249676 476700 249732 476756
rect 254492 568876 254548 568932
rect 253036 525196 253092 525252
rect 252812 476140 252868 476196
rect 252924 499548 252980 499604
rect 249452 464380 249508 464436
rect 249564 467180 249620 467236
rect 248108 456652 248164 456708
rect 252028 465500 252084 465556
rect 252028 457996 252084 458052
rect 249564 455196 249620 455252
rect 247772 455084 247828 455140
rect 222796 453516 222852 453572
rect 247772 452732 247828 452788
rect 222124 450268 222180 450324
rect 225932 450268 225988 450324
rect 205772 443660 205828 443716
rect 202412 442652 202468 442708
rect 225932 438620 225988 438676
rect 202412 432012 202468 432068
rect 230860 430556 230916 430612
rect 222124 430444 222180 430500
rect 211372 427084 211428 427140
rect 226828 430332 226884 430388
rect 223356 430220 223412 430276
rect 223356 429212 223412 429268
rect 224140 430108 224196 430164
rect 228172 430220 228228 430276
rect 229628 427196 229684 427252
rect 240268 428764 240324 428820
rect 222796 426412 222852 426468
rect 232204 426412 232260 426468
rect 200732 424620 200788 424676
rect 249564 447692 249620 447748
rect 249452 428540 249508 428596
rect 247772 421260 247828 421316
rect 247884 427196 247940 427252
rect 247884 414540 247940 414596
rect 247772 401100 247828 401156
rect 230860 385532 230916 385588
rect 253036 491820 253092 491876
rect 253148 498988 253204 499044
rect 254492 495740 254548 495796
rect 254604 509964 254660 510020
rect 254716 504924 254772 504980
rect 256172 494620 256228 494676
rect 256284 497868 256340 497924
rect 254716 490140 254772 490196
rect 254604 482860 254660 482916
rect 253148 466620 253204 466676
rect 256172 471100 256228 471156
rect 263004 571452 263060 571508
rect 261212 571340 261268 571396
rect 259756 569996 259812 570052
rect 257964 569884 258020 569940
rect 259532 569660 259588 569716
rect 258188 525084 258244 525140
rect 257964 494060 258020 494116
rect 258076 498316 258132 498372
rect 257852 480396 257908 480452
rect 256284 461020 256340 461076
rect 257852 468636 257908 468692
rect 256172 458108 256228 458164
rect 258188 481180 258244 481236
rect 258300 499212 258356 499268
rect 259756 527100 259812 527156
rect 259756 516684 259812 516740
rect 259532 491260 259588 491316
rect 259644 499100 259700 499156
rect 258300 468300 258356 468356
rect 259532 468860 259588 468916
rect 259532 456428 259588 456484
rect 258076 454860 258132 454916
rect 257852 453516 257908 453572
rect 252924 440300 252980 440356
rect 258076 444332 258132 444388
rect 253036 439292 253092 439348
rect 249788 430444 249844 430500
rect 249564 422940 249620 422996
rect 249676 426188 249732 426244
rect 252924 428652 252980 428708
rect 249788 409500 249844 409556
rect 252812 426972 252868 427028
rect 249676 402220 249732 402276
rect 257852 430556 257908 430612
rect 256172 428428 256228 428484
rect 253036 421820 253092 421876
rect 253148 425964 253204 426020
rect 253148 412300 253204 412356
rect 252924 405580 252980 405636
rect 252812 396060 252868 396116
rect 249452 394380 249508 394436
rect 222796 384412 222852 384468
rect 247772 385308 247828 385364
rect 249676 393820 249732 393876
rect 256284 427084 256340 427140
rect 256284 408380 256340 408436
rect 256172 391580 256228 391636
rect 256284 393260 256340 393316
rect 256284 384636 256340 384692
rect 249676 384524 249732 384580
rect 257964 426300 258020 426356
rect 258300 439404 258356 439460
rect 258076 422380 258132 422436
rect 258188 426860 258244 426916
rect 257964 392140 258020 392196
rect 258076 411740 258132 411796
rect 258300 417340 258356 417396
rect 259532 430332 259588 430388
rect 258188 399420 258244 399476
rect 258076 384412 258132 384468
rect 257852 383068 257908 383124
rect 229516 377580 229572 377636
rect 247772 380604 247828 380660
rect 197372 375340 197428 375396
rect 195692 372540 195748 372596
rect 187292 370860 187348 370916
rect 107548 366940 107604 366996
rect 100156 365820 100212 365876
rect 259756 483980 259812 484036
rect 259868 500892 259924 500948
rect 261660 511532 261716 511588
rect 261212 482300 261268 482356
rect 261324 500780 261380 500836
rect 259868 469420 259924 469476
rect 261548 499324 261604 499380
rect 261436 497756 261492 497812
rect 261772 508172 261828 508228
rect 261772 492380 261828 492436
rect 262892 500668 262948 500724
rect 261660 477260 261716 477316
rect 261548 458220 261604 458276
rect 261436 436940 261492 436996
rect 261660 437724 261716 437780
rect 261324 435820 261380 435876
rect 261212 430220 261268 430276
rect 259644 427420 259700 427476
rect 259756 428764 259812 428820
rect 259756 410060 259812 410116
rect 261324 426748 261380 426804
rect 264572 570444 264628 570500
rect 263116 569772 263172 569828
rect 263788 530460 263844 530516
rect 263788 527772 263844 527828
rect 265132 528108 265188 528164
rect 264572 506940 264628 506996
rect 264684 513212 264740 513268
rect 263116 496300 263172 496356
rect 263228 499436 263284 499492
rect 263004 487900 263060 487956
rect 264572 498092 264628 498148
rect 264572 488460 264628 488516
rect 264684 480620 264740 480676
rect 264796 506604 264852 506660
rect 263900 480396 263956 480452
rect 263788 479612 263844 479668
rect 263788 478380 263844 478436
rect 263900 474460 263956 474516
rect 265020 506492 265076 506548
rect 264908 503132 264964 503188
rect 265132 500780 265188 500836
rect 265132 496412 265188 496468
rect 265132 485660 265188 485716
rect 265020 480060 265076 480116
rect 264908 475580 264964 475636
rect 264796 473900 264852 473956
rect 263788 472220 263844 472276
rect 263788 468636 263844 468692
rect 263228 459340 263284 459396
rect 264572 447804 264628 447860
rect 265132 441196 265188 441252
rect 264572 430220 264628 430276
rect 265020 437836 265076 437892
rect 262892 417900 262948 417956
rect 263004 430108 263060 430164
rect 261660 416780 261716 416836
rect 261324 388780 261380 388836
rect 261436 411180 261492 411236
rect 261436 385532 261492 385588
rect 264684 429212 264740 429268
rect 264572 427644 264628 427700
rect 263116 426076 263172 426132
rect 263116 407820 263172 407876
rect 264684 398860 264740 398916
rect 264796 427532 264852 427588
rect 264572 389340 264628 389396
rect 264908 426636 264964 426692
rect 265356 439628 265412 439684
rect 265356 427980 265412 428036
rect 265132 426860 265188 426916
rect 265020 415660 265076 415716
rect 264908 397180 264964 397236
rect 264796 388220 264852 388276
rect 263004 380940 263060 380996
rect 263788 383068 263844 383124
rect 261212 379820 261268 379876
rect 261436 380492 261492 380548
rect 259532 379260 259588 379316
rect 247772 359100 247828 359156
rect 229516 358316 229572 358372
rect 158844 358204 158900 358260
rect 97468 358092 97524 358148
rect 81452 356300 81508 356356
rect 122668 358092 122724 358148
rect 100828 357980 100884 358036
rect 99484 356300 99540 356356
rect 104188 357868 104244 357924
rect 108220 356412 108276 356468
rect 107548 355628 107604 355684
rect 104860 355404 104916 355460
rect 122668 353836 122724 353892
rect 138572 357980 138628 358036
rect 100156 313852 100212 313908
rect 104860 311612 104916 311668
rect 104188 308700 104244 308756
rect 101500 307020 101556 307076
rect 99484 306460 99540 306516
rect 158172 356524 158228 356580
rect 186396 358204 186452 358260
rect 163548 358092 163604 358148
rect 166236 357980 166292 358036
rect 166908 356636 166964 356692
rect 168924 355852 168980 355908
rect 161532 355740 161588 355796
rect 225484 358204 225540 358260
rect 199052 358092 199108 358148
rect 186396 353948 186452 354004
rect 187292 356636 187348 356692
rect 187292 315420 187348 315476
rect 187516 355740 187572 355796
rect 166236 314636 166292 314692
rect 163548 314524 163604 314580
rect 187516 314188 187572 314244
rect 160188 313740 160244 313796
rect 167580 312396 167636 312452
rect 164220 312284 164276 312340
rect 224812 358092 224868 358148
rect 223356 355964 223412 356020
rect 228172 356636 228228 356692
rect 249452 358316 249508 358372
rect 248556 358204 248612 358260
rect 247996 357980 248052 358036
rect 247772 356524 247828 356580
rect 232204 356076 232260 356132
rect 248332 355852 248388 355908
rect 248556 349580 248612 349636
rect 248332 349020 248388 349076
rect 247996 348572 248052 348628
rect 247772 344540 247828 344596
rect 247772 319900 247828 319956
rect 225484 314412 225540 314468
rect 199052 313180 199108 313236
rect 168924 312172 168980 312228
rect 221452 311948 221508 312004
rect 224140 311836 224196 311892
rect 257964 358092 258020 358148
rect 252924 356300 252980 356356
rect 249564 356076 249620 356132
rect 252812 355964 252868 356020
rect 249788 355628 249844 355684
rect 249788 336140 249844 336196
rect 249564 324380 249620 324436
rect 256284 355292 256340 355348
rect 252924 337260 252980 337316
rect 256172 340060 256228 340116
rect 252812 321020 252868 321076
rect 249452 319340 249508 319396
rect 249452 318780 249508 318836
rect 247996 318220 248052 318276
rect 248556 317660 248612 317716
rect 248556 314524 248612 314580
rect 256284 329980 256340 330036
rect 257852 346780 257908 346836
rect 256172 313852 256228 313908
rect 249452 313740 249508 313796
rect 263788 378140 263844 378196
rect 263788 373772 263844 373828
rect 263788 369740 263844 369796
rect 261436 357980 261492 358036
rect 261660 357868 261716 357924
rect 258076 356412 258132 356468
rect 258076 334460 258132 334516
rect 259532 356300 259588 356356
rect 257964 323260 258020 323316
rect 258076 327180 258132 327236
rect 261324 356188 261380 356244
rect 259644 355404 259700 355460
rect 259644 338380 259700 338436
rect 261212 351260 261268 351316
rect 259532 314412 259588 314468
rect 258076 314076 258132 314132
rect 257852 312284 257908 312340
rect 247996 312172 248052 312228
rect 261324 329420 261380 329476
rect 261436 342860 261492 342916
rect 261324 326060 261380 326116
rect 261324 313964 261380 314020
rect 263788 356636 263844 356692
rect 264572 355516 264628 355572
rect 263788 353500 263844 353556
rect 264460 353948 264516 354004
rect 263788 348572 263844 348628
rect 261660 338940 261716 338996
rect 262892 348460 262948 348516
rect 264460 343420 264516 343476
rect 263788 341740 263844 341796
rect 265356 353836 265412 353892
rect 264908 353724 264964 353780
rect 264684 353612 264740 353668
rect 265356 337820 265412 337876
rect 264908 332220 264964 332276
rect 264684 328300 264740 328356
rect 264572 326620 264628 326676
rect 262892 314636 262948 314692
rect 261436 312396 261492 312452
rect 261212 311948 261268 312004
rect 247772 311836 247828 311892
rect 138572 310940 138628 310996
rect 166236 311612 166292 311668
rect 166236 309820 166292 309876
rect 106204 305900 106260 305956
rect 81452 303100 81508 303156
rect 263900 298060 263956 298116
rect 263788 297500 263844 297556
rect 257852 296940 257908 296996
rect 225932 296604 225988 296660
rect 224812 295260 224868 295316
rect 224140 294140 224196 294196
rect 187292 289660 187348 289716
rect 166908 287868 166964 287924
rect 98812 287756 98868 287812
rect 98140 287532 98196 287588
rect 122668 287756 122724 287812
rect 105532 287644 105588 287700
rect 102172 285852 102228 285908
rect 106204 285964 106260 286020
rect 102844 284508 102900 284564
rect 101500 284396 101556 284452
rect 162876 287756 162932 287812
rect 143612 287420 143668 287476
rect 160860 284732 160916 284788
rect 164220 286076 164276 286132
rect 169596 287420 169652 287476
rect 168924 286300 168980 286356
rect 170940 286860 170996 286916
rect 143612 283276 143668 283332
rect 122668 283052 122724 283108
rect 108892 242956 108948 243012
rect 94108 242844 94164 242900
rect 106204 241612 106260 241668
rect 163548 239708 163604 239764
rect 162204 239596 162260 239652
rect 166236 241388 166292 241444
rect 167132 242732 167188 242788
rect 170268 240156 170324 240212
rect 223468 287308 223524 287364
rect 197372 285180 197428 285236
rect 192332 284284 192388 284340
rect 192332 241500 192388 241556
rect 187292 240156 187348 240212
rect 167132 239820 167188 239876
rect 228844 296380 228900 296436
rect 225932 287308 225988 287364
rect 228172 287308 228228 287364
rect 230860 294812 230916 294868
rect 232876 291900 232932 291956
rect 249676 288540 249732 288596
rect 247772 287868 247828 287924
rect 248108 287756 248164 287812
rect 248108 267932 248164 267988
rect 249452 285964 249508 286020
rect 247772 256060 247828 256116
rect 248108 267260 248164 267316
rect 249564 284508 249620 284564
rect 249564 276220 249620 276276
rect 249452 249900 249508 249956
rect 249564 265020 249620 265076
rect 248556 246540 248612 246596
rect 248444 246092 248500 246148
rect 222124 243068 222180 243124
rect 222796 240156 222852 240212
rect 197372 239596 197428 239652
rect 247884 240156 247940 240212
rect 249564 243068 249620 243124
rect 248556 241724 248612 241780
rect 248444 239932 248500 239988
rect 230860 239596 230916 239652
rect 165564 239260 165620 239316
rect 249452 239372 249508 239428
rect 225484 233100 225540 233156
rect 199052 231980 199108 232036
rect 195692 230860 195748 230916
rect 166236 229180 166292 229236
rect 163548 228620 163604 228676
rect 158844 226940 158900 226996
rect 133532 224140 133588 224196
rect 105532 219660 105588 219716
rect 102172 219100 102228 219156
rect 101500 215852 101556 215908
rect 83804 215292 83860 215348
rect 98140 215180 98196 215236
rect 99484 215068 99540 215124
rect 98812 213724 98868 213780
rect 104188 217420 104244 217476
rect 103516 215292 103572 215348
rect 106204 217980 106260 218036
rect 106876 215404 106932 215460
rect 99484 213164 99540 213220
rect 102844 212828 102900 212884
rect 83804 210924 83860 210980
rect 125132 211260 125188 211316
rect 102844 171612 102900 171668
rect 100156 171164 100212 171220
rect 141932 216860 141988 216916
rect 159516 215068 159572 215124
rect 164220 215628 164276 215684
rect 186396 215068 186452 215124
rect 166908 213836 166964 213892
rect 160188 212828 160244 212884
rect 186396 211148 186452 211204
rect 186508 174300 186564 174356
rect 185612 173180 185668 173236
rect 164892 171724 164948 171780
rect 141932 171276 141988 171332
rect 133532 171164 133588 171220
rect 125132 169372 125188 169428
rect 166908 171276 166964 171332
rect 162876 169372 162932 169428
rect 167580 170492 167636 170548
rect 162204 169148 162260 169204
rect 125132 166460 125188 166516
rect 88060 159180 88116 159236
rect 81452 158060 81508 158116
rect 105532 150556 105588 150612
rect 102508 143612 102564 143668
rect 102844 143052 102900 143108
rect 106876 144844 106932 144900
rect 99484 142044 99540 142100
rect 98588 141932 98644 141988
rect 130172 165900 130228 165956
rect 125132 101612 125188 101668
rect 125244 160300 125300 160356
rect 81452 101052 81508 101108
rect 99484 100828 99540 100884
rect 102844 100716 102900 100772
rect 106876 100604 106932 100660
rect 101500 100492 101556 100548
rect 104188 98812 104244 98868
rect 105532 98924 105588 98980
rect 104860 98700 104916 98756
rect 135212 161980 135268 162036
rect 133532 154140 133588 154196
rect 133532 100940 133588 100996
rect 130172 100604 130228 100660
rect 162876 150668 162932 150724
rect 161532 147084 161588 147140
rect 164220 147196 164276 147252
rect 168252 169260 168308 169316
rect 168364 170604 168420 170660
rect 222796 215740 222852 215796
rect 223468 215516 223524 215572
rect 228508 215852 228564 215908
rect 228508 214284 228564 214340
rect 228844 215068 228900 215124
rect 247996 215068 248052 215124
rect 226828 212828 226884 212884
rect 231532 212828 231588 212884
rect 247884 212492 247940 212548
rect 247772 207900 247828 207956
rect 246428 172620 246484 172676
rect 199052 171724 199108 171780
rect 230860 171724 230916 171780
rect 195692 171276 195748 171332
rect 223468 171276 223524 171332
rect 186508 170604 186564 170660
rect 200732 170940 200788 170996
rect 185612 147196 185668 147252
rect 187292 170380 187348 170436
rect 160860 100940 160916 100996
rect 165564 100940 165620 100996
rect 169596 100716 169652 100772
rect 192332 142380 192388 142436
rect 187404 141820 187460 141876
rect 187404 101724 187460 101780
rect 187292 100716 187348 100772
rect 170268 100604 170324 100660
rect 192332 100604 192388 100660
rect 135212 98812 135268 98868
rect 125244 98700 125300 98756
rect 168924 98812 168980 98868
rect 166236 98700 166292 98756
rect 229516 171164 229572 171220
rect 228172 171052 228228 171108
rect 226156 169596 226212 169652
rect 225484 169036 225540 169092
rect 204204 165452 204260 165508
rect 200844 140700 200900 140756
rect 200844 100940 200900 100996
rect 204092 100940 204148 100996
rect 200732 98700 200788 98756
rect 135436 97580 135492 97636
rect 110012 96572 110068 96628
rect 106204 91756 106260 91812
rect 104188 86604 104244 86660
rect 98812 78092 98868 78148
rect 83916 74060 83972 74116
rect 83916 71820 83972 71876
rect 100828 74844 100884 74900
rect 100156 74732 100212 74788
rect 102844 73500 102900 73556
rect 105532 74620 105588 74676
rect 167356 95340 167412 95396
rect 165564 90076 165620 90132
rect 135436 79772 135492 79828
rect 160860 86716 160916 86772
rect 110012 74844 110068 74900
rect 125132 79100 125188 79156
rect 122668 31276 122724 31332
rect 78092 28364 78148 28420
rect 74732 26796 74788 26852
rect 73052 26572 73108 26628
rect 62972 26460 63028 26516
rect 103516 26572 103572 26628
rect 89404 26460 89460 26516
rect 61292 26348 61348 26404
rect 107548 26796 107604 26852
rect 104188 26348 104244 26404
rect 134428 76300 134484 76356
rect 134428 74732 134484 74788
rect 162876 79772 162932 79828
rect 163548 74732 163604 74788
rect 167356 84924 167412 84980
rect 168252 88396 168308 88452
rect 167132 84700 167188 84756
rect 167132 74732 167188 74788
rect 187292 81900 187348 81956
rect 160860 28252 160916 28308
rect 125132 26796 125188 26852
rect 122668 26348 122724 26404
rect 187292 28252 187348 28308
rect 230188 160412 230244 160468
rect 228172 158732 228228 158788
rect 204204 98812 204260 98868
rect 205772 150332 205828 150388
rect 204092 26460 204148 26516
rect 226156 148540 226212 148596
rect 224812 145740 224868 145796
rect 228844 157052 228900 157108
rect 229516 147196 229572 147252
rect 248556 213612 248612 213668
rect 247996 207340 248052 207396
rect 248108 212380 248164 212436
rect 248556 210140 248612 210196
rect 248108 203980 248164 204036
rect 247884 200060 247940 200116
rect 247772 171052 247828 171108
rect 256172 287532 256228 287588
rect 252924 287308 252980 287364
rect 252812 284396 252868 284452
rect 249788 249340 249844 249396
rect 252924 263900 252980 263956
rect 252812 248220 252868 248276
rect 252924 258860 252980 258916
rect 249788 242956 249844 243012
rect 256284 285852 256340 285908
rect 256284 277900 256340 277956
rect 256172 252140 256228 252196
rect 256284 273756 256340 273812
rect 253036 247660 253092 247716
rect 253036 241612 253092 241668
rect 256284 240044 256340 240100
rect 252924 239708 252980 239764
rect 263788 296604 263844 296660
rect 263900 294812 263956 294868
rect 259532 288204 259588 288260
rect 258636 287644 258692 287700
rect 258076 286076 258132 286132
rect 257964 278460 258020 278516
rect 258636 280140 258692 280196
rect 258076 254940 258132 254996
rect 259532 245980 259588 246036
rect 261212 285964 261268 286020
rect 261436 285740 261492 285796
rect 261212 243740 261268 243796
rect 261324 273420 261380 273476
rect 257964 242844 258020 242900
rect 262892 284732 262948 284788
rect 264908 284172 264964 284228
rect 264572 283052 264628 283108
rect 261436 268940 261492 268996
rect 262892 274540 262948 274596
rect 261324 241836 261380 241892
rect 261548 260540 261604 260596
rect 261548 241388 261604 241444
rect 257852 239596 257908 239652
rect 263004 254380 263060 254436
rect 264572 251580 264628 251636
rect 264684 271180 264740 271236
rect 263788 247100 263844 247156
rect 263788 246092 263844 246148
rect 264684 242732 264740 242788
rect 264796 270060 264852 270116
rect 265020 283276 265076 283332
rect 265020 270620 265076 270676
rect 264908 268380 264964 268436
rect 265132 267932 265188 267988
rect 265132 255500 265188 255556
rect 264796 241052 264852 241108
rect 262892 239484 262948 239540
rect 263788 240380 263844 240436
rect 263788 239372 263844 239428
rect 249676 239260 249732 239316
rect 262892 238140 262948 238196
rect 261212 237580 261268 237636
rect 259532 237020 259588 237076
rect 256284 215964 256340 216020
rect 249676 215740 249732 215796
rect 249564 213500 249620 213556
rect 253036 215628 253092 215684
rect 249676 202860 249732 202916
rect 249788 213724 249844 213780
rect 252812 212604 252868 212660
rect 249900 212268 249956 212324
rect 249900 203420 249956 203476
rect 249788 195020 249844 195076
rect 252812 193900 252868 193956
rect 252924 208460 252980 208516
rect 249564 184380 249620 184436
rect 249676 192220 249732 192276
rect 249452 169596 249508 169652
rect 249564 175420 249620 175476
rect 246428 150668 246484 150724
rect 237692 149100 237748 149156
rect 237692 147196 237748 147252
rect 247772 144956 247828 145012
rect 248108 144844 248164 144900
rect 247996 142828 248052 142884
rect 248108 137340 248164 137396
rect 249452 144620 249508 144676
rect 248108 126812 248164 126868
rect 248332 126140 248388 126196
rect 249452 125580 249508 125636
rect 247996 123452 248052 123508
rect 247884 113372 247940 113428
rect 247772 104972 247828 105028
rect 230188 100716 230244 100772
rect 232876 100716 232932 100772
rect 231532 100604 231588 100660
rect 227500 98812 227556 98868
rect 232204 98700 232260 98756
rect 229516 95004 229572 95060
rect 228172 94892 228228 94948
rect 226716 93660 226772 93716
rect 226716 89964 226772 90020
rect 227612 90300 227668 90356
rect 225484 89740 225540 89796
rect 224140 74956 224196 75012
rect 223468 74844 223524 74900
rect 224812 74732 224868 74788
rect 225932 88620 225988 88676
rect 225932 74844 225988 74900
rect 227612 74732 227668 74788
rect 228844 74844 228900 74900
rect 232204 84924 232260 84980
rect 226828 29820 226884 29876
rect 222124 28252 222180 28308
rect 230188 29260 230244 29316
rect 231532 28140 231588 28196
rect 227500 26796 227556 26852
rect 249452 122220 249508 122276
rect 247996 99036 248052 99092
rect 248108 108332 248164 108388
rect 248108 74844 248164 74900
rect 247884 74732 247940 74788
rect 248332 74172 248388 74228
rect 248332 66780 248388 66836
rect 249676 171612 249732 171668
rect 252812 177100 252868 177156
rect 252700 139132 252756 139188
rect 252700 138908 252756 138964
rect 249564 100716 249620 100772
rect 249676 115500 249732 115556
rect 249452 29820 249508 29876
rect 249564 90860 249620 90916
rect 254492 213836 254548 213892
rect 254492 201180 254548 201236
rect 256172 202300 256228 202356
rect 253036 199500 253092 199556
rect 256508 215516 256564 215572
rect 256508 204540 256564 204596
rect 258188 215292 258244 215348
rect 258188 194460 258244 194516
rect 256284 187740 256340 187796
rect 257852 180460 257908 180516
rect 256172 169148 256228 169204
rect 256284 174860 256340 174916
rect 252924 169036 252980 169092
rect 256284 160412 256340 160468
rect 256172 143052 256228 143108
rect 256172 135660 256228 135716
rect 254492 132860 254548 132916
rect 252812 100604 252868 100660
rect 252924 114940 252980 114996
rect 249676 86716 249732 86772
rect 249788 100380 249844 100436
rect 249564 28140 249620 28196
rect 247772 26796 247828 26852
rect 252812 89180 252868 89236
rect 252700 70476 252756 70532
rect 252700 70028 252756 70084
rect 253036 110460 253092 110516
rect 256284 117180 256340 117236
rect 254492 100492 254548 100548
rect 256172 112700 256228 112756
rect 253036 90076 253092 90132
rect 252924 88396 252980 88452
rect 252812 29148 252868 29204
rect 249788 26684 249844 26740
rect 205772 26460 205828 26516
rect 169596 26348 169652 26404
rect 167580 26236 167636 26292
rect 256284 95004 256340 95060
rect 256396 106540 256452 106596
rect 257964 176540 258020 176596
rect 259756 215404 259812 215460
rect 259532 171276 259588 171332
rect 259644 212380 259700 212436
rect 259756 190540 259812 190596
rect 259644 169484 259700 169540
rect 259756 181020 259812 181076
rect 257964 158732 258020 158788
rect 261548 215180 261604 215236
rect 261436 212940 261492 212996
rect 261212 171724 261268 171780
rect 261324 198380 261380 198436
rect 261548 195580 261604 195636
rect 261436 183260 261492 183316
rect 261324 169372 261380 169428
rect 261436 172060 261492 172116
rect 259756 157052 259812 157108
rect 264572 234332 264628 234388
rect 263116 213388 263172 213444
rect 262892 171164 262948 171220
rect 263004 201740 263060 201796
rect 263788 211148 263844 211204
rect 263788 200620 263844 200676
rect 263116 187180 263172 187236
rect 263228 188860 263284 188916
rect 263004 169260 263060 169316
rect 263788 171500 263844 171556
rect 263788 170492 263844 170548
rect 263228 168924 263284 168980
rect 263788 169260 263844 169316
rect 263788 165452 263844 165508
rect 261548 165340 261604 165396
rect 261548 150556 261604 150612
rect 263004 164780 263060 164836
rect 261436 147084 261492 147140
rect 259644 146076 259700 146132
rect 258076 127596 258132 127652
rect 257852 101724 257908 101780
rect 257964 107660 258020 107716
rect 257068 93100 257124 93156
rect 257068 88172 257124 88228
rect 256396 86604 256452 86660
rect 259532 109228 259588 109284
rect 258076 98924 258132 98980
rect 258188 105420 258244 105476
rect 258188 91756 258244 91812
rect 257964 78092 258020 78148
rect 261436 123340 261492 123396
rect 259644 98812 259700 98868
rect 261212 116620 261268 116676
rect 261324 111020 261380 111076
rect 261436 94892 261492 94948
rect 262892 105308 262948 105364
rect 261324 79772 261380 79828
rect 261212 28252 261268 28308
rect 263788 153580 263844 153636
rect 263788 152012 263844 152068
rect 263004 100828 263060 100884
rect 263116 147756 263172 147812
rect 263788 131740 263844 131796
rect 263788 127596 263844 127652
rect 263900 127260 263956 127316
rect 263788 126812 263844 126868
rect 263788 125020 263844 125076
rect 263900 123452 263956 123508
rect 263116 98700 263172 98756
rect 263228 117740 263284 117796
rect 262892 26572 262948 26628
rect 263116 91532 263172 91588
rect 263788 112140 263844 112196
rect 263788 109228 263844 109284
rect 263788 102620 263844 102676
rect 263788 96572 263844 96628
rect 263788 94220 263844 94276
rect 263788 93324 263844 93380
rect 263228 84924 263284 84980
rect 264684 215180 264740 215236
rect 264908 214284 264964 214340
rect 264796 210812 264852 210868
rect 264908 192780 264964 192836
rect 265020 210924 265076 210980
rect 265020 186060 265076 186116
rect 264796 182700 264852 182756
rect 264684 173852 264740 173908
rect 264684 143612 264740 143668
rect 265132 141932 265188 141988
rect 264908 141708 264964 141764
rect 265356 141932 265412 141988
rect 265356 141596 265412 141652
rect 265132 135100 265188 135156
rect 264908 132300 264964 132356
rect 264684 131180 264740 131236
rect 264684 123900 264740 123956
rect 264908 119420 264964 119476
rect 264796 118860 264852 118916
rect 264908 113372 264964 113428
rect 264796 108332 264852 108388
rect 265020 108220 265076 108276
rect 265020 105308 265076 105364
rect 264684 104972 264740 105028
rect 277004 571900 277060 571956
rect 268156 571788 268212 571844
rect 267932 571676 267988 571732
rect 266476 571452 266532 571508
rect 266364 568652 266420 568708
rect 266364 431900 266420 431956
rect 266252 93212 266308 93268
rect 266364 361228 266420 361284
rect 264684 78540 264740 78596
rect 264684 31276 264740 31332
rect 264908 66220 264964 66276
rect 264908 31164 264964 31220
rect 264572 28252 264628 28308
rect 265468 31052 265524 31108
rect 266588 569436 266644 569492
rect 266588 304892 266644 304948
rect 275884 571564 275940 571620
rect 273644 570556 273700 570612
rect 269164 570108 269220 570164
rect 274764 570220 274820 570276
rect 280364 577052 280420 577108
rect 283724 576156 283780 576212
rect 281484 575484 281540 575540
rect 282604 574364 282660 574420
rect 288092 590604 288148 590660
rect 287084 590492 287140 590548
rect 284732 574476 284788 574532
rect 284844 577164 284900 577220
rect 285964 574476 286020 574532
rect 289772 590492 289828 590548
rect 288092 574364 288148 574420
rect 288204 583772 288260 583828
rect 297836 590492 297892 590548
rect 303212 590492 303268 590548
rect 289772 576156 289828 576212
rect 303212 575484 303268 575540
rect 305004 588588 305060 588644
rect 299404 572236 299460 572292
rect 296492 572012 296548 572068
rect 296492 570668 296548 570724
rect 298284 570668 298340 570724
rect 294924 570444 294980 570500
rect 292684 570332 292740 570388
rect 290444 569772 290500 569828
rect 293804 569772 293860 569828
rect 296044 569884 296100 569940
rect 296940 569660 296996 569716
rect 291564 569212 291620 569268
rect 303660 569548 303716 569604
rect 307244 583772 307300 583828
rect 306124 573804 306180 573860
rect 311724 582204 311780 582260
rect 309484 578844 309540 578900
rect 308364 577164 308420 577220
rect 310604 574028 310660 574084
rect 364028 590604 364084 590660
rect 407372 591276 407428 591332
rect 341964 578844 342020 578900
rect 315084 578732 315140 578788
rect 312844 573916 312900 573972
rect 313964 573692 314020 573748
rect 408268 591276 408324 591332
rect 430220 590492 430276 590548
rect 432572 590492 432628 590548
rect 407372 577164 407428 577220
rect 496412 590492 496468 590548
rect 499772 590492 499828 590548
rect 474348 583772 474404 583828
rect 499772 582092 499828 582148
rect 432572 577052 432628 577108
rect 562604 590492 562660 590548
rect 540540 573804 540596 573860
rect 328524 572348 328580 572404
rect 325164 572012 325220 572068
rect 315756 571900 315812 571956
rect 315756 569996 315812 570052
rect 317324 571788 317380 571844
rect 315868 569548 315924 569604
rect 324044 571228 324100 571284
rect 322924 569436 322980 569492
rect 327404 571676 327460 571732
rect 326284 571452 326340 571508
rect 335244 572236 335300 572292
rect 329644 572124 329700 572180
rect 330764 571228 330820 571284
rect 333676 570220 333732 570276
rect 333452 570108 333508 570164
rect 317772 569324 317828 569380
rect 320684 569100 320740 569156
rect 321804 568988 321860 569044
rect 270284 568876 270340 568932
rect 271404 568876 271460 568932
rect 272524 568876 272580 568932
rect 289324 568876 289380 568932
rect 300524 568876 300580 568932
rect 301644 568876 301700 568932
rect 302764 568876 302820 568932
rect 319564 568876 319620 568932
rect 268156 516572 268212 516628
rect 267932 296492 267988 296548
rect 333564 567756 333620 567812
rect 335132 568540 335188 568596
rect 334460 518364 334516 518420
rect 334460 514220 334516 514276
rect 338716 571900 338772 571956
rect 336924 571788 336980 571844
rect 335468 571564 335524 571620
rect 336812 570444 336868 570500
rect 335468 528332 335524 528388
rect 335916 530012 335972 530068
rect 335916 527100 335972 527156
rect 335916 526652 335972 526708
rect 335916 524860 335972 524916
rect 335244 521612 335300 521668
rect 335132 509292 335188 509348
rect 335244 514892 335300 514948
rect 335132 501564 335188 501620
rect 335244 490700 335300 490756
rect 335132 482860 335188 482916
rect 335580 484652 335636 484708
rect 335580 475580 335636 475636
rect 335132 472780 335188 472836
rect 334460 472220 334516 472276
rect 334460 469532 334516 469588
rect 335132 453516 335188 453572
rect 333676 443212 333732 443268
rect 335804 444332 335860 444388
rect 334460 439292 334516 439348
rect 334460 435260 334516 435316
rect 335132 437724 335188 437780
rect 334460 426524 334516 426580
rect 334460 422380 334516 422436
rect 335804 436940 335860 436996
rect 335244 434252 335300 434308
rect 335244 417900 335300 417956
rect 335468 432684 335524 432740
rect 335468 416780 335524 416836
rect 335132 415660 335188 415716
rect 335132 413980 335188 414036
rect 335132 387548 335188 387604
rect 335356 410620 335412 410676
rect 335580 408380 335636 408436
rect 335580 387436 335636 387492
rect 336028 388780 336084 388836
rect 335356 387324 335412 387380
rect 336028 385644 336084 385700
rect 335916 384860 335972 384916
rect 335916 383852 335972 383908
rect 335916 362124 335972 362180
rect 335916 359100 335972 359156
rect 334348 356188 334404 356244
rect 335132 355628 335188 355684
rect 334348 353500 334404 353556
rect 334460 353612 334516 353668
rect 334460 349580 334516 349636
rect 335132 346220 335188 346276
rect 335244 353836 335300 353892
rect 335132 338492 335188 338548
rect 334460 325500 334516 325556
rect 334460 314188 334516 314244
rect 335468 353724 335524 353780
rect 335244 315980 335300 316036
rect 335356 350140 335412 350196
rect 335468 348460 335524 348516
rect 335356 314636 335412 314692
rect 335468 321020 335524 321076
rect 335468 313292 335524 313348
rect 335692 318332 335748 318388
rect 335692 312620 335748 312676
rect 335132 300300 335188 300356
rect 334460 298060 334516 298116
rect 334348 297500 334404 297556
rect 334460 296492 334516 296548
rect 334348 294812 334404 294868
rect 333564 284620 333620 284676
rect 335132 286412 335188 286468
rect 336028 284172 336084 284228
rect 336028 279020 336084 279076
rect 335132 257180 335188 257236
rect 335244 266700 335300 266756
rect 333452 244972 333508 245028
rect 335468 265580 335524 265636
rect 335356 263340 335412 263396
rect 335356 246092 335412 246148
rect 335468 240044 335524 240100
rect 335244 239596 335300 239652
rect 266476 234444 266532 234500
rect 334348 239260 334404 239316
rect 334460 238140 334516 238196
rect 334460 236012 334516 236068
rect 334348 232652 334404 232708
rect 337148 571676 337204 571732
rect 336924 485100 336980 485156
rect 337036 498204 337092 498260
rect 338492 571452 338548 571508
rect 337596 531580 337652 531636
rect 337596 525756 337652 525812
rect 337148 486220 337204 486276
rect 337260 503692 337316 503748
rect 337708 503132 337764 503188
rect 337708 500780 337764 500836
rect 337260 477820 337316 477876
rect 338492 476700 338548 476756
rect 338604 500780 338660 500836
rect 338492 469980 338548 470036
rect 338492 453292 338548 453348
rect 337036 453180 337092 453236
rect 336924 430332 336980 430388
rect 336924 407260 336980 407316
rect 338492 426860 338548 426916
rect 557564 571900 557620 571956
rect 433468 571788 433524 571844
rect 351932 571564 351988 571620
rect 341852 571340 341908 571396
rect 340172 570332 340228 570388
rect 339276 511756 339332 511812
rect 339276 508620 339332 508676
rect 338716 494620 338772 494676
rect 338828 499324 338884 499380
rect 338828 443660 338884 443716
rect 338604 418460 338660 418516
rect 338716 430220 338772 430276
rect 338716 406700 338772 406756
rect 338492 399980 338548 400036
rect 339276 358652 339332 358708
rect 337148 357084 337204 357140
rect 336924 356748 336980 356804
rect 339276 356188 339332 356244
rect 338604 355516 338660 355572
rect 337148 313740 337204 313796
rect 338492 351820 338548 351876
rect 338604 343980 338660 344036
rect 338492 311612 338548 311668
rect 336924 304780 336980 304836
rect 338604 287308 338660 287364
rect 338492 271740 338548 271796
rect 336924 260428 336980 260484
rect 338716 285628 338772 285684
rect 338716 267820 338772 267876
rect 338604 265020 338660 265076
rect 338492 243292 338548 243348
rect 336924 239708 336980 239764
rect 336812 231868 336868 231924
rect 338492 237580 338548 237636
rect 338492 227612 338548 227668
rect 336812 215740 336868 215796
rect 335244 215628 335300 215684
rect 335132 208460 335188 208516
rect 335244 207340 335300 207396
rect 335356 211036 335412 211092
rect 335132 177996 335188 178052
rect 335244 202860 335300 202916
rect 335916 210812 335972 210868
rect 335916 205660 335972 205716
rect 335356 198380 335412 198436
rect 335244 173964 335300 174020
rect 335356 179340 335412 179396
rect 335356 172172 335412 172228
rect 338492 215516 338548 215572
rect 339276 213612 339332 213668
rect 339276 209580 339332 209636
rect 338492 195580 338548 195636
rect 336812 171164 336868 171220
rect 338492 188300 338548 188356
rect 338716 177996 338772 178052
rect 338716 169484 338772 169540
rect 338492 169372 338548 169428
rect 334460 168700 334516 168756
rect 334460 167132 334516 167188
rect 336924 168140 336980 168196
rect 336028 154140 336084 154196
rect 336028 150332 336084 150388
rect 334460 147980 334516 148036
rect 334460 146972 334516 147028
rect 335244 143724 335300 143780
rect 335132 140700 335188 140756
rect 334460 140476 334516 140532
rect 334460 139020 334516 139076
rect 334348 113820 334404 113876
rect 336812 142044 336868 142100
rect 335244 137340 335300 137396
rect 335804 140700 335860 140756
rect 335804 135100 335860 135156
rect 335356 133980 335412 134036
rect 336812 129500 336868 129556
rect 335356 113372 335412 113428
rect 335692 116060 335748 116116
rect 335692 112812 335748 112868
rect 335132 110012 335188 110068
rect 334348 107436 334404 107492
rect 336812 107436 336868 107492
rect 267708 101612 267764 101668
rect 267708 101164 267764 101220
rect 335916 79100 335972 79156
rect 335916 78316 335972 78372
rect 335132 77420 335188 77476
rect 334460 68572 334516 68628
rect 334460 67788 334516 67844
rect 335356 72380 335412 72436
rect 335356 59612 335412 59668
rect 335132 31052 335188 31108
rect 270060 29932 270116 29988
rect 274316 29708 274372 29764
rect 278572 29596 278628 29652
rect 282828 29484 282884 29540
rect 291340 29372 291396 29428
rect 266364 29148 266420 29204
rect 295596 29260 295652 29316
rect 304108 29036 304164 29092
rect 299852 28476 299908 28532
rect 287084 28364 287140 28420
rect 308364 28252 308420 28308
rect 265468 26684 265524 26740
rect 263116 26572 263172 26628
rect 321132 26684 321188 26740
rect 316876 26572 316932 26628
rect 312620 26460 312676 26516
rect 259532 26348 259588 26404
rect 256172 26236 256228 26292
rect 10892 26124 10948 26180
rect 325388 26124 325444 26180
rect 4172 24332 4228 24388
rect 339276 153020 339332 153076
rect 350252 571228 350308 571284
rect 341852 531020 341908 531076
rect 345212 570108 345268 570164
rect 340284 521836 340340 521892
rect 342636 516796 342692 516852
rect 342636 511420 342692 511476
rect 342076 507052 342132 507108
rect 340284 480620 340340 480676
rect 340396 500668 340452 500724
rect 340284 469420 340340 469476
rect 340396 468300 340452 468356
rect 341852 499212 341908 499268
rect 340284 453180 340340 453236
rect 341964 497756 342020 497812
rect 345324 568876 345380 568932
rect 345324 506940 345380 506996
rect 349356 555212 349412 555268
rect 346892 503356 346948 503412
rect 345212 502460 345268 502516
rect 345548 503244 345604 503300
rect 342076 478940 342132 478996
rect 345212 501004 345268 501060
rect 341964 467180 342020 467236
rect 342076 469532 342132 469588
rect 342636 466060 342692 466116
rect 342636 457772 342692 457828
rect 342076 453404 342132 453460
rect 341852 448700 341908 448756
rect 345324 499436 345380 499492
rect 345436 498092 345492 498148
rect 346892 486780 346948 486836
rect 348572 499548 348628 499604
rect 345548 482300 345604 482356
rect 348572 467740 348628 467796
rect 350364 569548 350420 569604
rect 350364 506380 350420 506436
rect 350588 508172 350644 508228
rect 350252 484652 350308 484708
rect 350364 500892 350420 500948
rect 349356 483308 349412 483364
rect 345436 465500 345492 465556
rect 345436 464940 345492 464996
rect 345436 453068 345492 453124
rect 345324 445340 345380 445396
rect 345212 432684 345268 432740
rect 345436 444892 345492 444948
rect 345212 430108 345268 430164
rect 340284 428428 340340 428484
rect 342076 426748 342132 426804
rect 340284 404460 340340 404516
rect 341852 426188 341908 426244
rect 342076 406140 342132 406196
rect 341852 393260 341908 393316
rect 341852 389900 341908 389956
rect 341852 384188 341908 384244
rect 345324 428652 345380 428708
rect 345436 421820 345492 421876
rect 350252 463820 350308 463876
rect 350252 455084 350308 455140
rect 350252 446012 350308 446068
rect 350476 498988 350532 499044
rect 350588 492380 350644 492436
rect 374220 571452 374276 571508
rect 370860 571228 370916 571284
rect 407372 571452 407428 571508
rect 380268 570108 380324 570164
rect 374892 569548 374948 569604
rect 352044 568988 352100 569044
rect 372204 568988 372260 569044
rect 377580 568876 377636 568932
rect 400652 567644 400708 567700
rect 393932 567532 393988 567588
rect 357868 527772 357924 527828
rect 357868 527436 357924 527492
rect 368732 523404 368788 523460
rect 356188 521724 356244 521780
rect 356188 516460 356244 516516
rect 370188 507052 370244 507108
rect 372092 523516 372148 523572
rect 372092 505820 372148 505876
rect 368732 505260 368788 505316
rect 352044 504140 352100 504196
rect 372204 503692 372260 503748
rect 376908 523516 376964 523572
rect 377580 523404 377636 523460
rect 379708 523404 379764 523460
rect 379708 520380 379764 520436
rect 381388 516908 381444 516964
rect 381388 515340 381444 515396
rect 376236 503132 376292 503188
rect 370188 501004 370244 501060
rect 368172 499436 368228 499492
rect 352156 499100 352212 499156
rect 351932 489020 351988 489076
rect 352044 497868 352100 497924
rect 351036 462700 351092 462756
rect 351036 457884 351092 457940
rect 351932 462140 351988 462196
rect 351932 455196 351988 455252
rect 369516 499324 369572 499380
rect 368844 498988 368900 499044
rect 372876 500780 372932 500836
rect 374220 499212 374276 499268
rect 376236 497868 376292 497924
rect 352156 466620 352212 466676
rect 352492 463260 352548 463316
rect 352604 461580 352660 461636
rect 352604 456540 352660 456596
rect 352492 456428 352548 456484
rect 352044 448140 352100 448196
rect 350476 446460 350532 446516
rect 369628 451612 369684 451668
rect 370188 446012 370244 446068
rect 372092 451948 372148 452004
rect 369628 445900 369684 445956
rect 371308 444444 371364 444500
rect 371308 441980 371364 442036
rect 369516 437724 369572 437780
rect 373548 451948 373604 452004
rect 374220 451612 374276 451668
rect 375452 451052 375508 451108
rect 377580 444892 377636 444948
rect 375452 436380 375508 436436
rect 372092 434252 372148 434308
rect 350364 422940 350420 422996
rect 351932 430444 351988 430500
rect 350252 417340 350308 417396
rect 349356 411404 349412 411460
rect 348572 408940 348628 408996
rect 345324 394940 345380 394996
rect 345436 400540 345492 400596
rect 347788 391020 347844 391076
rect 347788 385756 347844 385812
rect 345436 385308 345492 385364
rect 348572 383964 348628 384020
rect 345212 361340 345268 361396
rect 342636 360332 342692 360388
rect 342636 358540 342692 358596
rect 340284 358316 340340 358372
rect 341852 357980 341908 358036
rect 340396 333900 340452 333956
rect 348684 357868 348740 357924
rect 341964 356636 342020 356692
rect 345436 356412 345492 356468
rect 345324 355292 345380 355348
rect 341964 330540 342020 330596
rect 345212 347340 345268 347396
rect 341852 324940 341908 324996
rect 340396 313740 340452 313796
rect 341852 318220 341908 318276
rect 345436 344540 345492 344596
rect 345324 331100 345380 331156
rect 348572 339500 348628 339556
rect 345212 314412 345268 314468
rect 345324 323260 345380 323316
rect 341852 313516 341908 313572
rect 349244 355852 349300 355908
rect 349244 355180 349300 355236
rect 348684 338492 348740 338548
rect 350252 403340 350308 403396
rect 350252 385420 350308 385476
rect 350364 397740 350420 397796
rect 350364 384412 350420 384468
rect 350588 390460 350644 390516
rect 350588 384300 350644 384356
rect 351148 387100 351204 387156
rect 351148 384076 351204 384132
rect 374892 430444 374948 430500
rect 376908 430108 376964 430164
rect 352044 426300 352100 426356
rect 352044 405020 352100 405076
rect 352044 401996 352100 402052
rect 352492 391580 352548 391636
rect 352492 385196 352548 385252
rect 352604 389340 352660 389396
rect 370860 385868 370916 385924
rect 370188 385644 370244 385700
rect 352604 385084 352660 385140
rect 352044 384524 352100 384580
rect 369068 385084 369124 385140
rect 374220 385756 374276 385812
rect 370860 384636 370916 384692
rect 368844 384188 368900 384244
rect 352716 383852 352772 383908
rect 352716 382956 352772 383012
rect 351932 362124 351988 362180
rect 372876 385308 372932 385364
rect 376908 384636 376964 384692
rect 375564 384300 375620 384356
rect 374892 384076 374948 384132
rect 373548 382956 373604 383012
rect 395164 504812 395220 504868
rect 395164 496300 395220 496356
rect 398972 501004 399028 501060
rect 394044 451164 394100 451220
rect 394044 434140 394100 434196
rect 412412 571228 412468 571284
rect 430780 571228 430836 571284
rect 412524 570108 412580 570164
rect 412524 510860 412580 510916
rect 414092 569548 414148 569604
rect 474684 571788 474740 571844
rect 438172 571676 438228 571732
rect 435484 570108 435540 570164
rect 435708 569548 435764 569604
rect 464492 571676 464548 571732
rect 428092 516796 428148 516852
rect 414092 509180 414148 509236
rect 430108 503356 430164 503412
rect 435484 521836 435540 521892
rect 440188 518364 440244 518420
rect 436828 516908 436884 516964
rect 471212 569996 471268 570052
rect 471212 523180 471268 523236
rect 474572 569660 474628 569716
rect 464492 514892 464548 514948
rect 442204 511756 442260 511812
rect 434812 503244 434868 503300
rect 412412 501564 412468 501620
rect 436156 501004 436212 501060
rect 407372 495180 407428 495236
rect 407484 500780 407540 500836
rect 412412 499212 412468 499268
rect 432796 499212 432852 499268
rect 438844 500892 438900 500948
rect 464492 499212 464548 499268
rect 434812 498204 434868 498260
rect 412412 457660 412468 457716
rect 430780 455980 430836 456036
rect 407484 438620 407540 438676
rect 412412 447916 412468 447972
rect 412412 434700 412468 434756
rect 464492 431340 464548 431396
rect 400652 430108 400708 430164
rect 412412 430444 412468 430500
rect 407372 426636 407428 426692
rect 398972 426524 399028 426580
rect 399196 426524 399252 426580
rect 399196 382060 399252 382116
rect 404012 426076 404068 426132
rect 407372 370860 407428 370916
rect 404012 368060 404068 368116
rect 436156 430444 436212 430500
rect 435484 428652 435540 428708
rect 467852 430444 467908 430500
rect 462812 428540 462868 428596
rect 436828 426972 436884 427028
rect 438172 426972 438228 427028
rect 430780 384412 430836 384468
rect 467852 382620 467908 382676
rect 462812 378140 462868 378196
rect 412412 365820 412468 365876
rect 393932 363916 393988 363972
rect 377580 360332 377636 360388
rect 372204 359660 372260 359716
rect 402332 358428 402388 358484
rect 370860 358316 370916 358372
rect 349356 341628 349412 341684
rect 348572 313628 348628 313684
rect 348684 322140 348740 322196
rect 345324 312284 345380 312340
rect 348684 311948 348740 312004
rect 340284 301420 340340 301476
rect 340284 288540 340340 288596
rect 341852 287756 341908 287812
rect 340284 241724 340340 241780
rect 340396 262220 340452 262276
rect 342076 287532 342132 287588
rect 348684 285852 348740 285908
rect 345324 284284 345380 284340
rect 345212 281260 345268 281316
rect 342076 249900 342132 249956
rect 342188 277340 342244 277396
rect 341852 243180 341908 243236
rect 342188 242956 342244 243012
rect 345324 276220 345380 276276
rect 348572 280140 348628 280196
rect 345212 241612 345268 241668
rect 347788 246092 347844 246148
rect 340396 239932 340452 239988
rect 348684 277900 348740 277956
rect 348572 243068 348628 243124
rect 350252 358204 350308 358260
rect 352716 358092 352772 358148
rect 352716 356860 352772 356916
rect 369516 357868 369572 357924
rect 352380 356524 352436 356580
rect 352156 356188 352212 356244
rect 351932 355964 351988 356020
rect 351932 349020 351988 349076
rect 350252 318332 350308 318388
rect 350364 347900 350420 347956
rect 351932 346780 351988 346836
rect 350588 328300 350644 328356
rect 350364 313964 350420 314020
rect 350476 319340 350532 319396
rect 351932 314524 351988 314580
rect 352044 342860 352100 342916
rect 350588 314076 350644 314132
rect 393148 358316 393204 358372
rect 372876 356748 372932 356804
rect 378252 356636 378308 356692
rect 374220 356188 374276 356244
rect 374892 355292 374948 355348
rect 393148 353836 393204 353892
rect 398972 356748 399028 356804
rect 352380 341740 352436 341796
rect 352156 332220 352212 332276
rect 352268 332780 352324 332836
rect 352044 313852 352100 313908
rect 352156 317660 352212 317716
rect 350476 312172 350532 312228
rect 359436 314076 359492 314132
rect 352268 313404 352324 313460
rect 352156 311724 352212 311780
rect 370188 303100 370244 303156
rect 374220 313404 374276 313460
rect 398972 310940 399028 310996
rect 400652 356636 400708 356692
rect 400652 310380 400708 310436
rect 439516 358428 439572 358484
rect 410732 357868 410788 357924
rect 404796 314188 404852 314244
rect 404796 311836 404852 311892
rect 402332 309820 402388 309876
rect 435484 357868 435540 357924
rect 432124 356748 432180 356804
rect 410732 308140 410788 308196
rect 412412 356188 412468 356244
rect 430780 356188 430836 356244
rect 436156 356636 436212 356692
rect 430108 309260 430164 309316
rect 412412 307020 412468 307076
rect 434812 313628 434868 313684
rect 436156 312060 436212 312116
rect 444220 313740 444276 313796
rect 437500 311500 437556 311556
rect 501564 571788 501620 571844
rect 498204 571676 498260 571732
rect 496188 571564 496244 571620
rect 476252 569660 476308 569716
rect 474684 521500 474740 521556
rect 474796 569548 474852 569604
rect 492268 569660 492324 569716
rect 494844 569548 494900 569604
rect 500892 569996 500948 570052
rect 533372 571564 533428 571620
rect 555548 571340 555604 571396
rect 533372 530012 533428 530068
rect 536732 571228 536788 571284
rect 475468 523292 475524 523348
rect 476140 520940 476196 520996
rect 475468 519820 475524 519876
rect 474796 517580 474852 517636
rect 498204 523404 498260 523460
rect 554204 571228 554260 571284
rect 558236 571564 558292 571620
rect 558908 571452 558964 571508
rect 590492 570668 590548 570724
rect 580636 570556 580692 570612
rect 580412 569772 580468 569828
rect 539196 529340 539252 529396
rect 539196 527772 539252 527828
rect 556892 527772 556948 527828
rect 536732 526652 536788 526708
rect 559580 527660 559636 527716
rect 557564 527436 557620 527492
rect 554876 525756 554932 525812
rect 562268 525420 562324 525476
rect 499548 523292 499604 523348
rect 494844 521724 494900 521780
rect 493500 508172 493556 508228
rect 564284 524300 564340 524356
rect 563612 504812 563668 504868
rect 536732 501004 536788 501060
rect 476252 500892 476308 500948
rect 474684 497868 474740 497924
rect 474684 458220 474740 458276
rect 498876 500892 498932 500948
rect 493500 499212 493556 499268
rect 530012 500892 530068 500948
rect 492828 498092 492884 498148
rect 494172 497868 494228 497924
rect 496860 457100 496916 457156
rect 494844 456540 494900 456596
rect 493500 455084 493556 455140
rect 496188 456428 496244 456484
rect 498876 453068 498932 453124
rect 494172 451164 494228 451220
rect 501564 455196 501620 455252
rect 499548 447916 499604 447972
rect 530012 440860 530068 440916
rect 533372 497868 533428 497924
rect 476252 439292 476308 439348
rect 558908 501004 558964 501060
rect 558236 500780 558292 500836
rect 554876 500668 554932 500724
rect 556220 499100 556276 499156
rect 562268 500892 562324 500948
rect 562940 499548 562996 499604
rect 555548 497868 555604 497924
rect 564284 497756 564340 497812
rect 558908 456988 558964 457044
rect 555548 453292 555604 453348
rect 556220 453180 556276 453236
rect 562268 453516 562324 453572
rect 562940 453404 562996 453460
rect 561596 451052 561652 451108
rect 559580 444444 559636 444500
rect 536732 444332 536788 444388
rect 533372 437500 533428 437556
rect 561596 430444 561652 430500
rect 494172 430332 494228 430388
rect 503580 430220 503636 430276
rect 500892 428428 500948 428484
rect 560252 428540 560308 428596
rect 474684 426972 474740 427028
rect 556220 426972 556276 427028
rect 493500 426860 493556 426916
rect 500220 426748 500276 426804
rect 497532 426636 497588 426692
rect 557564 426524 557620 426580
rect 502908 426412 502964 426468
rect 535836 408716 535892 408772
rect 495516 385420 495572 385476
rect 474684 380380 474740 380436
rect 493500 374220 493556 374276
rect 499548 385308 499604 385364
rect 498876 384524 498932 384580
rect 498204 373100 498260 373156
rect 498204 358316 498260 358372
rect 493500 358204 493556 358260
rect 475468 357868 475524 357924
rect 494844 357868 494900 357924
rect 497532 356412 497588 356468
rect 495628 355964 495684 356020
rect 500220 357084 500276 357140
rect 500892 356524 500948 356580
rect 501116 355628 501172 355684
rect 499548 355516 499604 355572
rect 475468 353724 475524 353780
rect 535948 387548 536004 387604
rect 537740 387436 537796 387492
rect 537628 387324 537684 387380
rect 537628 382956 537684 383012
rect 535948 382844 536004 382900
rect 537740 382732 537796 382788
rect 559580 383964 559636 384020
rect 558908 382956 558964 383012
rect 554204 382844 554260 382900
rect 553532 382732 553588 382788
rect 560252 378700 560308 378756
rect 558908 358652 558964 358708
rect 539196 358204 539252 358260
rect 557564 357980 557620 358036
rect 566972 358204 567028 358260
rect 562940 358092 562996 358148
rect 539196 353612 539252 353668
rect 535836 341628 535892 341684
rect 561036 314636 561092 314692
rect 500892 314524 500948 314580
rect 493500 314412 493556 314468
rect 496188 313852 496244 313908
rect 499772 313964 499828 314020
rect 499548 313516 499604 313572
rect 553532 311948 553588 312004
rect 558124 313292 558180 313348
rect 557788 312284 557844 312340
rect 554876 311836 554932 311892
rect 496860 311724 496916 311780
rect 562940 314076 562996 314132
rect 562268 312172 562324 312228
rect 560924 311612 560980 311668
rect 474572 311052 474628 311108
rect 433468 308700 433524 308756
rect 430780 306460 430836 306516
rect 376236 304220 376292 304276
rect 373548 303660 373604 303716
rect 372204 301980 372260 302036
rect 400652 298620 400708 298676
rect 351932 288092 351988 288148
rect 349356 268380 349412 268436
rect 347788 239820 347844 239876
rect 348572 215292 348628 215348
rect 340284 215180 340340 215236
rect 345548 213500 345604 213556
rect 342076 212940 342132 212996
rect 340284 206780 340340 206836
rect 341852 212380 341908 212436
rect 340284 205100 340340 205156
rect 342076 203980 342132 204036
rect 345212 199500 345268 199556
rect 341852 186060 341908 186116
rect 341964 190988 342020 191044
rect 340284 169596 340340 169652
rect 340396 182140 340452 182196
rect 341852 178220 341908 178276
rect 345212 171276 345268 171332
rect 345324 192780 345380 192836
rect 348572 200060 348628 200116
rect 345548 191660 345604 191716
rect 350252 287644 350308 287700
rect 350476 287420 350532 287476
rect 350476 259420 350532 259476
rect 350252 249340 350308 249396
rect 350364 253260 350420 253316
rect 349468 245420 349524 245476
rect 349468 241836 349524 241892
rect 376236 287756 376292 287812
rect 352268 285964 352324 286020
rect 352156 284396 352212 284452
rect 351932 242844 351988 242900
rect 352044 271180 352100 271236
rect 350364 241388 350420 241444
rect 375564 285964 375620 286020
rect 368844 285628 368900 285684
rect 376908 284396 376964 284452
rect 352268 270620 352324 270676
rect 352156 269500 352212 269556
rect 352156 252140 352212 252196
rect 374892 243292 374948 243348
rect 352156 243180 352212 243236
rect 352044 241276 352100 241332
rect 359548 242060 359604 242116
rect 370188 241836 370244 241892
rect 359548 240156 359604 240212
rect 563724 296940 563780 296996
rect 504812 296492 504868 296548
rect 499772 294812 499828 294868
rect 518252 296380 518308 296436
rect 560364 295820 560420 295876
rect 518252 289772 518308 289828
rect 559468 289772 559524 289828
rect 504812 288204 504868 288260
rect 556108 288204 556164 288260
rect 499772 288092 499828 288148
rect 498876 287980 498932 288036
rect 436828 287644 436884 287700
rect 433468 285852 433524 285908
rect 438732 287532 438788 287588
rect 477148 287532 477204 287588
rect 477148 286412 477204 286468
rect 498204 287420 498260 287476
rect 475468 285740 475524 285796
rect 434812 284284 434868 284340
rect 432796 284172 432852 284228
rect 501564 287532 501620 287588
rect 500220 286300 500276 286356
rect 499548 285628 499604 285684
rect 500892 285740 500948 285796
rect 554428 287308 554484 287364
rect 561708 288092 561764 288148
rect 475468 283500 475524 283556
rect 438844 243180 438900 243236
rect 436828 243068 436884 243124
rect 448924 242956 448980 243012
rect 400652 241836 400708 241892
rect 432124 241612 432180 241668
rect 493500 242844 493556 242900
rect 494172 241724 494228 241780
rect 434812 241388 434868 241444
rect 375564 241276 375620 241332
rect 372876 240156 372932 240212
rect 496188 239708 496244 239764
rect 503132 240380 503188 240436
rect 350252 233100 350308 233156
rect 437612 232540 437668 232596
rect 427532 224700 427588 224756
rect 414092 224140 414148 224196
rect 350252 222572 350308 222628
rect 406588 223020 406644 223076
rect 398972 220220 399028 220276
rect 372876 216860 372932 216916
rect 352156 215404 352212 215460
rect 350364 215068 350420 215124
rect 349356 198492 349412 198548
rect 345324 169260 345380 169316
rect 348572 181580 348628 181636
rect 341964 169148 342020 169204
rect 341852 162092 341908 162148
rect 341964 167020 342020 167076
rect 340396 160412 340452 160468
rect 341964 158844 342020 158900
rect 340172 152460 340228 152516
rect 340284 153580 340340 153636
rect 339276 152124 339332 152180
rect 338492 151900 338548 151956
rect 338604 144508 338660 144564
rect 338604 136780 338660 136836
rect 338492 101724 338548 101780
rect 340172 112812 340228 112868
rect 336924 100940 336980 100996
rect 338604 100380 338660 100436
rect 338492 94220 338548 94276
rect 336812 26796 336868 26852
rect 337036 69580 337092 69636
rect 338604 89964 338660 90020
rect 338716 93100 338772 93156
rect 338716 29596 338772 29652
rect 338492 29372 338548 29428
rect 340284 101836 340340 101892
rect 340396 143500 340452 143556
rect 342076 142828 342132 142884
rect 341964 130620 342020 130676
rect 340396 98812 340452 98868
rect 340508 111020 340564 111076
rect 340508 94892 340564 94948
rect 341852 108220 341908 108276
rect 342076 128940 342132 128996
rect 345212 142156 345268 142212
rect 345212 125020 345268 125076
rect 345324 123900 345380 123956
rect 342188 117740 342244 117796
rect 341964 100604 342020 100660
rect 342076 114940 342132 114996
rect 345212 115500 345268 115556
rect 343532 110012 343588 110068
rect 343532 98700 343588 98756
rect 342188 96684 342244 96740
rect 342076 86492 342132 86548
rect 341852 29260 341908 29316
rect 346892 113372 346948 113428
rect 348684 144732 348740 144788
rect 348684 136220 348740 136276
rect 350252 212492 350308 212548
rect 351932 213724 351988 213780
rect 350476 213388 350532 213444
rect 350476 196700 350532 196756
rect 350364 188860 350420 188916
rect 352044 213276 352100 213332
rect 350252 183820 350308 183876
rect 350588 187180 350644 187236
rect 349356 127932 349412 127988
rect 348572 98924 348628 98980
rect 348684 119420 348740 119476
rect 346892 98588 346948 98644
rect 345324 93212 345380 93268
rect 348684 78092 348740 78148
rect 348572 74172 348628 74228
rect 348572 66780 348628 66836
rect 345212 28476 345268 28532
rect 348572 59612 348628 59668
rect 340172 26684 340228 26740
rect 337036 26460 337092 26516
rect 350252 180460 350308 180516
rect 368172 215068 368228 215124
rect 366716 213612 366772 213668
rect 376236 213724 376292 213780
rect 370860 212828 370916 212884
rect 378252 212828 378308 212884
rect 352156 201180 352212 201236
rect 351932 195356 351988 195412
rect 351820 184940 351876 184996
rect 352044 187740 352100 187796
rect 350588 171612 350644 171668
rect 351932 178780 351988 178836
rect 352156 182700 352212 182756
rect 393932 173964 393988 174020
rect 352156 171724 352212 171780
rect 368844 171724 368900 171780
rect 375564 171612 375620 171668
rect 376908 171164 376964 171220
rect 373548 169372 373604 169428
rect 352044 169036 352100 169092
rect 406588 219324 406644 219380
rect 398972 171164 399028 171220
rect 412412 218540 412468 218596
rect 427532 218092 427588 218148
rect 429212 221900 429268 221956
rect 434140 219324 434196 219380
rect 429212 217756 429268 217812
rect 433468 218092 433524 218148
rect 430780 213500 430836 213556
rect 473116 230860 473172 230916
rect 440972 230300 441028 230356
rect 437612 217644 437668 217700
rect 439516 217756 439572 217812
rect 436156 217420 436212 217476
rect 437500 215516 437556 215572
rect 464492 226380 464548 226436
rect 440972 217756 441028 217812
rect 461132 225820 461188 225876
rect 436828 213276 436884 213332
rect 414092 171612 414148 171668
rect 432124 171612 432180 171668
rect 412412 171052 412468 171108
rect 393932 169372 393988 169428
rect 438508 171164 438564 171220
rect 461132 171164 461188 171220
rect 440300 171052 440356 171108
rect 464492 171052 464548 171108
rect 474684 227500 474740 227556
rect 473116 170940 473172 170996
rect 474572 174300 474628 174356
rect 439068 169260 439124 169316
rect 472892 169820 472948 169876
rect 432348 169148 432404 169204
rect 377580 169036 377636 169092
rect 414092 165900 414148 165956
rect 398972 164220 399028 164276
rect 351932 152012 351988 152068
rect 372652 152348 372708 152404
rect 376908 152124 376964 152180
rect 372652 147084 372708 147140
rect 372876 150332 372932 150388
rect 352716 144844 352772 144900
rect 352716 143724 352772 143780
rect 350588 143164 350644 143220
rect 350364 137900 350420 137956
rect 369516 143164 369572 143220
rect 351932 143052 351988 143108
rect 351036 141708 351092 141764
rect 351036 138460 351092 138516
rect 350588 126140 350644 126196
rect 352156 142940 352212 142996
rect 352044 142268 352100 142324
rect 368172 142268 368228 142324
rect 372204 142828 372260 142884
rect 374220 147084 374276 147140
rect 373548 143052 373604 143108
rect 393148 142828 393204 142884
rect 375564 142156 375620 142212
rect 376236 142044 376292 142100
rect 393148 139580 393204 139636
rect 352156 135660 352212 135716
rect 352044 128604 352100 128660
rect 351932 124460 351988 124516
rect 352044 114380 352100 114436
rect 350364 100492 350420 100548
rect 350476 107660 350532 107716
rect 350252 99036 350308 99092
rect 350476 96908 350532 96964
rect 351932 102620 351988 102676
rect 349356 57036 349412 57092
rect 350252 96460 350308 96516
rect 350252 29708 350308 29764
rect 352044 88172 352100 88228
rect 352492 107100 352548 107156
rect 351932 29484 351988 29540
rect 352044 78540 352100 78596
rect 410732 163660 410788 163716
rect 398972 101724 399028 101780
rect 407372 160860 407428 160916
rect 407372 100828 407428 100884
rect 368172 100716 368228 100772
rect 368844 100716 368900 100772
rect 376908 100604 376964 100660
rect 412412 161420 412468 161476
rect 410844 159180 410900 159236
rect 410844 101948 410900 102004
rect 413980 144956 414036 145012
rect 413980 140700 414036 140756
rect 412412 101836 412468 101892
rect 414092 101612 414148 101668
rect 414204 159740 414260 159796
rect 410732 100604 410788 100660
rect 437612 146972 437668 147028
rect 437612 145292 437668 145348
rect 435484 144956 435540 145012
rect 434812 144844 434868 144900
rect 432796 144732 432852 144788
rect 435036 143052 435092 143108
rect 435036 142380 435092 142436
rect 437500 144508 437556 144564
rect 438172 142940 438228 142996
rect 444220 100828 444276 100884
rect 472892 100828 472948 100884
rect 422044 100716 422100 100772
rect 429436 100716 429492 100772
rect 434140 100716 434196 100772
rect 438844 100716 438900 100772
rect 435484 100604 435540 100660
rect 501564 217756 501620 217812
rect 500892 217644 500948 217700
rect 475468 215516 475524 215572
rect 496860 215516 496916 215572
rect 495516 215404 495572 215460
rect 492156 215292 492212 215348
rect 555548 240044 555604 240100
rect 553532 239820 553588 239876
rect 562268 241836 562324 241892
rect 560252 239932 560308 239988
rect 557564 239596 557620 239652
rect 536732 236012 536788 236068
rect 503132 217532 503188 217588
rect 523292 234780 523348 234836
rect 496188 213388 496244 213444
rect 475468 211036 475524 211092
rect 493500 171276 493556 171332
rect 494172 170940 494228 170996
rect 474684 170828 474740 170884
rect 533484 232652 533540 232708
rect 523292 171276 523348 171332
rect 533372 172172 533428 172228
rect 496188 171164 496244 171220
rect 495516 171052 495572 171108
rect 494844 170828 494900 170884
rect 493500 167132 493556 167188
rect 475468 144508 475524 144564
rect 494172 158844 494228 158900
rect 497532 144508 497588 144564
rect 500892 143052 500948 143108
rect 498204 142828 498260 142884
rect 492828 141708 492884 141764
rect 475468 140476 475524 140532
rect 498876 100940 498932 100996
rect 499548 100828 499604 100884
rect 474572 100604 474628 100660
rect 495516 100604 495572 100660
rect 420028 100492 420084 100548
rect 420476 100492 420532 100548
rect 414204 100268 414260 100324
rect 428764 100268 428820 100324
rect 492828 98812 492884 98868
rect 500892 100492 500948 100548
rect 533484 169260 533540 169316
rect 560364 235900 560420 235956
rect 560252 227612 560308 227668
rect 555548 217532 555604 217588
rect 539196 215292 539252 215348
rect 558908 215292 558964 215348
rect 564284 222572 564340 222628
rect 560364 216636 560420 216692
rect 562268 216636 562324 216692
rect 562940 215628 562996 215684
rect 563612 215180 563668 215236
rect 557564 212940 557620 212996
rect 539196 210812 539252 210868
rect 580636 403564 580692 403620
rect 582092 569884 582148 569940
rect 587132 569212 587188 569268
rect 582204 567420 582260 567476
rect 582204 548940 582260 548996
rect 585452 567308 585508 567364
rect 585452 469868 585508 469924
rect 582092 271404 582148 271460
rect 580412 192108 580468 192164
rect 536732 169148 536788 169204
rect 556108 169484 556164 169540
rect 571676 171276 571732 171332
rect 562828 169596 562884 169652
rect 559580 169372 559636 169428
rect 558236 169260 558292 169316
rect 554876 169148 554932 169204
rect 556892 162092 556948 162148
rect 556220 152012 556276 152068
rect 536732 150780 536788 150836
rect 557564 160412 557620 160468
rect 561596 145740 561652 145796
rect 560252 145292 560308 145348
rect 587244 566972 587300 567028
rect 590604 569324 590660 569380
rect 590604 535836 590660 535892
rect 590716 528108 590772 528164
rect 590604 521612 590660 521668
rect 590716 496300 590772 496356
rect 590604 390572 590660 390628
rect 590492 350924 590548 350980
rect 587244 324492 587300 324548
rect 587132 113036 587188 113092
rect 536732 101052 536788 101108
rect 556892 101052 556948 101108
rect 533372 98812 533428 98868
rect 564284 99036 564340 99092
rect 558908 98924 558964 98980
rect 556220 98812 556276 98868
rect 494172 98700 494228 98756
rect 430108 98588 430164 98644
rect 438172 96908 438228 96964
rect 355292 94780 355348 94836
rect 355292 79996 355348 80052
rect 372204 89964 372260 90020
rect 352492 78428 352548 78484
rect 371308 78316 371364 78372
rect 371308 75068 371364 75124
rect 352716 74060 352772 74116
rect 352268 70588 352324 70644
rect 359548 73948 359604 74004
rect 368844 73948 368900 74004
rect 432572 89180 432628 89236
rect 403228 87500 403284 87556
rect 393932 85820 393988 85876
rect 375452 84700 375508 84756
rect 375452 74844 375508 74900
rect 379596 79996 379652 80052
rect 376908 74172 376964 74228
rect 372876 74060 372932 74116
rect 403228 81452 403284 81508
rect 407372 81900 407428 81956
rect 404796 80780 404852 80836
rect 404796 78316 404852 78372
rect 404012 77980 404068 78036
rect 393932 74956 393988 75012
rect 402332 76300 402388 76356
rect 402332 74732 402388 74788
rect 359548 70700 359604 70756
rect 371196 70700 371252 70756
rect 377580 70588 377636 70644
rect 352716 68460 352772 68516
rect 352268 66892 352324 66948
rect 372204 29708 372260 29764
rect 370860 29596 370916 29652
rect 404012 29596 404068 29652
rect 377580 29372 377636 29428
rect 432124 74732 432180 74788
rect 436156 78428 436212 78484
rect 432572 74732 432628 74788
rect 433468 75068 433524 75124
rect 556892 96684 556948 96740
rect 504252 94892 504308 94948
rect 461916 91420 461972 91476
rect 461916 84924 461972 84980
rect 464492 90300 464548 90356
rect 461132 83580 461188 83636
rect 407372 29372 407428 29428
rect 414092 31052 414148 31108
rect 352044 26572 352100 26628
rect 348572 26348 348628 26404
rect 376908 26460 376964 26516
rect 434812 29596 434868 29652
rect 434140 29484 434196 29540
rect 436828 29260 436884 29316
rect 432796 26572 432852 26628
rect 414092 26460 414148 26516
rect 461132 29260 461188 29316
rect 494844 88172 494900 88228
rect 492156 81340 492212 81396
rect 494172 78316 494228 78372
rect 498204 86492 498260 86548
rect 497532 74956 497588 75012
rect 499772 85260 499828 85316
rect 501564 74844 501620 74900
rect 499772 74620 499828 74676
rect 500892 74620 500948 74676
rect 554204 93212 554260 93268
rect 560252 84924 560308 84980
rect 557564 78092 557620 78148
rect 560924 81452 560980 81508
rect 562268 74732 562324 74788
rect 498204 29372 498260 29428
rect 499548 29260 499604 29316
rect 495516 28476 495572 28532
rect 494172 26796 494228 26852
rect 492156 26684 492212 26740
rect 464492 26572 464548 26628
rect 562268 26572 562324 26628
rect 438844 26460 438900 26516
rect 374892 26348 374948 26404
rect 329644 24332 329700 24388
rect 4172 22876 4228 22932
rect 11564 5068 11620 5124
<< metal3 >>
rect 407362 591276 407372 591332
rect 407428 591276 408268 591332
rect 408324 591276 408334 591332
rect 165666 590604 165676 590660
rect 165732 590604 284732 590660
rect 284788 590604 284798 590660
rect 288082 590604 288092 590660
rect 288148 590604 364028 590660
rect 364084 590604 364094 590660
rect 33282 590492 33292 590548
rect 33348 590492 46172 590548
rect 46228 590492 46238 590548
rect 99474 590492 99484 590548
rect 99540 590492 287084 590548
rect 287140 590492 287150 590548
rect 289762 590492 289772 590548
rect 289828 590492 297836 590548
rect 297892 590492 297902 590548
rect 303202 590492 303212 590548
rect 303268 590492 430220 590548
rect 430276 590492 430286 590548
rect 432562 590492 432572 590548
rect 432628 590492 496412 590548
rect 496468 590492 496478 590548
rect 499762 590492 499772 590548
rect 499828 590492 562604 590548
rect 562660 590492 562670 590548
rect 595560 588644 597000 588840
rect 304994 588588 305004 588644
rect 305060 588616 597000 588644
rect 305060 588588 595672 588616
rect -960 587160 480 587384
rect 46162 583772 46172 583828
rect 46228 583772 288204 583828
rect 288260 583772 288270 583828
rect 307234 583772 307244 583828
rect 307300 583772 474348 583828
rect 474404 583772 474414 583828
rect 209570 582204 209580 582260
rect 209636 582204 311724 582260
rect 311780 582204 311790 582260
rect 279234 582092 279244 582148
rect 279300 582092 499772 582148
rect 499828 582092 499838 582148
rect 309474 578844 309484 578900
rect 309540 578844 341964 578900
rect 342020 578844 342030 578900
rect 10994 578732 11004 578788
rect 11060 578732 315084 578788
rect 315140 578732 315150 578788
rect 231634 577164 231644 577220
rect 231700 577164 284844 577220
rect 284900 577164 284910 577220
rect 308354 577164 308364 577220
rect 308420 577164 407372 577220
rect 407428 577164 407438 577220
rect 280354 577052 280364 577108
rect 280420 577052 432572 577108
rect 432628 577052 432638 577108
rect 283714 576156 283724 576212
rect 283780 576156 289772 576212
rect 289828 576156 289838 576212
rect 281474 575484 281484 575540
rect 281540 575484 303212 575540
rect 303268 575484 303278 575540
rect 595560 575428 597000 575624
rect 278114 575372 278124 575428
rect 278180 575400 597000 575428
rect 278180 575372 595672 575400
rect 284722 574476 284732 574532
rect 284788 574476 285964 574532
rect 286020 574476 286030 574532
rect 282594 574364 282604 574420
rect 282660 574364 288092 574420
rect 288148 574364 288158 574420
rect 275762 574028 275772 574084
rect 275828 574028 310604 574084
rect 310660 574028 310670 574084
rect 143378 573916 143388 573972
rect 143444 573916 312844 573972
rect 312900 573916 312910 573972
rect 306114 573804 306124 573860
rect 306180 573804 540540 573860
rect 540596 573804 540606 573860
rect 77298 573692 77308 573748
rect 77364 573692 313964 573748
rect 314020 573692 314030 573748
rect -960 573076 480 573272
rect -960 573048 76412 573076
rect 392 573020 76412 573048
rect 76468 573020 76478 573076
rect 266242 572348 266252 572404
rect 266308 572348 328524 572404
rect 328580 572348 328590 572404
rect 299394 572236 299404 572292
rect 299460 572236 335244 572292
rect 335300 572236 335310 572292
rect 249442 572124 249452 572180
rect 249508 572124 329644 572180
rect 329700 572124 329710 572180
rect 296482 572012 296492 572068
rect 296548 572012 325164 572068
rect 325220 572012 325230 572068
rect 40226 571900 40236 571956
rect 40292 571900 257852 571956
rect 257908 571900 257918 571956
rect 276994 571900 277004 571956
rect 277060 571900 315756 571956
rect 315812 571900 315822 571956
rect 338706 571900 338716 571956
rect 338772 571900 557564 571956
rect 557620 571900 557630 571956
rect 160178 571788 160188 571844
rect 160244 571788 187292 571844
rect 187348 571788 187358 571844
rect 224802 571788 224812 571844
rect 224868 571788 256172 571844
rect 256228 571788 256238 571844
rect 268146 571788 268156 571844
rect 268212 571788 317324 571844
rect 317380 571788 317390 571844
rect 336914 571788 336924 571844
rect 336980 571788 433468 571844
rect 433524 571788 433534 571844
rect 474674 571788 474684 571844
rect 474740 571788 501564 571844
rect 501620 571788 501630 571844
rect 44258 571676 44268 571732
rect 44324 571676 62972 571732
rect 63028 571676 63038 571732
rect 170258 571676 170268 571732
rect 170324 571676 247996 571732
rect 248052 571676 248062 571732
rect 267922 571676 267932 571732
rect 267988 571676 327404 571732
rect 327460 571676 327470 571732
rect 337138 571676 337148 571732
rect 337204 571676 438172 571732
rect 438228 571676 438238 571732
rect 464482 571676 464492 571732
rect 464548 571676 498204 571732
rect 498260 571676 498270 571732
rect 45602 571564 45612 571620
rect 45668 571564 69692 571620
rect 69748 571564 69758 571620
rect 104850 571564 104860 571620
rect 104916 571564 130172 571620
rect 130228 571564 130238 571620
rect 164210 571564 164220 571620
rect 164276 571564 247772 571620
rect 247828 571564 247838 571620
rect 275874 571564 275884 571620
rect 275940 571564 335468 571620
rect 335524 571564 335534 571620
rect 351922 571564 351932 571620
rect 351988 571564 496188 571620
rect 496244 571564 496254 571620
rect 533362 571564 533372 571620
rect 533428 571564 558236 571620
rect 558292 571564 558302 571620
rect 41570 571452 41580 571508
rect 41636 571452 73052 571508
rect 73108 571452 73118 571508
rect 100146 571452 100156 571508
rect 100212 571452 136892 571508
rect 136948 571452 136958 571508
rect 160850 571452 160860 571508
rect 160916 571452 263004 571508
rect 263060 571452 263070 571508
rect 266466 571452 266476 571508
rect 266532 571452 326284 571508
rect 326340 571452 326350 571508
rect 338482 571452 338492 571508
rect 338548 571452 374220 571508
rect 374276 571452 374286 571508
rect 407362 571452 407372 571508
rect 407428 571452 558908 571508
rect 558964 571452 558974 571508
rect 38882 571340 38892 571396
rect 38948 571340 78092 571396
rect 78148 571340 78158 571396
rect 107538 571340 107548 571396
rect 107604 571340 261212 571396
rect 261268 571340 261278 571396
rect 341842 571340 341852 571396
rect 341908 571340 555548 571396
rect 555604 571340 555614 571396
rect 46946 571228 46956 571284
rect 47012 571228 63196 571284
rect 63252 571228 63262 571284
rect 224130 571228 224140 571284
rect 224196 571228 249676 571284
rect 249732 571228 249742 571284
rect 319106 571228 319116 571284
rect 319172 571228 324044 571284
rect 324100 571228 324110 571284
rect 330726 571228 330764 571284
rect 330820 571228 330830 571284
rect 350242 571228 350252 571284
rect 350308 571228 370860 571284
rect 370916 571228 370926 571284
rect 412402 571228 412412 571284
rect 412468 571228 430780 571284
rect 430836 571228 430846 571284
rect 536722 571228 536732 571284
rect 536788 571228 554204 571284
rect 554260 571228 554270 571284
rect 4274 570668 4284 570724
rect 4340 570668 296492 570724
rect 296548 570668 296558 570724
rect 298274 570668 298284 570724
rect 298340 570668 590492 570724
rect 590548 570668 590558 570724
rect 273634 570556 273644 570612
rect 273700 570556 580636 570612
rect 580692 570556 580702 570612
rect 40226 570444 40236 570500
rect 40292 570444 264572 570500
rect 264628 570444 264638 570500
rect 294914 570444 294924 570500
rect 294980 570444 336812 570500
rect 336868 570444 336878 570500
rect 292674 570332 292684 570388
rect 292740 570332 340172 570388
rect 340228 570332 340238 570388
rect 274754 570220 274764 570276
rect 274820 570220 333676 570276
rect 333732 570220 333742 570276
rect 269154 570108 269164 570164
rect 269220 570108 333452 570164
rect 333508 570108 333518 570164
rect 345202 570108 345212 570164
rect 345268 570108 380268 570164
rect 380324 570108 380334 570164
rect 412514 570108 412524 570164
rect 412580 570108 435484 570164
rect 435540 570108 435550 570164
rect 169586 569996 169596 570052
rect 169652 569996 187404 570052
rect 187460 569996 187470 570052
rect 231522 569996 231532 570052
rect 231588 569996 259756 570052
rect 259812 569996 259822 570052
rect 315746 569996 315756 570052
rect 315812 569996 317996 570052
rect 318052 569996 318062 570052
rect 471202 569996 471212 570052
rect 471268 569996 500892 570052
rect 500948 569996 500958 570052
rect 162866 569884 162876 569940
rect 162932 569884 192332 569940
rect 192388 569884 192398 569940
rect 228162 569884 228172 569940
rect 228228 569884 257964 569940
rect 258020 569884 258030 569940
rect 296034 569884 296044 569940
rect 296100 569884 582092 569940
rect 582148 569884 582158 569940
rect 168914 569772 168924 569828
rect 168980 569772 199052 569828
rect 199108 569772 199118 569828
rect 226146 569772 226156 569828
rect 226212 569772 263116 569828
rect 263172 569772 263182 569828
rect 290406 569772 290444 569828
rect 290500 569772 290510 569828
rect 293794 569772 293804 569828
rect 293860 569772 580412 569828
rect 580468 569772 580478 569828
rect 46722 569660 46732 569716
rect 46788 569660 125132 569716
rect 125188 569660 125198 569716
rect 166450 569660 166460 569716
rect 166516 569660 259532 569716
rect 259588 569660 259598 569716
rect 296930 569660 296940 569716
rect 296996 569660 474572 569716
rect 474628 569660 474638 569716
rect 476242 569660 476252 569716
rect 476308 569660 492268 569716
rect 492324 569660 492334 569716
rect 36866 569548 36876 569604
rect 36932 569548 252812 569604
rect 252868 569548 252878 569604
rect 303622 569548 303660 569604
rect 303716 569548 303726 569604
rect 315746 569548 315756 569604
rect 315812 569548 315868 569604
rect 315924 569548 315934 569604
rect 350354 569548 350364 569604
rect 350420 569548 374892 569604
rect 374948 569548 374958 569604
rect 414082 569548 414092 569604
rect 414148 569548 435708 569604
rect 435764 569548 435774 569604
rect 474786 569548 474796 569604
rect 474852 569548 494844 569604
rect 494900 569548 494910 569604
rect 266578 569436 266588 569492
rect 266644 569436 322924 569492
rect 322980 569436 322990 569492
rect 4498 569324 4508 569380
rect 4564 569324 317772 569380
rect 317828 569324 317838 569380
rect 317986 569324 317996 569380
rect 318052 569324 590604 569380
rect 590660 569324 590670 569380
rect 291554 569212 291564 569268
rect 291620 569212 587132 569268
rect 587188 569212 587198 569268
rect 15922 569100 15932 569156
rect 15988 569100 320684 569156
rect 320740 569100 320750 569156
rect 7634 568988 7644 569044
rect 7700 568988 321804 569044
rect 321860 568988 321870 569044
rect 352034 568988 352044 569044
rect 352100 568988 372204 569044
rect 372260 568988 372270 569044
rect 230850 568876 230860 568932
rect 230916 568876 254492 568932
rect 254548 568876 254558 568932
rect 270246 568876 270284 568932
rect 270340 568876 270350 568932
rect 271366 568876 271404 568932
rect 271460 568876 271470 568932
rect 272486 568876 272524 568932
rect 272580 568876 272590 568932
rect 289286 568876 289324 568932
rect 289380 568876 289390 568932
rect 300486 568876 300524 568932
rect 300580 568876 300590 568932
rect 301606 568876 301644 568932
rect 301700 568876 301710 568932
rect 302726 568876 302764 568932
rect 302820 568876 302830 568932
rect 314132 568876 319564 568932
rect 319620 568876 319630 568932
rect 345314 568876 345324 568932
rect 345380 568876 377580 568932
rect 377636 568876 377646 568932
rect 314132 568820 314188 568876
rect 290612 568764 314188 568820
rect 290612 568708 290668 568764
rect 266354 568652 266364 568708
rect 266420 568652 290668 568708
rect 302754 568652 302764 568708
rect 302820 568652 302830 568708
rect 302764 568596 302820 568652
rect 302764 568540 335132 568596
rect 335188 568540 335198 568596
rect 270274 567756 270284 567812
rect 270340 567756 333564 567812
rect 333620 567756 333630 567812
rect 300514 567644 300524 567700
rect 300580 567644 400652 567700
rect 400708 567644 400718 567700
rect 272514 567532 272524 567588
rect 272580 567532 393932 567588
rect 393988 567532 393998 567588
rect 303650 567420 303660 567476
rect 303716 567420 582204 567476
rect 582260 567420 582270 567476
rect 301634 567308 301644 567364
rect 301700 567308 585452 567364
rect 585508 567308 585518 567364
rect 4162 567196 4172 567252
rect 4228 567196 315756 567252
rect 315812 567196 315822 567252
rect 4386 567084 4396 567140
rect 4452 567084 319116 567140
rect 319172 567084 319182 567140
rect 271394 566972 271404 567028
rect 271460 566972 587244 567028
rect 587300 566972 587310 567028
rect 141026 563948 141036 564004
rect 141092 563948 144088 564004
rect 579880 563948 583212 564004
rect 583268 563948 583278 564004
rect 595560 562184 597000 562408
rect 392 559160 4172 559188
rect -960 559132 4172 559160
rect 4228 559132 4238 559188
rect -960 558936 480 559132
rect 141026 556108 141036 556164
rect 141092 556108 141932 556164
rect 141988 556108 141998 556164
rect 18386 555884 18396 555940
rect 18452 555884 20104 555940
rect 141026 555884 141036 555940
rect 141092 555912 144088 555940
rect 141092 555884 144116 555912
rect 144060 555268 144116 555884
rect 80098 555212 80108 555268
rect 80164 555212 82040 555268
rect 144050 555212 144060 555268
rect 144116 555212 144126 555268
rect 349346 555212 349356 555268
rect 349412 555212 352716 555268
rect 352772 555212 352782 555268
rect 473666 555212 473676 555268
rect 473732 555240 476056 555268
rect 473732 555212 476084 555240
rect 414642 555100 414652 555156
rect 414708 555100 414718 555156
rect 80434 554540 80444 554596
rect 80500 554540 82040 554596
rect 123928 554540 126924 554596
rect 126980 554540 126990 554596
rect 201618 554540 201628 554596
rect 201684 554540 206136 554596
rect 414652 554568 414708 555100
rect 476028 554820 476084 555212
rect 476018 554764 476028 554820
rect 476084 554764 476094 554820
rect 18358 554428 18396 554484
rect 18452 554428 18462 554484
rect 82674 553868 82684 553924
rect 82740 553868 82750 553924
rect 247912 553868 252812 553924
rect 252868 553868 252878 553924
rect 347778 553868 347788 553924
rect 347844 553868 352072 553924
rect 410946 553868 410956 553924
rect 411012 553868 414120 553924
rect 473442 553868 473452 553924
rect 473508 553868 476056 553924
rect 519026 553868 519036 553924
rect 519092 553868 538104 553924
rect 18274 553196 18284 553252
rect 18340 553196 20104 553252
rect 340274 553196 340284 553252
rect 340340 553196 352072 553252
rect 410722 553196 410732 553252
rect 410788 553196 414120 553252
rect 455896 553196 458780 553252
rect 458836 553196 458846 553252
rect 472882 553196 472892 553252
rect 472948 553196 476056 553252
rect 579880 553196 583436 553252
rect 583492 553196 583502 553252
rect 61880 552524 65100 552580
rect 65156 552524 65166 552580
rect 123928 552524 127260 552580
rect 127316 552524 127326 552580
rect 204866 552524 204876 552580
rect 204932 552524 206136 552580
rect 247912 552524 261324 552580
rect 261380 552524 261390 552580
rect 473218 552524 473228 552580
rect 473284 552524 476056 552580
rect 535490 552524 535500 552580
rect 535556 552524 538104 552580
rect 579880 552524 583324 552580
rect 583380 552524 583390 552580
rect 18386 551852 18396 551908
rect 18452 551852 20104 551908
rect 141026 551852 141036 551908
rect 141092 551852 144088 551908
rect 203186 551852 203196 551908
rect 203252 551852 206136 551908
rect 393960 551852 396844 551908
rect 396900 551852 396910 551908
rect 455896 551852 458668 551908
rect 458724 551852 458734 551908
rect 517944 551852 521276 551908
rect 521332 551852 521342 551908
rect 341954 551628 341964 551684
rect 342020 551628 347788 551684
rect 347844 551628 347854 551684
rect 579852 551348 579908 551880
rect 579852 551292 582484 551348
rect 80322 551180 80332 551236
rect 80388 551180 82040 551236
rect 140914 551180 140924 551236
rect 140980 551180 144088 551236
rect 185864 551180 189084 551236
rect 189140 551180 189150 551236
rect 247912 551180 262892 551236
rect 262948 551180 262958 551236
rect 348562 551180 348572 551236
rect 348628 551180 352072 551236
rect 393960 551180 394828 551236
rect 394884 551180 394894 551236
rect 455896 551180 459004 551236
rect 459060 551180 459070 551236
rect 517916 551124 517972 551208
rect 535266 551180 535276 551236
rect 535332 551180 538104 551236
rect 579618 551180 579628 551236
rect 579684 551180 579694 551236
rect 582428 551124 582484 551292
rect 517916 551068 518252 551124
rect 518308 551068 518318 551124
rect 582418 551068 582428 551124
rect 582484 551068 582494 551124
rect 206108 550004 206164 550536
rect 345202 550508 345212 550564
rect 345268 550508 352072 550564
rect 473106 550508 473116 550564
rect 473172 550508 476056 550564
rect 205762 549948 205772 550004
rect 205828 549948 206164 550004
rect 61880 549836 74732 549892
rect 74788 549836 74798 549892
rect 185864 549836 188972 549892
rect 189028 549836 189038 549892
rect 348674 549836 348684 549892
rect 348740 549836 352072 549892
rect 410834 549836 410844 549892
rect 410900 549836 414120 549892
rect 517944 549836 520940 549892
rect 520996 549836 521006 549892
rect 534258 549836 534268 549892
rect 534324 549836 538104 549892
rect 61880 549164 74844 549220
rect 74900 549164 74910 549220
rect 82002 549164 82012 549220
rect 82068 549164 82078 549220
rect 338482 549164 338492 549220
rect 338548 549164 352072 549220
rect 455896 549164 458892 549220
rect 458948 549164 458958 549220
rect 595560 548996 597000 549192
rect 582194 548940 582204 548996
rect 582260 548968 597000 548996
rect 582260 548940 595672 548968
rect 61880 548492 64652 548548
rect 64708 548492 64718 548548
rect 123928 548492 143612 548548
rect 143668 548492 143678 548548
rect 185864 548492 189196 548548
rect 189252 548492 189262 548548
rect 247912 548492 257852 548548
rect 257908 548492 257918 548548
rect 402322 548492 402332 548548
rect 402388 548492 414120 548548
rect 455896 548492 456988 548548
rect 457044 548492 457054 548548
rect 461122 548492 461132 548548
rect 461188 548492 473228 548548
rect 473284 548492 473294 548548
rect 476028 547876 476084 548520
rect 523282 548492 523292 548548
rect 523348 548492 534268 548548
rect 534324 548492 534334 548548
rect 579880 548492 583100 548548
rect 583156 548492 583166 548548
rect 123928 547820 126812 547876
rect 126868 547820 126878 547876
rect 247912 547820 264572 547876
rect 264628 547820 264638 547876
rect 473218 547820 473228 547876
rect 473284 547820 476084 547876
rect 535154 547820 535164 547876
rect 535220 547820 538104 547876
rect 456082 547708 456092 547764
rect 456148 547708 458668 547764
rect 458724 547708 458734 547764
rect 82226 547148 82236 547204
rect 82292 547148 82302 547204
rect 123928 547148 127036 547204
rect 127092 547148 127102 547204
rect 247912 547148 251916 547204
rect 251972 547148 251982 547204
rect 393362 547148 393372 547204
rect 393428 547148 393438 547204
rect 517944 547148 521052 547204
rect 521108 547148 521118 547204
rect 535042 547148 535052 547204
rect 535108 547148 538104 547204
rect 82114 546476 82124 546532
rect 82180 546476 82190 546532
rect 123928 546476 142044 546532
rect 142100 546476 142110 546532
rect 411058 546476 411068 546532
rect 411124 546476 414120 546532
rect 455896 546476 458668 546532
rect 458724 546476 458734 546532
rect 472994 546476 473004 546532
rect 473060 546476 476056 546532
rect 517944 546476 519260 546532
rect 519316 546476 519326 546532
rect 579880 546476 581308 546532
rect 581364 546476 581374 546532
rect 141026 546028 141036 546084
rect 141092 546028 143724 546084
rect 143780 546028 143790 546084
rect 457762 546028 457772 546084
rect 457828 546028 458780 546084
rect 458836 546028 458846 546084
rect 20066 545804 20076 545860
rect 20132 545804 20142 545860
rect 61880 545804 64764 545860
rect 64820 545804 64830 545860
rect 123928 545804 127148 545860
rect 127204 545804 127214 545860
rect 185864 545804 197372 545860
rect 197428 545804 197438 545860
rect 247912 545804 254492 545860
rect 254548 545804 254558 545860
rect 473330 545804 473340 545860
rect 473396 545804 476056 545860
rect 18162 545132 18172 545188
rect 18228 545132 20104 545188
rect 123928 545132 138572 545188
rect 138628 545132 138638 545188
rect 140802 545132 140812 545188
rect 140868 545132 144088 545188
rect 185864 545132 189420 545188
rect 189476 545132 189486 545188
rect 247912 545132 259980 545188
rect 260036 545132 260046 545188
rect 341842 545132 341852 545188
rect 341908 545132 352072 545188
rect 455896 545132 458780 545188
rect 458836 545132 458846 545188
rect 517916 545076 517972 545832
rect 579880 545804 581420 545860
rect 581476 545804 581486 545860
rect -960 544824 480 545048
rect 517916 545020 519988 545076
rect 519932 544852 519988 545020
rect 519922 544796 519932 544852
rect 519988 544796 519998 544852
rect 61880 544460 64988 544516
rect 65044 544460 65054 544516
rect 80210 544460 80220 544516
rect 80276 544460 82040 544516
rect 141026 544460 141036 544516
rect 141092 544460 144088 544516
rect 203074 544460 203084 544516
rect 203140 544460 206136 544516
rect 247912 544460 256284 544516
rect 256340 544460 256350 544516
rect 393960 544460 394940 544516
rect 394996 544460 395006 544516
rect 517944 544460 519148 544516
rect 519204 544460 519214 544516
rect 203186 544348 203196 544404
rect 203252 544348 204092 544404
rect 204148 544348 204158 544404
rect 18050 543788 18060 543844
rect 18116 543788 20104 543844
rect 203074 543788 203084 543844
rect 203140 543788 206136 543844
rect 247912 543788 261212 543844
rect 261268 543788 261278 543844
rect 340162 543788 340172 543844
rect 340228 543788 352072 543844
rect 393932 543284 393988 543816
rect 398962 543788 398972 543844
rect 399028 543788 414120 543844
rect 535378 543788 535388 543844
rect 535444 543788 538104 543844
rect 393932 543228 395612 543284
rect 395668 543228 395678 543284
rect 142706 543116 142716 543172
rect 142772 543116 144088 543172
rect 393932 542724 393988 543144
rect 517944 543116 520828 543172
rect 520884 543116 520894 543172
rect 393932 542668 396732 542724
rect 396788 542668 396798 542724
rect 393960 542444 396620 542500
rect 396676 542444 396686 542500
rect 455298 542444 455308 542500
rect 455364 542444 455374 542500
rect 517944 541772 521164 541828
rect 521220 541772 521230 541828
rect 61880 538412 64876 538468
rect 64932 538412 64942 538468
rect 464482 536732 464492 536788
rect 464548 536732 473452 536788
rect 473508 536732 473518 536788
rect 595560 535892 597000 535976
rect 590594 535836 590604 535892
rect 590660 535836 597000 535892
rect 595560 535752 597000 535836
rect 252802 533372 252812 533428
rect 252868 533372 263900 533428
rect 263956 533372 263966 533428
rect 519026 533372 519036 533428
rect 519092 533372 535388 533428
rect 535444 533372 535454 533428
rect 254482 531580 254492 531636
rect 254548 531580 268072 531636
rect 331912 531580 337596 531636
rect 337652 531580 337662 531636
rect 263778 531020 263788 531076
rect 263844 531020 268072 531076
rect 331912 531020 341852 531076
rect 341908 531020 341918 531076
rect -960 530740 480 530936
rect -960 530712 12572 530740
rect 392 530684 12572 530712
rect 12628 530684 12638 530740
rect 263778 530460 263788 530516
rect 263844 530460 268072 530516
rect 331912 530460 523292 530516
rect 523348 530460 523358 530516
rect 140802 530236 140812 530292
rect 140868 530236 205996 530292
rect 206052 530236 206062 530292
rect 65090 530124 65100 530180
rect 65156 530124 259532 530180
rect 259588 530124 259598 530180
rect 456866 530124 456876 530180
rect 456932 530124 583212 530180
rect 583268 530124 583278 530180
rect 18162 530012 18172 530068
rect 18228 530012 256172 530068
rect 256228 530012 256238 530068
rect 335906 530012 335916 530068
rect 335972 530012 533372 530068
rect 533428 530012 533438 530068
rect 205762 529900 205772 529956
rect 205828 529900 268072 529956
rect 331912 529900 582428 529956
rect 582484 529900 582494 529956
rect 263890 529340 263900 529396
rect 263956 529340 268072 529396
rect 331912 529340 539196 529396
rect 539252 529340 539262 529396
rect 140914 529116 140924 529172
rect 140980 529116 146076 529172
rect 146132 529116 146142 529172
rect 261314 528780 261324 528836
rect 261380 528780 268072 528836
rect 331884 528388 331940 528808
rect 335244 528444 344428 528500
rect 331884 528332 332668 528388
rect 332724 528332 332734 528388
rect 18050 528220 18060 528276
rect 18116 528220 261548 528276
rect 261604 528220 261614 528276
rect 63186 528108 63196 528164
rect 63252 528108 265132 528164
rect 265188 528108 265198 528164
rect 80210 527996 80220 528052
rect 80276 527996 252812 528052
rect 252868 527996 252878 528052
rect 268044 527940 268100 528248
rect 331884 528052 331940 528248
rect 335244 528164 335300 528444
rect 335458 528332 335468 528388
rect 335524 528332 339332 528388
rect 332332 528108 335300 528164
rect 339276 528164 339332 528332
rect 344372 528276 344428 528444
rect 344372 528220 519036 528276
rect 519092 528220 519102 528276
rect 339276 528108 590716 528164
rect 590772 528108 590782 528164
rect 332332 528052 332388 528108
rect 331884 527996 332388 528052
rect 354386 527996 354396 528052
rect 354452 527996 535500 528052
rect 535556 527996 535566 528052
rect 227490 527884 227500 527940
rect 227556 527884 268100 527940
rect 357746 527884 357756 527940
rect 357812 527884 520828 527940
rect 520884 527884 520894 527940
rect 224018 527772 224028 527828
rect 224084 527772 263788 527828
rect 263844 527772 263854 527828
rect 332658 527772 332668 527828
rect 332724 527772 357868 527828
rect 357924 527772 357934 527828
rect 539186 527772 539196 527828
rect 539252 527772 556892 527828
rect 556948 527772 556958 527828
rect 224802 527660 224812 527716
rect 224868 527660 268072 527716
rect 331912 527660 559580 527716
rect 559636 527660 559646 527716
rect 357858 527436 357868 527492
rect 357924 527436 557564 527492
rect 557620 527436 557630 527492
rect 259746 527100 259756 527156
rect 259812 527100 268072 527156
rect 331912 527100 335916 527156
rect 335972 527100 335982 527156
rect 127250 526652 127260 526708
rect 127316 526652 249452 526708
rect 249508 526652 249518 526708
rect 335906 526652 335916 526708
rect 335972 526652 536732 526708
rect 536788 526652 536798 526708
rect 259970 526540 259980 526596
rect 260036 526540 268072 526596
rect 331912 526540 456876 526596
rect 456932 526540 456942 526596
rect 224690 525980 224700 526036
rect 224756 525980 268072 526036
rect 331912 525980 354396 526036
rect 354452 525980 354462 526036
rect 337586 525756 337596 525812
rect 337652 525756 554876 525812
rect 554932 525756 554942 525812
rect 249666 525420 249676 525476
rect 249732 525420 268072 525476
rect 331912 525420 562268 525476
rect 562324 525420 562334 525476
rect 230178 525308 230188 525364
rect 230244 525308 244412 525364
rect 244468 525308 244478 525364
rect 164210 525196 164220 525252
rect 164276 525196 253036 525252
rect 253092 525196 253102 525252
rect 98802 525084 98812 525140
rect 98868 525084 258188 525140
rect 258244 525084 258254 525140
rect 36194 524972 36204 525028
rect 36260 524972 249900 525028
rect 249956 524972 249966 525028
rect 256274 524860 256284 524916
rect 256340 524860 268072 524916
rect 331912 524860 335916 524916
rect 335972 524860 335982 524916
rect 251906 524300 251916 524356
rect 251972 524300 268072 524356
rect 331912 524300 564284 524356
rect 564340 524300 564350 524356
rect 162866 523740 162876 523796
rect 162932 523740 268072 523796
rect 331912 523740 521164 523796
rect 521220 523740 521230 523796
rect 168914 523628 168924 523684
rect 168980 523628 198156 523684
rect 198212 523628 198222 523684
rect 100146 523516 100156 523572
rect 100212 523516 170492 523572
rect 170548 523516 170558 523572
rect 203074 523516 203084 523572
rect 203140 523516 246092 523572
rect 246148 523516 246158 523572
rect 372082 523516 372092 523572
rect 372148 523516 376908 523572
rect 376964 523516 376974 523572
rect 40226 523404 40236 523460
rect 40292 523404 249676 523460
rect 249732 523404 249742 523460
rect 368722 523404 368732 523460
rect 368788 523404 377580 523460
rect 377636 523404 377646 523460
rect 379698 523404 379708 523460
rect 379764 523404 498204 523460
rect 498260 523404 498270 523460
rect 4162 523292 4172 523348
rect 4228 523292 249452 523348
rect 249508 523292 249518 523348
rect 348786 523292 348796 523348
rect 348852 523292 473340 523348
rect 473396 523292 473406 523348
rect 475458 523292 475468 523348
rect 475524 523292 499548 523348
rect 499604 523292 499614 523348
rect 146066 523180 146076 523236
rect 146132 523180 268072 523236
rect 331912 523180 471212 523236
rect 471268 523180 471278 523236
rect 197362 522620 197372 522676
rect 197428 522620 268072 522676
rect 331912 522620 518252 522676
rect 518308 522620 518318 522676
rect 595560 522536 597000 522760
rect 189186 522060 189196 522116
rect 189252 522060 268072 522116
rect 331912 522060 357756 522116
rect 357812 522060 357822 522116
rect 106866 521948 106876 522004
rect 106932 521948 188076 522004
rect 188132 521948 188142 522004
rect 351922 521948 351932 522004
rect 351988 521948 396732 522004
rect 396788 521948 396798 522004
rect 107538 521836 107548 521892
rect 107604 521836 192444 521892
rect 192500 521836 192510 521892
rect 340274 521836 340284 521892
rect 340340 521836 435484 521892
rect 435540 521836 435550 521892
rect 126914 521724 126924 521780
rect 126980 521724 256508 521780
rect 256564 521724 256574 521780
rect 356178 521724 356188 521780
rect 356244 521724 494844 521780
rect 494900 521724 494910 521780
rect 18274 521612 18284 521668
rect 18340 521612 256284 521668
rect 256340 521612 256350 521668
rect 335234 521612 335244 521668
rect 335300 521612 590604 521668
rect 590660 521612 590670 521668
rect 189410 521500 189420 521556
rect 189476 521500 268072 521556
rect 331912 521500 474684 521556
rect 474740 521500 474750 521556
rect 205986 520940 205996 520996
rect 206052 520940 268072 520996
rect 331912 520940 476140 520996
rect 476196 520940 476206 520996
rect 142706 520380 142716 520436
rect 142772 520380 268072 520436
rect 331912 520380 379708 520436
rect 379764 520380 379774 520436
rect 355282 520156 355292 520212
rect 355348 520156 411068 520212
rect 411124 520156 411134 520212
rect 80434 520044 80444 520100
rect 80500 520044 247772 520100
rect 247828 520044 247838 520100
rect 380482 520044 380492 520100
rect 380548 520044 459004 520100
rect 459060 520044 459070 520100
rect 82226 519932 82236 519988
rect 82292 519932 263788 519988
rect 263844 519932 263854 519988
rect 336802 519932 336812 519988
rect 336868 519932 521052 519988
rect 521108 519932 521118 519988
rect 143714 519820 143724 519876
rect 143780 519820 268072 519876
rect 331912 519820 475468 519876
rect 475524 519820 475534 519876
rect 192322 519260 192332 519316
rect 192388 519260 268072 519316
rect 331912 519260 519260 519316
rect 519316 519260 519326 519316
rect 168242 518700 168252 518756
rect 168308 518700 268072 518756
rect 331912 518700 461132 518756
rect 461188 518700 461198 518756
rect 40898 518476 40908 518532
rect 40964 518476 157052 518532
rect 157108 518476 157118 518532
rect 82114 518364 82124 518420
rect 82180 518364 264908 518420
rect 264964 518364 264974 518420
rect 334450 518364 334460 518420
rect 334516 518364 440188 518420
rect 440244 518364 440254 518420
rect 80322 518252 80332 518308
rect 80388 518252 263116 518308
rect 263172 518252 263182 518308
rect 353602 518252 353612 518308
rect 353668 518252 583324 518308
rect 583380 518252 583390 518308
rect 187394 518140 187404 518196
rect 187460 518140 268072 518196
rect 331912 518140 519932 518196
rect 519988 518140 519998 518196
rect 199042 517580 199052 517636
rect 199108 517580 268072 517636
rect 331912 517580 474796 517636
rect 474852 517580 474862 517636
rect 198146 517020 198156 517076
rect 198212 517020 268072 517076
rect 331912 517020 464492 517076
rect 464548 517020 464558 517076
rect 381378 516908 381388 516964
rect 381444 516908 436828 516964
rect 436884 516908 436894 516964
rect -960 516628 480 516824
rect 342626 516796 342636 516852
rect 342692 516796 428092 516852
rect 428148 516796 428158 516852
rect 103506 516684 103516 516740
rect 103572 516684 259756 516740
rect 259812 516684 259822 516740
rect 353714 516684 353724 516740
rect 353780 516684 535276 516740
rect 535332 516684 535342 516740
rect -960 516600 268156 516628
rect 392 516572 268156 516600
rect 268212 516572 268222 516628
rect 335234 516572 335244 516628
rect 335300 516572 519148 516628
rect 519204 516572 519214 516628
rect 141922 516460 141932 516516
rect 141988 516460 268072 516516
rect 331912 516460 356188 516516
rect 356244 516460 356254 516516
rect 82002 515900 82012 515956
rect 82068 515900 268072 515956
rect 331912 515900 398972 515956
rect 399028 515900 399038 515956
rect 188066 515340 188076 515396
rect 188132 515340 268072 515396
rect 331912 515340 381388 515396
rect 381444 515340 381454 515396
rect 80098 514892 80108 514948
rect 80164 514892 257964 514948
rect 258020 514892 258030 514948
rect 335234 514892 335244 514948
rect 335300 514892 464492 514948
rect 464548 514892 464558 514948
rect 142034 514780 142044 514836
rect 142100 514780 268072 514836
rect 331912 514780 456988 514836
rect 457044 514780 457054 514836
rect 263778 514220 263788 514276
rect 263844 514220 268072 514276
rect 331912 514220 334460 514276
rect 334516 514220 334526 514276
rect 127026 513660 127036 513716
rect 127092 513660 268072 513716
rect 331912 513660 380492 513716
rect 380548 513660 380558 513716
rect 160178 513324 160188 513380
rect 160244 513324 249564 513380
rect 249620 513324 249630 513380
rect 342066 513324 342076 513380
rect 342132 513324 473228 513380
rect 473284 513324 473294 513380
rect 130162 513212 130172 513268
rect 130228 513212 264684 513268
rect 264740 513212 264750 513268
rect 345538 513212 345548 513268
rect 345604 513212 583100 513268
rect 583156 513212 583166 513268
rect 126802 513100 126812 513156
rect 126868 513100 268072 513156
rect 331912 513100 456092 513156
rect 456148 513100 456158 513156
rect 264898 512540 264908 512596
rect 264964 512540 268072 512596
rect 331912 512540 457772 512596
rect 457828 512540 457838 512596
rect 99474 511980 99484 512036
rect 99540 511980 268072 512036
rect 331912 511980 355292 512036
rect 355348 511980 355358 512036
rect 334450 511868 334460 511924
rect 334516 511868 402332 511924
rect 402388 511868 402398 511924
rect 339266 511756 339276 511812
rect 339332 511756 442204 511812
rect 442260 511756 442270 511812
rect 141026 511644 141036 511700
rect 141092 511644 247884 511700
rect 247940 511644 247950 511700
rect 354386 511644 354396 511700
rect 354452 511644 458892 511700
rect 458948 511644 458958 511700
rect 38210 511532 38220 511588
rect 38276 511532 261660 511588
rect 261716 511532 261726 511588
rect 340386 511532 340396 511588
rect 340452 511532 520940 511588
rect 520996 511532 521006 511588
rect 102834 511420 102844 511476
rect 102900 511420 268072 511476
rect 331912 511420 342636 511476
rect 342692 511420 342702 511476
rect 127138 510860 127148 510916
rect 127204 510860 268072 510916
rect 331912 510860 412524 510916
rect 412580 510860 412590 510916
rect 170482 510300 170492 510356
rect 170548 510300 268072 510356
rect 331912 510300 354396 510356
rect 354452 510300 354462 510356
rect 334338 510188 334348 510244
rect 334404 510188 394828 510244
rect 394884 510188 394894 510244
rect 335458 510076 335468 510132
rect 335524 510076 455308 510132
rect 455364 510076 455374 510132
rect 102162 509964 102172 510020
rect 102228 509964 254604 510020
rect 254660 509964 254670 510020
rect 345314 509964 345324 510020
rect 345380 509964 473116 510020
rect 473172 509964 473182 510020
rect 74834 509852 74844 509908
rect 74900 509852 263788 509908
rect 263844 509852 263854 509908
rect 353826 509852 353836 509908
rect 353892 509852 535164 509908
rect 535220 509852 535230 509908
rect 192434 509740 192444 509796
rect 192500 509740 268072 509796
rect 331912 509740 334460 509796
rect 334516 509740 334526 509796
rect 595560 509348 597000 509544
rect 335122 509292 335132 509348
rect 335188 509320 597000 509348
rect 335188 509292 595672 509320
rect 138562 509180 138572 509236
rect 138628 509180 268072 509236
rect 331912 509180 414092 509236
rect 414148 509180 414158 509236
rect 143602 508620 143612 508676
rect 143668 508620 268072 508676
rect 331912 508620 339276 508676
rect 339332 508620 339342 508676
rect 342178 508284 342188 508340
rect 342244 508284 410844 508340
rect 410900 508284 410910 508340
rect 167570 508172 167580 508228
rect 167636 508172 261772 508228
rect 261828 508172 261838 508228
rect 350578 508172 350588 508228
rect 350644 508172 493500 508228
rect 493556 508172 493566 508228
rect 263778 508060 263788 508116
rect 263844 508060 268072 508116
rect 331912 508060 341964 508116
rect 342020 508060 342030 508116
rect 261538 507500 261548 507556
rect 261604 507500 268072 507556
rect 331912 507500 334348 507556
rect 334404 507500 334414 507556
rect 342066 507052 342076 507108
rect 342132 507052 370188 507108
rect 370244 507052 370254 507108
rect 264562 506940 264572 506996
rect 264628 506940 268072 506996
rect 331912 506940 345324 506996
rect 345380 506940 345390 506996
rect 350578 506828 350588 506884
rect 350644 506828 410956 506884
rect 411012 506828 411022 506884
rect 189074 506716 189084 506772
rect 189140 506716 247996 506772
rect 248052 506716 248062 506772
rect 352146 506716 352156 506772
rect 352212 506716 458668 506772
rect 458724 506716 458734 506772
rect 73042 506604 73052 506660
rect 73108 506604 264796 506660
rect 264852 506604 264862 506660
rect 335122 506604 335132 506660
rect 335188 506604 393372 506660
rect 393428 506604 393438 506660
rect 402322 506604 402332 506660
rect 402388 506604 535052 506660
rect 535108 506604 535118 506660
rect 62962 506492 62972 506548
rect 63028 506492 265020 506548
rect 265076 506492 265086 506548
rect 338706 506492 338716 506548
rect 338772 506492 521276 506548
rect 521332 506492 521342 506548
rect 64642 506380 64652 506436
rect 64708 506380 268072 506436
rect 331912 506380 350364 506436
rect 350420 506380 350430 506436
rect 69682 505820 69692 505876
rect 69748 505820 268072 505876
rect 331912 505820 372092 505876
rect 372148 505820 372158 505876
rect 337698 505372 337708 505428
rect 337764 505372 396620 505428
rect 396676 505372 396686 505428
rect 64754 505260 64764 505316
rect 64820 505260 268072 505316
rect 331912 505260 368732 505316
rect 368788 505260 368798 505316
rect 348898 505148 348908 505204
rect 348964 505148 410732 505204
rect 410788 505148 410798 505204
rect 338594 505036 338604 505092
rect 338660 505036 458780 505092
rect 458836 505036 458846 505092
rect 169586 504924 169596 504980
rect 169652 504924 254716 504980
rect 254772 504924 254782 504980
rect 352258 504924 352268 504980
rect 352324 504924 473004 504980
rect 473060 504924 473070 504980
rect 74722 504812 74732 504868
rect 74788 504812 264684 504868
rect 264740 504812 264750 504868
rect 335346 504812 335356 504868
rect 335412 504812 394940 504868
rect 394996 504812 395006 504868
rect 395154 504812 395164 504868
rect 395220 504812 563612 504868
rect 563668 504812 563678 504868
rect 64978 504700 64988 504756
rect 65044 504700 268072 504756
rect 331912 504700 340284 504756
rect 340340 504700 340350 504756
rect 18386 504140 18396 504196
rect 18452 504140 268072 504196
rect 331912 504140 352044 504196
rect 352100 504140 352110 504196
rect 337250 503692 337260 503748
rect 337316 503692 372204 503748
rect 372260 503692 372270 503748
rect 125122 503580 125132 503636
rect 125188 503580 268072 503636
rect 331912 503580 338492 503636
rect 338548 503580 338558 503636
rect 335906 503468 335916 503524
rect 335972 503468 348684 503524
rect 348740 503468 348750 503524
rect 349010 503468 349020 503524
rect 349076 503468 396844 503524
rect 396900 503468 396910 503524
rect 346882 503356 346892 503412
rect 346948 503356 430108 503412
rect 430164 503356 430174 503412
rect 188962 503244 188972 503300
rect 189028 503244 251916 503300
rect 251972 503244 251982 503300
rect 345538 503244 345548 503300
rect 345604 503244 434812 503300
rect 434868 503244 434878 503300
rect 78082 503132 78092 503188
rect 78148 503132 264908 503188
rect 264964 503132 264974 503188
rect 337698 503132 337708 503188
rect 337764 503132 376236 503188
rect 376292 503132 376302 503188
rect 393922 503132 393932 503188
rect 393988 503132 583436 503188
rect 583492 503132 583502 503188
rect 39554 503020 39564 503076
rect 39620 503020 268072 503076
rect 331912 503020 395612 503076
rect 395668 503020 395678 503076
rect -960 502488 480 502712
rect 64866 502460 64876 502516
rect 64932 502460 268072 502516
rect 331912 502460 345212 502516
rect 345268 502460 345278 502516
rect 20066 501900 20076 501956
rect 20132 501900 268072 501956
rect 331912 501900 335916 501956
rect 335972 501900 335982 501956
rect 335122 501564 335132 501620
rect 335188 501564 412412 501620
rect 412468 501564 412478 501620
rect 203186 501452 203196 501508
rect 203252 501452 246876 501508
rect 246932 501452 246942 501508
rect 344082 501452 344092 501508
rect 344148 501452 472892 501508
rect 472948 501452 472958 501508
rect 157042 501340 157052 501396
rect 157108 501340 268072 501396
rect 331912 501340 337708 501396
rect 337764 501340 337774 501396
rect 98802 501116 98812 501172
rect 98868 501116 125132 501172
rect 125188 501116 125198 501172
rect 100146 501004 100156 501060
rect 100212 501004 130172 501060
rect 130228 501004 130238 501060
rect 166226 501004 166236 501060
rect 166292 501004 187404 501060
rect 187460 501004 187470 501060
rect 345202 501004 345212 501060
rect 345268 501004 370188 501060
rect 370244 501004 370254 501060
rect 398962 501004 398972 501060
rect 399028 501004 436156 501060
rect 436212 501004 436222 501060
rect 536722 501004 536732 501060
rect 536788 501004 558908 501060
rect 558964 501004 558974 501060
rect 36194 500892 36204 500948
rect 36260 500892 62972 500948
rect 63028 500892 63038 500948
rect 100818 500892 100828 500948
rect 100884 500892 135212 500948
rect 135268 500892 135278 500948
rect 170930 500892 170940 500948
rect 170996 500892 195692 500948
rect 195748 500892 195758 500948
rect 230178 500892 230188 500948
rect 230244 500892 259868 500948
rect 259924 500892 259934 500948
rect 350354 500892 350364 500948
rect 350420 500892 438844 500948
rect 438900 500892 438910 500948
rect 476242 500892 476252 500948
rect 476308 500892 498876 500948
rect 498932 500892 498942 500948
rect 530002 500892 530012 500948
rect 530068 500892 562268 500948
rect 562324 500892 562334 500948
rect 40898 500780 40908 500836
rect 40964 500780 74732 500836
rect 74788 500780 74798 500836
rect 104850 500780 104860 500836
rect 104916 500780 200732 500836
rect 200788 500780 200798 500836
rect 226146 500780 226156 500836
rect 226212 500780 261324 500836
rect 261380 500780 261390 500836
rect 265122 500780 265132 500836
rect 265188 500780 268072 500836
rect 331912 500780 337708 500836
rect 337764 500780 337774 500836
rect 338594 500780 338604 500836
rect 338660 500780 372876 500836
rect 372932 500780 372942 500836
rect 407474 500780 407484 500836
rect 407540 500780 558236 500836
rect 558292 500780 558302 500836
rect 36866 500668 36876 500724
rect 36932 500668 262892 500724
rect 262948 500668 262958 500724
rect 340386 500668 340396 500724
rect 340452 500668 554876 500724
rect 554932 500668 554942 500724
rect 257842 500220 257852 500276
rect 257908 500220 268072 500276
rect 331912 500220 581420 500276
rect 581476 500220 581486 500276
rect 262882 500108 262892 500164
rect 262948 500108 263900 500164
rect 263956 500108 263966 500164
rect 264562 499660 264572 499716
rect 264628 499660 268072 499716
rect 331912 499660 353836 499716
rect 353892 499660 353902 499716
rect 222786 499548 222796 499604
rect 222852 499548 252924 499604
rect 252980 499548 252990 499604
rect 348562 499548 348572 499604
rect 348628 499548 562940 499604
rect 562996 499548 563006 499604
rect 164210 499436 164220 499492
rect 164276 499436 263228 499492
rect 263284 499436 263294 499492
rect 345314 499436 345324 499492
rect 345380 499436 368172 499492
rect 368228 499436 368238 499492
rect 155474 499324 155484 499380
rect 155540 499324 261548 499380
rect 261604 499324 261614 499380
rect 338818 499324 338828 499380
rect 338884 499324 369516 499380
rect 369572 499324 369582 499380
rect 46946 499212 46956 499268
rect 47012 499212 197372 499268
rect 197428 499212 197438 499268
rect 231522 499212 231532 499268
rect 231588 499212 258300 499268
rect 258356 499212 258366 499268
rect 341842 499212 341852 499268
rect 341908 499212 374220 499268
rect 374276 499212 374286 499268
rect 412402 499212 412412 499268
rect 412468 499212 432796 499268
rect 432852 499212 432862 499268
rect 464482 499212 464492 499268
rect 464548 499212 493500 499268
rect 493556 499212 493566 499268
rect 104178 499100 104188 499156
rect 104244 499100 259644 499156
rect 259700 499100 259710 499156
rect 261202 499100 261212 499156
rect 261268 499100 268072 499156
rect 331912 499100 345548 499156
rect 345604 499100 345614 499156
rect 352146 499100 352156 499156
rect 352212 499100 556220 499156
rect 556276 499100 556286 499156
rect 37538 498988 37548 499044
rect 37604 498988 205772 499044
rect 205828 498988 205838 499044
rect 232194 498988 232204 499044
rect 232260 498988 253148 499044
rect 253204 498988 253214 499044
rect 350466 498988 350476 499044
rect 350532 498988 368844 499044
rect 368900 498988 368910 499044
rect 244402 498540 244412 498596
rect 244468 498540 268072 498596
rect 331912 498540 581308 498596
rect 581364 498540 581374 498596
rect 162866 498428 162876 498484
rect 162932 498428 249452 498484
rect 249508 498428 249518 498484
rect 103506 498316 103516 498372
rect 103572 498316 258076 498372
rect 258132 498316 258142 498372
rect 166898 498204 166908 498260
rect 166964 498204 187516 498260
rect 187572 498204 187582 498260
rect 337026 498204 337036 498260
rect 337092 498204 434812 498260
rect 434868 498204 434878 498260
rect 187282 498092 187292 498148
rect 187348 498092 264572 498148
rect 264628 498092 264638 498148
rect 345426 498092 345436 498148
rect 345492 498092 492828 498148
rect 492884 498092 492894 498148
rect 164882 497980 164892 498036
rect 164948 497980 192332 498036
rect 192388 497980 192398 498036
rect 263890 497980 263900 498036
rect 263956 497980 268072 498036
rect 331912 497980 579628 498036
rect 579684 497980 579694 498036
rect 178994 497868 179004 497924
rect 179060 497868 256284 497924
rect 256340 497868 256350 497924
rect 352034 497868 352044 497924
rect 352100 497868 376236 497924
rect 376292 497868 376302 497924
rect 474674 497868 474684 497924
rect 474740 497868 494172 497924
rect 494228 497868 494238 497924
rect 533362 497868 533372 497924
rect 533428 497868 555548 497924
rect 555604 497868 555614 497924
rect 43586 497756 43596 497812
rect 43652 497756 199052 497812
rect 199108 497756 199118 497812
rect 226818 497756 226828 497812
rect 226884 497756 261436 497812
rect 261492 497756 261502 497812
rect 341954 497756 341964 497812
rect 342020 497756 564284 497812
rect 564340 497756 564350 497812
rect 246866 497532 246876 497588
rect 246932 497532 268100 497588
rect 268044 497448 268100 497532
rect 331912 497420 353724 497476
rect 353780 497420 353790 497476
rect 204082 496860 204092 496916
rect 204148 496860 268072 496916
rect 331912 496860 402332 496916
rect 402388 496860 402398 496916
rect 136882 496412 136892 496468
rect 136948 496412 265132 496468
rect 265188 496412 265198 496468
rect 263106 496300 263116 496356
rect 263172 496300 268072 496356
rect 331912 496300 395164 496356
rect 395220 496300 395230 496356
rect 590706 496300 590716 496356
rect 590772 496328 595672 496356
rect 590772 496300 597000 496328
rect 595560 496104 597000 496300
rect 254482 495740 254492 495796
rect 254548 495740 268072 495796
rect 331912 495740 393932 495796
rect 393988 495740 393998 495796
rect 246082 495180 246092 495236
rect 246148 495180 268072 495236
rect 331912 495180 407372 495236
rect 407428 495180 407438 495236
rect 349412 494956 353612 495012
rect 353668 494956 353678 495012
rect 256162 494620 256172 494676
rect 256228 494620 268072 494676
rect 331912 494620 338716 494676
rect 338772 494620 338782 494676
rect 349412 494452 349468 494956
rect 331884 494396 349468 494452
rect 257954 494060 257964 494116
rect 258020 494060 268072 494116
rect 331884 494088 331940 494396
rect 249554 493500 249564 493556
rect 249620 493500 268072 493556
rect 331912 493500 348796 493556
rect 348852 493500 348862 493556
rect 123928 493388 143612 493444
rect 143668 493388 143678 493444
rect 455896 493388 459228 493444
rect 459284 493388 459294 493444
rect 247874 492940 247884 492996
rect 247940 492940 268072 492996
rect 331912 492940 336812 492996
rect 336868 492940 336878 492996
rect 61880 492716 69692 492772
rect 69748 492716 69758 492772
rect 140914 492716 140924 492772
rect 140980 492716 144088 492772
rect 261762 492380 261772 492436
rect 261828 492380 268072 492436
rect 331912 492380 350588 492436
rect 350644 492380 350654 492436
rect 253026 491820 253036 491876
rect 253092 491820 268072 491876
rect 331912 491820 345324 491876
rect 345380 491820 345390 491876
rect 259522 491260 259532 491316
rect 259588 491260 268072 491316
rect 331912 491260 352268 491316
rect 352324 491260 352334 491316
rect 247986 490700 247996 490756
rect 248052 490700 268072 490756
rect 331912 490700 335244 490756
rect 335300 490700 335310 490756
rect 254706 490140 254716 490196
rect 254772 490140 268072 490196
rect 331912 490140 342076 490196
rect 342132 490140 342142 490196
rect 247986 489580 247996 489636
rect 248052 489580 268072 489636
rect 331912 489580 344092 489636
rect 344148 489580 344158 489636
rect 247762 489020 247772 489076
rect 247828 489020 268072 489076
rect 331912 489020 351932 489076
rect 351988 489020 351998 489076
rect -960 488404 480 488600
rect 264562 488460 264572 488516
rect 264628 488460 268072 488516
rect 331912 488460 335244 488516
rect 335300 488460 335310 488516
rect -960 488376 14252 488404
rect 392 488348 14252 488376
rect 14308 488348 14318 488404
rect 335570 488012 335580 488068
rect 335636 488012 345212 488068
rect 345268 488012 345278 488068
rect 262994 487900 263004 487956
rect 263060 487900 268072 487956
rect 331912 487900 340396 487956
rect 340452 487900 340462 487956
rect 251906 487340 251916 487396
rect 251972 487340 268072 487396
rect 331912 487340 338716 487396
rect 338772 487340 338782 487396
rect 247762 486780 247772 486836
rect 247828 486780 268072 486836
rect 331912 486780 346892 486836
rect 346948 486780 346958 486836
rect 257954 486220 257964 486276
rect 258020 486220 268072 486276
rect 331912 486220 337148 486276
rect 337204 486220 337214 486276
rect 265122 485660 265132 485716
rect 265188 485660 268072 485716
rect 331912 485660 348908 485716
rect 348964 485660 348974 485716
rect 256498 485100 256508 485156
rect 256564 485100 268072 485156
rect 331912 485100 336924 485156
rect 336980 485100 336990 485156
rect 335570 484652 335580 484708
rect 335636 484652 350252 484708
rect 350308 484652 350318 484708
rect 534258 484652 534268 484708
rect 534324 484652 538104 484708
rect 249442 484540 249452 484596
rect 249508 484540 268072 484596
rect 331912 484540 350588 484596
rect 350644 484540 350654 484596
rect 476018 484316 476028 484372
rect 476084 484316 476094 484372
rect 476028 484036 476084 484316
rect 18358 483980 18396 484036
rect 18452 483980 20076 484036
rect 20132 483980 20142 484036
rect 141036 483980 144088 484036
rect 259746 483980 259756 484036
rect 259812 483980 268072 484036
rect 331912 483980 342188 484036
rect 342244 483980 342254 484036
rect 473666 483980 473676 484036
rect 473732 484008 476084 484036
rect 473732 483980 476056 484008
rect 141036 483812 141092 483980
rect 141026 483756 141036 483812
rect 141092 483756 141102 483812
rect 335794 483756 335804 483812
rect 335860 483756 340172 483812
rect 340228 483756 340238 483812
rect 252802 483420 252812 483476
rect 252868 483420 268072 483476
rect 331912 483420 335468 483476
rect 335524 483420 335534 483476
rect 61880 483308 64764 483364
rect 64820 483308 64830 483364
rect 82674 483308 82684 483364
rect 82740 483308 82750 483364
rect 201618 483308 201628 483364
rect 201684 483308 206136 483364
rect 349346 483308 349356 483364
rect 349412 483308 352716 483364
rect 352772 483308 352782 483364
rect 393960 483308 396844 483364
rect 396900 483308 396910 483364
rect 455896 483308 458668 483364
rect 458724 483308 458734 483364
rect 517944 483308 519148 483364
rect 519204 483308 519214 483364
rect 254594 482860 254604 482916
rect 254660 482860 268072 482916
rect 331912 482860 335132 482916
rect 335188 482860 335198 482916
rect 595560 482888 597000 483112
rect 123928 482636 126028 482692
rect 185864 482636 189084 482692
rect 189140 482636 189150 482692
rect 125972 482132 126028 482636
rect 206556 482356 206612 482664
rect 247912 482636 259644 482692
rect 259700 482636 259710 482692
rect 393960 482636 396732 482692
rect 396788 482636 396798 482692
rect 410834 482636 410844 482692
rect 410900 482636 414120 482692
rect 455896 482636 458780 482692
rect 458836 482636 458846 482692
rect 472098 482636 472108 482692
rect 472164 482636 476056 482692
rect 206556 482300 206668 482356
rect 206724 482300 206734 482356
rect 261202 482300 261212 482356
rect 261268 482300 268072 482356
rect 331912 482300 345548 482356
rect 345604 482300 345614 482356
rect 125972 482076 136892 482132
rect 136948 482076 136958 482132
rect 82226 481964 82236 482020
rect 82292 481964 82302 482020
rect 123928 481964 127596 482020
rect 127652 481964 127662 482020
rect 247912 481964 262892 482020
rect 262948 481964 262958 482020
rect 411170 481964 411180 482020
rect 411236 481964 414120 482020
rect 455896 481964 456988 482020
rect 457044 481964 457054 482020
rect 472210 481964 472220 482020
rect 472276 481964 476056 482020
rect 517916 481908 517972 482664
rect 579880 482636 581308 482692
rect 581364 482636 581374 482692
rect 534258 481964 534268 482020
rect 534324 481964 538104 482020
rect 517916 481852 518252 481908
rect 518308 481852 518318 481908
rect 263106 481740 263116 481796
rect 263172 481740 268072 481796
rect 331912 481740 352156 481796
rect 352212 481740 352222 481796
rect 461122 481404 461132 481460
rect 461188 481404 472108 481460
rect 472164 481404 472174 481460
rect 61880 481292 64876 481348
rect 64932 481292 64942 481348
rect 123928 481292 142044 481348
rect 142100 481292 142110 481348
rect 203186 481292 203196 481348
rect 203252 481292 206136 481348
rect 410946 481292 410956 481348
rect 411012 481292 414120 481348
rect 455896 481292 459004 481348
rect 459060 481292 459070 481348
rect 462802 481292 462812 481348
rect 462868 481292 476056 481348
rect 535042 481292 535052 481348
rect 535108 481292 538104 481348
rect 258178 481180 258188 481236
rect 258244 481180 268072 481236
rect 331912 481180 338604 481236
rect 338660 481180 338670 481236
rect 414642 481068 414652 481124
rect 414708 481068 414718 481124
rect 18162 480620 18172 480676
rect 18228 480620 20104 480676
rect 141026 480620 141036 480676
rect 141092 480620 144088 480676
rect 247912 480620 261324 480676
rect 261380 480620 261390 480676
rect 264674 480620 264684 480676
rect 264740 480620 268072 480676
rect 331912 480620 340284 480676
rect 340340 480620 340350 480676
rect 414652 480648 414708 481068
rect 455896 480620 458892 480676
rect 458948 480620 458958 480676
rect 579880 480620 583324 480676
rect 583380 480620 583390 480676
rect 127586 480396 127596 480452
rect 127652 480396 130172 480452
rect 130228 480396 130238 480452
rect 140914 480396 140924 480452
rect 140980 480396 143724 480452
rect 143780 480396 143790 480452
rect 257842 480396 257852 480452
rect 257908 480396 263900 480452
rect 263956 480396 263966 480452
rect 265010 480060 265020 480116
rect 265076 480060 268072 480116
rect 331912 480060 349020 480116
rect 349076 480060 349086 480116
rect 18274 479948 18284 480004
rect 18340 479948 20104 480004
rect 123928 479948 133532 480004
rect 133588 479948 133598 480004
rect 185864 479948 197372 480004
rect 197428 479948 197438 480004
rect 348786 479948 348796 480004
rect 348852 479948 352072 480004
rect 393960 479948 394828 480004
rect 394884 479948 394894 480004
rect 455298 479948 455308 480004
rect 455364 479948 455374 480004
rect 472882 479948 472892 480004
rect 472948 479948 476056 480004
rect 517458 479948 517468 480004
rect 517524 479948 517534 480004
rect 249890 479612 249900 479668
rect 249956 479612 263788 479668
rect 263844 479612 263854 479668
rect 523282 479612 523292 479668
rect 523348 479612 534268 479668
rect 534324 479612 534334 479668
rect 259522 479500 259532 479556
rect 259588 479500 268072 479556
rect 331912 479500 348572 479556
rect 348628 479500 348638 479556
rect 61880 479276 65100 479332
rect 65156 479276 65166 479332
rect 80546 479276 80556 479332
rect 80612 479276 82040 479332
rect 185864 479276 204204 479332
rect 204260 479276 204270 479332
rect 206556 478660 206612 479304
rect 348674 479276 348684 479332
rect 348740 479276 352072 479332
rect 393960 479276 394940 479332
rect 394996 479276 395006 479332
rect 455410 479276 455420 479332
rect 455476 479276 455486 479332
rect 473106 479276 473116 479332
rect 473172 479276 476056 479332
rect 517944 479276 521164 479332
rect 521220 479276 521230 479332
rect 579880 479276 581420 479332
rect 581476 479276 581486 479332
rect 264674 478940 264684 478996
rect 264740 478940 268072 478996
rect 331912 478940 342076 478996
rect 342132 478940 342142 478996
rect 61880 478604 73164 478660
rect 73220 478604 73230 478660
rect 80322 478604 80332 478660
rect 80388 478604 82040 478660
rect 123928 478604 127596 478660
rect 127652 478604 127662 478660
rect 185864 478604 188972 478660
rect 189028 478604 189038 478660
rect 206546 478604 206556 478660
rect 206612 478604 206622 478660
rect 247912 478604 251020 478660
rect 251076 478604 251086 478660
rect 342066 478604 342076 478660
rect 342132 478604 352072 478660
rect 393960 478604 396508 478660
rect 396564 478604 396574 478660
rect 455896 478604 459116 478660
rect 459172 478604 459182 478660
rect 579880 478604 582988 478660
rect 583044 478604 583054 478660
rect 263778 478380 263788 478436
rect 263844 478380 268072 478436
rect 331912 478380 341852 478436
rect 341908 478380 341918 478436
rect 579618 478380 579628 478436
rect 579684 478380 579694 478436
rect 185864 477932 194908 477988
rect 194964 477932 194974 477988
rect 247912 477932 250908 477988
rect 250964 477932 250974 477988
rect 404002 477932 404012 477988
rect 404068 477932 414120 477988
rect 455896 477932 457324 477988
rect 457380 477932 457390 477988
rect 467842 477932 467852 477988
rect 467908 477932 476056 477988
rect 579628 477960 579684 478380
rect 256162 477820 256172 477876
rect 256228 477820 268072 477876
rect 331912 477820 337260 477876
rect 337316 477820 337326 477876
rect 17938 477260 17948 477316
rect 18004 477260 20104 477316
rect 140914 477260 140924 477316
rect 140980 477260 144088 477316
rect 247912 477260 252812 477316
rect 252868 477260 252878 477316
rect 261650 477260 261660 477316
rect 261716 477260 268072 477316
rect 331912 477260 335356 477316
rect 335412 477260 335422 477316
rect 517944 477260 518532 477316
rect 518476 477204 518532 477260
rect 518466 477148 518476 477204
rect 518532 477148 518542 477204
rect 249666 476700 249676 476756
rect 249732 476700 268072 476756
rect 331912 476700 338492 476756
rect 338548 476700 338558 476756
rect 61880 476588 78316 476644
rect 78372 476588 78382 476644
rect 80434 476588 80444 476644
rect 80500 476588 82040 476644
rect 123928 476588 135212 476644
rect 135268 476588 135278 476644
rect 140802 476588 140812 476644
rect 140868 476588 144088 476644
rect 247912 476588 259532 476644
rect 259588 476588 259598 476644
rect 340162 476588 340172 476644
rect 340228 476588 352072 476644
rect 393960 476588 396620 476644
rect 396676 476588 396686 476644
rect 517944 476588 519260 476644
rect 519316 476588 519326 476644
rect 127586 476252 127596 476308
rect 127652 476252 138572 476308
rect 138628 476252 138638 476308
rect 251010 476252 251020 476308
rect 251076 476252 264572 476308
rect 264628 476252 264638 476308
rect 252802 476140 252812 476196
rect 252868 476140 268072 476196
rect 331912 476140 335132 476196
rect 335188 476140 335198 476196
rect 18050 475916 18060 475972
rect 18116 475916 20104 475972
rect 61880 475916 64652 475972
rect 64708 475916 64718 475972
rect 185864 475916 189532 475972
rect 189588 475916 189598 475972
rect 247912 475916 261212 475972
rect 261268 475916 261278 475972
rect 393362 475916 393372 475972
rect 393428 475916 393438 475972
rect 400642 475916 400652 475972
rect 400708 475916 414120 475972
rect 455522 475916 455532 475972
rect 455588 475916 455598 475972
rect 517944 475916 520940 475972
rect 520996 475916 521006 475972
rect 579394 475916 579404 475972
rect 579460 475916 579470 475972
rect 264898 475580 264908 475636
rect 264964 475580 268072 475636
rect 331912 475580 335580 475636
rect 335636 475580 335646 475636
rect 141026 475468 141036 475524
rect 141092 475468 141932 475524
rect 141988 475468 141998 475524
rect 335346 475468 335356 475524
rect 335412 475468 339388 475524
rect 339444 475468 339454 475524
rect 457762 475468 457772 475524
rect 457828 475468 458668 475524
rect 458724 475468 458734 475524
rect 395602 475356 395612 475412
rect 395668 475356 396844 475412
rect 396900 475356 396910 475412
rect 20066 475244 20076 475300
rect 20132 475244 20142 475300
rect 256274 475020 256284 475076
rect 256340 475020 268072 475076
rect 331912 475020 351932 475076
rect 351988 475020 351998 475076
rect 455868 474852 455924 475272
rect 250898 474796 250908 474852
rect 250964 474796 256508 474852
rect 256564 474796 256574 474852
rect 455868 474796 456148 474852
rect 123928 474572 126812 474628
rect 126868 474572 126878 474628
rect 392 474488 4508 474516
rect -960 474460 4508 474488
rect 4564 474460 4574 474516
rect 263890 474460 263900 474516
rect 263956 474460 268072 474516
rect 331912 474460 335580 474516
rect 335636 474460 335646 474516
rect -960 474264 480 474460
rect 455868 474180 455924 474600
rect 456092 474516 456148 474796
rect 579628 474628 579684 475272
rect 535154 474572 535164 474628
rect 535220 474572 538104 474628
rect 579618 474572 579628 474628
rect 579684 474572 579694 474628
rect 456082 474460 456092 474516
rect 456148 474460 456158 474516
rect 455868 474124 457268 474180
rect 457212 474068 457268 474124
rect 457202 474012 457212 474068
rect 457268 474012 457278 474068
rect 82114 473900 82124 473956
rect 82180 473900 82190 473956
rect 123928 473900 127036 473956
rect 127092 473900 127102 473956
rect 185864 473900 189532 473956
rect 189588 473900 189598 473956
rect 247912 473900 262108 473956
rect 262164 473900 262174 473956
rect 264786 473900 264796 473956
rect 264852 473900 268072 473956
rect 331912 473900 335804 473956
rect 335860 473900 335870 473956
rect 348562 473900 348572 473956
rect 348628 473900 352072 473956
rect 402322 473900 402332 473956
rect 402388 473900 414120 473956
rect 455896 473900 457100 473956
rect 457156 473900 457166 473956
rect 517944 473900 521052 473956
rect 521108 473900 521118 473956
rect 345202 473788 345212 473844
rect 345268 473788 348684 473844
rect 348740 473788 348750 473844
rect 263778 473340 263788 473396
rect 263844 473340 268072 473396
rect 331912 473340 334460 473396
rect 334516 473340 334526 473396
rect 61880 473228 69804 473284
rect 69860 473228 69870 473284
rect 185864 473228 199052 473284
rect 199108 473228 199118 473284
rect 247912 473228 257852 473284
rect 257908 473228 257918 473284
rect 393960 473228 396844 473284
rect 396900 473228 396910 473284
rect 410722 473228 410732 473284
rect 410788 473228 414120 473284
rect 248098 472780 248108 472836
rect 248164 472780 268072 472836
rect 331912 472780 335132 472836
rect 335188 472780 335198 472836
rect 61880 472556 73052 472612
rect 73108 472556 73118 472612
rect 263778 472220 263788 472276
rect 263844 472220 268072 472276
rect 331912 472220 334460 472276
rect 334516 472220 334526 472276
rect 144396 471268 144452 471912
rect 393960 471884 395052 471940
rect 395108 471884 395118 471940
rect 247986 471660 247996 471716
rect 248052 471660 268072 471716
rect 331912 471660 351036 471716
rect 351092 471660 351102 471716
rect 61880 471212 64988 471268
rect 65044 471212 65054 471268
rect 144386 471212 144396 471268
rect 144452 471212 144462 471268
rect 256162 471100 256172 471156
rect 256228 471100 268072 471156
rect 331912 471100 334348 471156
rect 334404 471100 334414 471156
rect 247762 470540 247772 470596
rect 247828 470540 268072 470596
rect 331912 470540 334460 470596
rect 334516 470540 334526 470596
rect 262098 469980 262108 470036
rect 262164 469980 268072 470036
rect 331912 469980 338492 470036
rect 338548 469980 338558 470036
rect 579282 469868 579292 469924
rect 579348 469868 579358 469924
rect 585442 469868 585452 469924
rect 585508 469896 595672 469924
rect 585508 469868 597000 469896
rect 595560 469672 597000 469868
rect 334450 469532 334460 469588
rect 334516 469532 342076 469588
rect 342132 469532 342142 469588
rect 259858 469420 259868 469476
rect 259924 469420 268072 469476
rect 331912 469420 340284 469476
rect 340340 469420 340350 469476
rect 259522 468860 259532 468916
rect 259588 468860 268072 468916
rect 331912 468860 334460 468916
rect 334516 468860 334526 468916
rect 257842 468636 257852 468692
rect 257908 468636 263788 468692
rect 263844 468636 263854 468692
rect 258290 468300 258300 468356
rect 258356 468300 268072 468356
rect 331912 468300 340396 468356
rect 340452 468300 340462 468356
rect 189074 467852 189084 467908
rect 189140 467852 204092 467908
rect 204148 467852 204158 467908
rect 261314 467740 261324 467796
rect 261380 467740 268072 467796
rect 331912 467740 348572 467796
rect 348628 467740 348638 467796
rect 249554 467180 249564 467236
rect 249620 467180 268072 467236
rect 331912 467180 341964 467236
rect 342020 467180 342030 467236
rect 253138 466620 253148 466676
rect 253204 466620 268072 466676
rect 331912 466620 352156 466676
rect 352212 466620 352222 466676
rect 249442 466172 249452 466228
rect 249508 466172 263900 466228
rect 263956 466172 263966 466228
rect 259522 466060 259532 466116
rect 259588 466060 268072 466116
rect 331912 466060 342636 466116
rect 342692 466060 342702 466116
rect 252018 465500 252028 465556
rect 252084 465500 268072 465556
rect 331912 465500 345436 465556
rect 345492 465500 345502 465556
rect 61880 465164 81452 465220
rect 81508 465164 81518 465220
rect 263778 464940 263788 464996
rect 263844 464940 268072 464996
rect 331912 464940 345436 464996
rect 345492 464940 345502 464996
rect 249442 464380 249452 464436
rect 249508 464380 268072 464436
rect 331912 464380 334460 464436
rect 334516 464380 334526 464436
rect 264674 463820 264684 463876
rect 264740 463820 268072 463876
rect 331912 463820 350252 463876
rect 350308 463820 350318 463876
rect 263890 463260 263900 463316
rect 263956 463260 268072 463316
rect 331912 463260 352492 463316
rect 352548 463260 352558 463316
rect 398962 462812 398972 462868
rect 399028 462812 410844 462868
rect 410900 462812 410910 462868
rect 263778 462700 263788 462756
rect 263844 462700 268072 462756
rect 331912 462700 351036 462756
rect 351092 462700 351102 462756
rect 249554 462140 249564 462196
rect 249620 462140 268072 462196
rect 331912 462140 351932 462196
rect 351988 462140 351998 462196
rect 264002 461580 264012 461636
rect 264068 461580 268072 461636
rect 331912 461580 352604 461636
rect 352660 461580 352670 461636
rect 82002 461132 82012 461188
rect 82068 461132 82078 461188
rect 123928 461132 142156 461188
rect 142212 461132 142222 461188
rect 188962 461132 188972 461188
rect 189028 461132 205772 461188
rect 205828 461132 205838 461188
rect 256274 461020 256284 461076
rect 256340 461020 268072 461076
rect 331912 461020 334460 461076
rect 334516 461020 334526 461076
rect 264114 460460 264124 460516
rect 264180 460460 268072 460516
rect 331912 460460 334348 460516
rect 334404 460460 334414 460516
rect -960 460152 480 460376
rect 268044 459508 268100 459928
rect 331912 459900 335356 459956
rect 335412 459900 335422 459956
rect 255332 459452 268100 459508
rect 255332 459172 255388 459452
rect 263218 459340 263228 459396
rect 263284 459340 268072 459396
rect 331912 459340 518252 459396
rect 518308 459340 518318 459396
rect 143714 459116 143724 459172
rect 143780 459116 255388 459172
rect 204194 458780 204204 458836
rect 204260 458780 268072 458836
rect 331912 458780 518476 458836
rect 518532 458780 518542 458836
rect 261538 458220 261548 458276
rect 261604 458220 268072 458276
rect 331912 458220 474684 458276
rect 474740 458220 474750 458276
rect 230850 458108 230860 458164
rect 230916 458108 256172 458164
rect 256228 458108 256238 458164
rect 354386 458108 354396 458164
rect 354452 458108 459116 458164
rect 459172 458108 459182 458164
rect 160850 457996 160860 458052
rect 160916 457996 252028 458052
rect 252084 457996 252094 458052
rect 336018 457996 336028 458052
rect 336084 457996 459004 458052
rect 459060 457996 459070 458052
rect 142034 457884 142044 457940
rect 142100 457884 263900 457940
rect 263956 457884 263966 457940
rect 351026 457884 351036 457940
rect 351092 457884 493724 457940
rect 493780 457884 493790 457940
rect 495068 457884 502348 457940
rect 495068 457828 495124 457884
rect 69682 457772 69692 457828
rect 69748 457772 264684 457828
rect 264740 457772 264750 457828
rect 342626 457772 342636 457828
rect 342692 457772 495124 457828
rect 502292 457828 502348 457884
rect 502292 457772 558964 457828
rect 130162 457660 130172 457716
rect 130228 457660 268072 457716
rect 331912 457660 412412 457716
rect 412468 457660 412478 457716
rect 268044 457044 268100 457128
rect 133522 456988 133532 457044
rect 133588 456988 268100 457044
rect 331884 457044 331940 457128
rect 392466 457100 392476 457156
rect 392532 457100 396732 457156
rect 396788 457100 396798 457156
rect 493714 457100 493724 457156
rect 493780 457100 496860 457156
rect 496916 457100 496926 457156
rect 558908 457044 558964 457772
rect 331884 456988 457324 457044
rect 457380 456988 457390 457044
rect 558898 456988 558908 457044
rect 558964 456988 558974 457044
rect 160822 456876 160860 456932
rect 160916 456876 160926 456932
rect 230822 456876 230860 456932
rect 230916 456876 230926 456932
rect 229506 456652 229516 456708
rect 229572 456652 248108 456708
rect 248164 456652 248174 456708
rect 331884 456652 354396 456708
rect 354452 456652 354462 456708
rect 125122 456540 125132 456596
rect 125188 456540 268072 456596
rect 331884 456568 331940 456652
rect 352594 456540 352604 456596
rect 352660 456540 494844 456596
rect 494900 456540 494910 456596
rect 227490 456428 227500 456484
rect 227556 456428 259532 456484
rect 259588 456428 259598 456484
rect 352482 456428 352492 456484
rect 352548 456428 496188 456484
rect 496244 456428 496254 456484
rect 595560 456456 597000 456680
rect 336130 456316 336140 456372
rect 336196 456316 411180 456372
rect 411236 456316 411246 456372
rect 354386 456204 354396 456260
rect 354452 456204 459228 456260
rect 459284 456204 459294 456260
rect 82002 456092 82012 456148
rect 82068 456092 263788 456148
rect 263844 456092 263854 456148
rect 337698 456092 337708 456148
rect 337764 456092 458892 456148
rect 458948 456092 458958 456148
rect 135202 455980 135212 456036
rect 135268 455980 268072 456036
rect 331912 455980 430780 456036
rect 430836 455980 430846 456036
rect 136882 455420 136892 455476
rect 136948 455420 268072 455476
rect 331912 455420 455532 455476
rect 455588 455420 455598 455476
rect 226146 455196 226156 455252
rect 226212 455196 249564 455252
rect 249620 455196 249630 455252
rect 351922 455196 351932 455252
rect 351988 455196 501564 455252
rect 501620 455196 501630 455252
rect 231522 455084 231532 455140
rect 231588 455084 247772 455140
rect 247828 455084 247838 455140
rect 350242 455084 350252 455140
rect 350308 455084 493500 455140
rect 493556 455084 493566 455140
rect 258066 454860 258076 454916
rect 258132 454860 268072 454916
rect 331912 454860 457212 454916
rect 457268 454860 457278 454916
rect 138562 454300 138572 454356
rect 138628 454300 268072 454356
rect 331912 454300 456092 454356
rect 456148 454300 456158 454356
rect 263890 453740 263900 453796
rect 263956 453740 268072 453796
rect 331912 453740 337708 453796
rect 337764 453740 337774 453796
rect 222786 453516 222796 453572
rect 222852 453516 257852 453572
rect 257908 453516 257918 453572
rect 335122 453516 335132 453572
rect 335188 453516 562268 453572
rect 562324 453516 562334 453572
rect 342066 453404 342076 453460
rect 342132 453404 562940 453460
rect 562996 453404 563006 453460
rect 338482 453292 338492 453348
rect 338548 453292 555548 453348
rect 555604 453292 555614 453348
rect 103506 453180 103516 453236
rect 103572 453180 268072 453236
rect 331912 453180 337036 453236
rect 337092 453180 337102 453236
rect 340274 453180 340284 453236
rect 340340 453180 556220 453236
rect 556276 453180 556286 453236
rect 345426 453068 345436 453124
rect 345492 453068 498876 453124
rect 498932 453068 498942 453124
rect 80322 452844 80332 452900
rect 80388 452844 258188 452900
rect 258244 452844 258254 452900
rect 40226 452732 40236 452788
rect 40292 452732 247772 452788
rect 247828 452732 247838 452788
rect 263778 452620 263788 452676
rect 263844 452620 268072 452676
rect 331912 452620 336140 452676
rect 336196 452620 336206 452676
rect 104178 452060 104188 452116
rect 104244 452060 268072 452116
rect 331912 452060 336028 452116
rect 336084 452060 336094 452116
rect 372082 451948 372092 452004
rect 372148 451948 373548 452004
rect 373604 451948 373614 452004
rect 369618 451612 369628 451668
rect 369684 451612 374220 451668
rect 374276 451612 374286 451668
rect 82114 451500 82124 451556
rect 82180 451500 268072 451556
rect 331912 451500 457772 451556
rect 457828 451500 457838 451556
rect 335122 451164 335132 451220
rect 335188 451164 393372 451220
rect 393428 451164 393438 451220
rect 394034 451164 394044 451220
rect 394100 451164 494172 451220
rect 494228 451164 494238 451220
rect 20066 451052 20076 451108
rect 20132 451052 264908 451108
rect 264964 451052 264974 451108
rect 375442 451052 375452 451108
rect 375508 451052 561596 451108
rect 561652 451052 561662 451108
rect 142146 450940 142156 450996
rect 142212 450940 268072 450996
rect 331912 450940 398972 450996
rect 399028 450940 399038 450996
rect 143602 450380 143612 450436
rect 143668 450380 268072 450436
rect 331912 450380 354396 450436
rect 354452 450380 354462 450436
rect 222114 450268 222124 450324
rect 222180 450268 225932 450324
rect 225988 450268 225998 450324
rect 197362 449820 197372 449876
rect 197428 449820 268072 449876
rect 331912 449820 345212 449876
rect 345268 449820 345278 449876
rect 351922 449708 351932 449764
rect 351988 449708 396620 449764
rect 396676 449708 396686 449764
rect 342178 449596 342188 449652
rect 342244 449596 396844 449652
rect 396900 449596 396910 449652
rect 162866 449484 162876 449540
rect 162932 449484 170492 449540
rect 170548 449484 170558 449540
rect 392354 449484 392364 449540
rect 392420 449484 535052 449540
rect 535108 449484 535118 449540
rect 17938 449372 17948 449428
rect 18004 449372 247772 449428
rect 247828 449372 247838 449428
rect 352146 449372 352156 449428
rect 352212 449372 520940 449428
rect 520996 449372 521006 449428
rect 64754 449260 64764 449316
rect 64820 449260 268072 449316
rect 331912 449260 395052 449316
rect 395108 449260 395118 449316
rect 65090 448700 65100 448756
rect 65156 448700 268072 448756
rect 331912 448700 341852 448756
rect 341908 448700 341918 448756
rect 18162 448140 18172 448196
rect 18228 448140 268072 448196
rect 331912 448140 352044 448196
rect 352100 448140 352110 448196
rect 412402 447916 412412 447972
rect 412468 447916 499548 447972
rect 499604 447916 499614 447972
rect 195682 447804 195692 447860
rect 195748 447804 264572 447860
rect 264628 447804 264638 447860
rect 336802 447804 336812 447860
rect 336868 447804 458780 447860
rect 458836 447804 458846 447860
rect 102834 447692 102844 447748
rect 102900 447692 249564 447748
rect 249620 447692 249630 447748
rect 355282 447692 355292 447748
rect 355348 447692 535164 447748
rect 535220 447692 535230 447748
rect 64866 447580 64876 447636
rect 64932 447580 268072 447636
rect 331912 447580 392476 447636
rect 392532 447580 392542 447636
rect 199042 447020 199052 447076
rect 199108 447020 268072 447076
rect 331912 447020 395612 447076
rect 395668 447020 395678 447076
rect 344418 446572 344428 446628
rect 344484 446572 396508 446628
rect 396564 446572 396574 446628
rect 73154 446460 73164 446516
rect 73220 446460 268072 446516
rect 331912 446460 350476 446516
rect 350532 446460 350542 446516
rect 353602 446348 353612 446404
rect 353668 446348 410732 446404
rect 410788 446348 410798 446404
rect -960 446068 480 446264
rect 342290 446236 342300 446292
rect 342356 446236 410956 446292
rect 411012 446236 411022 446292
rect 370402 446124 370412 446180
rect 370468 446124 521164 446180
rect 521220 446124 521230 446180
rect -960 446040 78092 446068
rect 392 446012 78092 446040
rect 78148 446012 78158 446068
rect 127026 446012 127036 446068
rect 127092 446012 261324 446068
rect 261380 446012 261390 446068
rect 335794 446012 335804 446068
rect 335860 446012 348796 446068
rect 348852 446012 348862 446068
rect 350242 446012 350252 446068
rect 350308 446012 370188 446068
rect 370244 446012 370254 446068
rect 391346 446012 391356 446068
rect 391412 446012 583324 446068
rect 583380 446012 583390 446068
rect 78306 445900 78316 445956
rect 78372 445900 268072 445956
rect 331912 445900 369628 445956
rect 369684 445900 369694 445956
rect 62962 445340 62972 445396
rect 63028 445340 268072 445396
rect 331912 445340 345324 445396
rect 345380 445340 345390 445396
rect 345426 444892 345436 444948
rect 345492 444892 377580 444948
rect 377636 444892 377646 444948
rect 18050 444780 18060 444836
rect 18116 444780 268072 444836
rect 331912 444780 344428 444836
rect 344484 444780 344494 444836
rect 335906 444668 335916 444724
rect 335972 444668 394940 444724
rect 394996 444668 395006 444724
rect 338482 444556 338492 444612
rect 338548 444556 472892 444612
rect 472948 444556 472958 444612
rect 140802 444444 140812 444500
rect 140868 444444 253148 444500
rect 253204 444444 253214 444500
rect 371298 444444 371308 444500
rect 371364 444444 559580 444500
rect 559636 444444 559646 444500
rect 100818 444332 100828 444388
rect 100884 444332 258076 444388
rect 258132 444332 258142 444388
rect 335794 444332 335804 444388
rect 335860 444332 536732 444388
rect 536788 444332 536798 444388
rect 81442 444220 81452 444276
rect 81508 444220 268072 444276
rect 331912 444220 342076 444276
rect 342132 444220 342142 444276
rect 205762 443660 205772 443716
rect 205828 443660 268072 443716
rect 331912 443660 338828 443716
rect 338884 443660 338894 443716
rect 595560 443268 597000 443464
rect 333666 443212 333676 443268
rect 333732 443240 597000 443268
rect 333732 443212 595672 443240
rect 264898 443100 264908 443156
rect 264964 443100 268072 443156
rect 331912 443100 335916 443156
rect 335972 443100 335982 443156
rect 166226 442652 166236 442708
rect 166292 442652 202412 442708
rect 202468 442652 202478 442708
rect 264674 442540 264684 442596
rect 264740 442540 268072 442596
rect 331912 442540 335804 442596
rect 335860 442540 335870 442596
rect 203186 441980 203196 442036
rect 203252 441980 268072 442036
rect 331912 441980 371308 442036
rect 371364 441980 371374 442036
rect 261202 441868 261212 441924
rect 261268 441868 264292 441924
rect 264236 441812 264292 441868
rect 264236 441756 268100 441812
rect 268044 441448 268100 441756
rect 331912 441420 581308 441476
rect 581364 441420 581374 441476
rect 135202 441196 135212 441252
rect 135268 441196 265132 441252
rect 265188 441196 265198 441252
rect 64978 441084 64988 441140
rect 65044 441084 256172 441140
rect 256228 441084 256238 441140
rect 64642 440972 64652 441028
rect 64708 440972 259532 441028
rect 259588 440972 259598 441028
rect 256498 440860 256508 440916
rect 256564 440860 268072 440916
rect 331912 440860 530012 440916
rect 530068 440860 530078 440916
rect 252914 440300 252924 440356
rect 252980 440300 268072 440356
rect 331912 440300 391356 440356
rect 391412 440300 391422 440356
rect 252802 439740 252812 439796
rect 252868 439740 268072 439796
rect 331912 439740 392364 439796
rect 392420 439740 392430 439796
rect 130162 439628 130172 439684
rect 130228 439628 265356 439684
rect 265412 439628 265422 439684
rect 69794 439516 69804 439572
rect 69860 439516 264684 439572
rect 264740 439516 264750 439572
rect 44930 439404 44940 439460
rect 44996 439404 258300 439460
rect 258356 439404 258366 439460
rect 38210 439292 38220 439348
rect 38276 439292 253036 439348
rect 253092 439292 253102 439348
rect 334450 439292 334460 439348
rect 334516 439292 476252 439348
rect 476308 439292 476318 439348
rect 257842 439180 257852 439236
rect 257908 439180 268072 439236
rect 331912 439180 581420 439236
rect 581476 439180 581486 439236
rect 225922 438620 225932 438676
rect 225988 438620 268072 438676
rect 331912 438620 407484 438676
rect 407540 438620 407550 438676
rect 259634 438060 259644 438116
rect 259700 438060 268072 438116
rect 331912 438060 523292 438116
rect 523348 438060 523358 438116
rect 126802 437948 126812 438004
rect 126868 437948 247884 438004
rect 247940 437948 247950 438004
rect 74722 437836 74732 437892
rect 74788 437836 265020 437892
rect 265076 437836 265086 437892
rect 42914 437724 42924 437780
rect 42980 437724 261660 437780
rect 261716 437724 261726 437780
rect 335122 437724 335132 437780
rect 335188 437724 369516 437780
rect 369572 437724 369582 437780
rect 18274 437612 18284 437668
rect 18340 437612 261212 437668
rect 261268 437612 261278 437668
rect 335346 437612 335356 437668
rect 335412 437612 394828 437668
rect 394884 437612 394894 437668
rect 262882 437500 262892 437556
rect 262948 437500 268072 437556
rect 331912 437500 533372 437556
rect 533428 437500 533438 437556
rect 261426 436940 261436 436996
rect 261492 436940 268072 436996
rect 331912 436940 335804 436996
rect 335860 436940 335870 436996
rect 264562 436380 264572 436436
rect 264628 436380 268072 436436
rect 331912 436380 375452 436436
rect 375508 436380 375518 436436
rect 261314 435820 261324 435876
rect 261380 435820 268072 435876
rect 331912 435820 355292 435876
rect 355348 435820 355358 435876
rect 168914 435260 168924 435316
rect 168980 435260 268072 435316
rect 331912 435260 334460 435316
rect 334516 435260 334526 435316
rect 205762 434700 205772 434756
rect 205828 434700 268072 434756
rect 331912 434700 412412 434756
rect 412468 434700 412478 434756
rect 80546 434364 80556 434420
rect 80612 434364 263340 434420
rect 263396 434364 263406 434420
rect 73042 434252 73052 434308
rect 73108 434252 264572 434308
rect 264628 434252 264638 434308
rect 335234 434252 335244 434308
rect 335300 434252 372092 434308
rect 372148 434252 372158 434308
rect 166898 434140 166908 434196
rect 166964 434140 268072 434196
rect 331912 434140 394044 434196
rect 394100 434140 394110 434196
rect 204082 433580 204092 433636
rect 204148 433580 268072 433636
rect 331912 433580 519260 433636
rect 519316 433580 519326 433636
rect 141922 433020 141932 433076
rect 141988 433020 268072 433076
rect 331912 433020 519148 433076
rect 519204 433020 519214 433076
rect 335458 432684 335468 432740
rect 335524 432684 345212 432740
rect 345268 432684 345278 432740
rect 80434 432572 80444 432628
rect 80500 432572 255612 432628
rect 255668 432572 255678 432628
rect 335794 432572 335804 432628
rect 335860 432572 455420 432628
rect 455476 432572 455486 432628
rect 170482 432460 170492 432516
rect 170548 432460 268072 432516
rect 331912 432460 517468 432516
rect 517524 432460 517534 432516
rect -960 431956 480 432152
rect 202402 432012 202412 432068
rect 202468 432012 268100 432068
rect -960 431928 266364 431956
rect 392 431900 266364 431928
rect 266420 431900 266430 431956
rect 268044 431928 268100 432012
rect 331912 431900 467852 431956
rect 467908 431900 467918 431956
rect 187506 431340 187516 431396
rect 187572 431340 268072 431396
rect 331912 431340 464492 431396
rect 464548 431340 464558 431396
rect 192322 430780 192332 430836
rect 192388 430780 268072 430836
rect 331912 430780 461132 430836
rect 461188 430780 461198 430836
rect 38882 430668 38892 430724
rect 38948 430668 171388 430724
rect 171444 430668 171454 430724
rect 162866 430556 162876 430612
rect 162932 430556 187292 430612
rect 187348 430556 187358 430612
rect 230850 430556 230860 430612
rect 230916 430556 257852 430612
rect 257908 430556 257918 430612
rect 331884 430556 352156 430612
rect 352212 430556 352222 430612
rect 105522 430444 105532 430500
rect 105588 430444 130172 430500
rect 130228 430444 130238 430500
rect 168914 430444 168924 430500
rect 168980 430444 197372 430500
rect 197428 430444 197438 430500
rect 222114 430444 222124 430500
rect 222180 430444 249788 430500
rect 249844 430444 249854 430500
rect 103506 430332 103516 430388
rect 103572 430332 174636 430388
rect 174692 430332 174702 430388
rect 226818 430332 226828 430388
rect 226884 430332 259532 430388
rect 259588 430332 259598 430388
rect 39554 430220 39564 430276
rect 39620 430220 69692 430276
rect 69748 430220 69758 430276
rect 98130 430220 98140 430276
rect 98196 430220 223356 430276
rect 223412 430220 223422 430276
rect 228162 430220 228172 430276
rect 228228 430220 261212 430276
rect 261268 430220 261278 430276
rect 264562 430220 264572 430276
rect 264628 430220 268072 430276
rect 331884 430248 331940 430556
rect 351922 430444 351932 430500
rect 351988 430444 374892 430500
rect 374948 430444 374958 430500
rect 412402 430444 412412 430500
rect 412468 430444 436156 430500
rect 436212 430444 436222 430500
rect 467842 430444 467852 430500
rect 467908 430444 561596 430500
rect 561652 430444 561662 430500
rect 336914 430332 336924 430388
rect 336980 430332 494172 430388
rect 494228 430332 494238 430388
rect 338706 430220 338716 430276
rect 338772 430220 503580 430276
rect 503636 430220 503646 430276
rect 595560 430164 597000 430248
rect 161522 430108 161532 430164
rect 161588 430108 195692 430164
rect 195748 430108 195758 430164
rect 224130 430108 224140 430164
rect 224196 430108 263004 430164
rect 263060 430108 263070 430164
rect 345202 430108 345212 430164
rect 345268 430108 376908 430164
rect 376964 430108 376974 430164
rect 400642 430108 400652 430164
rect 400708 430108 597000 430164
rect 595560 430024 597000 430108
rect 187394 429660 187404 429716
rect 187460 429660 268072 429716
rect 331912 429660 370412 429716
rect 370468 429660 370478 429716
rect 223346 429212 223356 429268
rect 223412 429212 264684 429268
rect 264740 429212 264750 429268
rect 253138 429100 253148 429156
rect 253204 429100 268072 429156
rect 331912 429100 338492 429156
rect 338548 429100 338558 429156
rect 165554 428764 165564 428820
rect 165620 428764 192332 428820
rect 192388 428764 192398 428820
rect 240258 428764 240268 428820
rect 240324 428764 259756 428820
rect 259812 428764 259822 428820
rect 164210 428652 164220 428708
rect 164276 428652 252924 428708
rect 252980 428652 252990 428708
rect 345314 428652 345324 428708
rect 345380 428652 435484 428708
rect 435540 428652 435550 428708
rect 102834 428540 102844 428596
rect 102900 428540 249452 428596
rect 249508 428540 249518 428596
rect 255602 428540 255612 428596
rect 255668 428540 268072 428596
rect 331912 428540 404012 428596
rect 404068 428540 404078 428596
rect 462802 428540 462812 428596
rect 462868 428540 560252 428596
rect 560308 428540 560318 428596
rect 42914 428428 42924 428484
rect 42980 428428 256172 428484
rect 256228 428428 256238 428484
rect 340274 428428 340284 428484
rect 340340 428428 500892 428484
rect 500948 428428 500958 428484
rect 265346 427980 265356 428036
rect 265412 427980 268072 428036
rect 331912 427980 402332 428036
rect 402388 427980 402398 428036
rect 171378 427644 171388 427700
rect 171444 427644 264572 427700
rect 264628 427644 264638 427700
rect 38546 427532 38556 427588
rect 38612 427532 264796 427588
rect 264852 427532 264862 427588
rect 334450 427532 334460 427588
rect 334516 427532 455308 427588
rect 455364 427532 455374 427588
rect 259634 427420 259644 427476
rect 259700 427420 268072 427476
rect 331912 427420 457100 427476
rect 457156 427420 457166 427476
rect 229618 427196 229628 427252
rect 229684 427196 247884 427252
rect 247940 427196 247950 427252
rect 167570 427084 167580 427140
rect 167636 427084 188972 427140
rect 189028 427084 189038 427140
rect 211362 427084 211372 427140
rect 211428 427084 256284 427140
rect 256340 427084 256350 427140
rect 99474 426972 99484 427028
rect 99540 426972 252812 427028
rect 252868 426972 252878 427028
rect 436790 426972 436828 427028
rect 436884 426972 436894 427028
rect 438134 426972 438172 427028
rect 438228 426972 438238 427028
rect 474674 426972 474684 427028
rect 474740 426972 556220 427028
rect 556276 426972 556286 427028
rect 102162 426860 102172 426916
rect 102228 426860 258188 426916
rect 258244 426860 258254 426916
rect 265122 426860 265132 426916
rect 265188 426860 268072 426916
rect 331912 426860 335804 426916
rect 335860 426860 335870 426916
rect 338482 426860 338492 426916
rect 338548 426860 493500 426916
rect 493556 426860 493566 426916
rect 40226 426748 40236 426804
rect 40292 426748 261324 426804
rect 261380 426748 261390 426804
rect 342066 426748 342076 426804
rect 342132 426748 500220 426804
rect 500276 426748 500286 426804
rect 166226 426636 166236 426692
rect 166292 426636 173852 426692
rect 173908 426636 173918 426692
rect 174626 426636 174636 426692
rect 174692 426636 264908 426692
rect 264964 426636 264974 426692
rect 331884 426636 400652 426692
rect 400708 426636 400718 426692
rect 407362 426636 407372 426692
rect 407428 426636 497532 426692
rect 497588 426636 497598 426692
rect 44258 426524 44268 426580
rect 44324 426524 73052 426580
rect 73108 426524 73118 426580
rect 82226 426524 82236 426580
rect 82292 426524 268100 426580
rect 88050 426412 88060 426468
rect 88116 426412 90748 426468
rect 160850 426412 160860 426468
rect 160916 426412 167860 426468
rect 170230 426412 170268 426468
rect 170324 426412 170334 426468
rect 222758 426412 222796 426468
rect 222852 426412 222862 426468
rect 232166 426412 232204 426468
rect 232260 426412 232270 426468
rect 90692 426356 90748 426412
rect 90692 426300 156268 426356
rect 156212 426132 156268 426300
rect 167804 426244 167860 426412
rect 167972 426300 170212 426356
rect 173730 426300 173740 426356
rect 173796 426300 257964 426356
rect 258020 426300 258030 426356
rect 268044 426328 268100 426524
rect 331884 426328 331940 426636
rect 334450 426524 334460 426580
rect 334516 426524 398972 426580
rect 399028 426524 399038 426580
rect 399186 426524 399196 426580
rect 399252 426524 557564 426580
rect 557620 426524 557630 426580
rect 478772 426412 502908 426468
rect 502964 426412 502974 426468
rect 478772 426356 478828 426412
rect 352034 426300 352044 426356
rect 352100 426300 478828 426356
rect 167972 426244 168028 426300
rect 167804 426188 168028 426244
rect 170156 426244 170212 426300
rect 170156 426188 249676 426244
rect 249732 426188 249742 426244
rect 341842 426188 341852 426244
rect 341908 426188 436828 426244
rect 436884 426188 436894 426244
rect 438162 426188 438172 426244
rect 438228 426188 438238 426244
rect 438172 426132 438228 426188
rect 156212 426076 168028 426132
rect 170258 426076 170268 426132
rect 170324 426076 170334 426132
rect 173842 426076 173852 426132
rect 173908 426076 189084 426132
rect 189140 426076 189150 426132
rect 222786 426076 222796 426132
rect 222852 426076 263116 426132
rect 263172 426076 263182 426132
rect 404002 426076 404012 426132
rect 404068 426076 438228 426132
rect 167972 425908 168028 426076
rect 170268 426020 170324 426076
rect 170268 425964 187404 426020
rect 187460 425964 187470 426020
rect 232194 425964 232204 426020
rect 232260 425964 253148 426020
rect 253204 425964 253214 426020
rect 167972 425852 173740 425908
rect 173796 425852 173806 425908
rect 263330 425740 263340 425796
rect 263396 425740 268072 425796
rect 331912 425740 353612 425796
rect 353668 425740 353678 425796
rect 258178 425180 258188 425236
rect 258244 425180 268072 425236
rect 331912 425180 342300 425236
rect 342356 425180 342366 425236
rect 200722 424620 200732 424676
rect 200788 424620 268072 424676
rect 331912 424620 456988 424676
rect 457044 424620 457054 424676
rect 247874 424060 247884 424116
rect 247940 424060 268072 424116
rect 331912 424060 336812 424116
rect 336868 424060 336878 424116
rect 261314 423500 261324 423556
rect 261380 423500 268072 423556
rect 331912 423500 334460 423556
rect 334516 423500 334526 423556
rect 249554 422940 249564 422996
rect 249620 422940 268072 422996
rect 331912 422940 350364 422996
rect 350420 422940 350430 422996
rect 258066 422380 258076 422436
rect 258132 422380 268072 422436
rect 331912 422380 334460 422436
rect 334516 422380 334526 422436
rect 253026 421820 253036 421876
rect 253092 421820 268072 421876
rect 331912 421820 345436 421876
rect 345492 421820 345502 421876
rect 348786 421484 348796 421540
rect 348852 421484 352072 421540
rect 393960 421484 396620 421540
rect 396676 421484 396686 421540
rect 410722 421484 410732 421540
rect 410788 421484 414120 421540
rect 472098 421484 472108 421540
rect 472164 421484 476056 421540
rect 247762 421260 247772 421316
rect 247828 421260 268072 421316
rect 331912 421260 348572 421316
rect 348628 421260 348638 421316
rect 259522 420700 259532 420756
rect 259588 420700 268072 420756
rect 331912 420700 335132 420756
rect 335188 420700 335198 420756
rect 261202 420140 261212 420196
rect 261268 420140 268072 420196
rect 331912 420140 340172 420196
rect 340228 420140 340238 420196
rect 393932 420084 393988 420840
rect 393932 420028 395668 420084
rect 395612 419972 395668 420028
rect 395602 419916 395612 419972
rect 395668 419916 395678 419972
rect 247762 419580 247772 419636
rect 247828 419580 268072 419636
rect 331912 419580 342188 419636
rect 342244 419580 342254 419636
rect 256162 419020 256172 419076
rect 256228 419020 268072 419076
rect 331912 419020 335356 419076
rect 335412 419020 335422 419076
rect 264562 418460 264572 418516
rect 264628 418460 268072 418516
rect 331912 418460 338604 418516
rect 338660 418460 338670 418516
rect -960 417816 480 418040
rect 262882 417900 262892 417956
rect 262948 417900 268072 417956
rect 331912 417900 335244 417956
rect 335300 417900 335310 417956
rect 258290 417340 258300 417396
rect 258356 417340 268072 417396
rect 331912 417340 350252 417396
rect 350308 417340 350318 417396
rect 261650 416780 261660 416836
rect 261716 416780 268072 416836
rect 331912 416780 335468 416836
rect 335524 416780 335534 416836
rect 595560 416808 597000 417032
rect 264674 416220 264684 416276
rect 264740 416220 268072 416276
rect 331912 416220 351932 416276
rect 351988 416220 351998 416276
rect 265010 415660 265020 415716
rect 265076 415660 268072 415716
rect 331912 415660 335132 415716
rect 335188 415660 335198 415716
rect 206556 415044 206612 415464
rect 263890 415100 263900 415156
rect 263956 415100 268072 415156
rect 331912 415100 334460 415156
rect 334516 415100 334526 415156
rect 206556 414988 206668 415044
rect 206724 414988 206734 415044
rect 247874 414540 247884 414596
rect 247940 414540 268072 414596
rect 331912 414540 334460 414596
rect 334516 414540 334526 414596
rect 262882 413980 262892 414036
rect 262948 413980 268072 414036
rect 331912 413980 335132 414036
rect 335188 413980 335198 414036
rect 263330 413420 263340 413476
rect 263396 413420 268072 413476
rect 331912 413420 334460 413476
rect 334516 413420 334526 413476
rect 472098 413420 472108 413476
rect 472164 413420 476056 413476
rect 263778 412860 263788 412916
rect 263844 412860 268072 412916
rect 331912 412860 351036 412916
rect 351092 412860 351102 412916
rect 82674 412748 82684 412804
rect 82740 412748 82750 412804
rect 141026 412748 141036 412804
rect 141092 412748 144060 412804
rect 144116 412748 144126 412804
rect 253138 412300 253148 412356
rect 253204 412300 268072 412356
rect 331912 412300 334348 412356
rect 334404 412300 334414 412356
rect 18358 411740 18396 411796
rect 18452 411740 18462 411796
rect 20076 411684 20132 412104
rect 201618 412076 201628 412132
rect 201684 412076 206136 412132
rect 247912 412076 262108 412132
rect 262164 412076 262174 412132
rect 472098 412076 472108 412132
rect 472164 412076 476056 412132
rect 258066 411740 258076 411796
rect 258132 411740 268072 411796
rect 331912 411740 334460 411796
rect 334516 411740 334526 411796
rect 19954 411628 19964 411684
rect 20020 411628 20132 411684
rect 18050 411404 18060 411460
rect 18116 411404 20104 411460
rect 123928 411404 135212 411460
rect 135268 411404 135278 411460
rect 349346 411404 349356 411460
rect 349412 411404 352716 411460
rect 352772 411404 352782 411460
rect 411506 411404 411516 411460
rect 411572 411404 414652 411460
rect 414708 411404 414718 411460
rect 464482 411404 464492 411460
rect 464548 411404 476056 411460
rect 534370 411404 534380 411460
rect 534436 411404 538104 411460
rect 261426 411180 261436 411236
rect 261492 411180 268072 411236
rect 331912 411180 334460 411236
rect 334516 411180 334526 411236
rect 19842 410732 19852 410788
rect 19908 410732 20104 410788
rect 61880 410732 69692 410788
rect 69748 410732 69758 410788
rect 123928 410732 127036 410788
rect 127092 410732 127102 410788
rect 455896 410732 457324 410788
rect 457380 410732 457390 410788
rect 473106 410732 473116 410788
rect 473172 410732 476056 410788
rect 530002 410732 530012 410788
rect 530068 410732 538104 410788
rect 579282 410732 579292 410788
rect 579348 410732 579358 410788
rect 262098 410620 262108 410676
rect 262164 410620 268072 410676
rect 331912 410620 335356 410676
rect 335412 410620 335422 410676
rect 579618 410620 579628 410676
rect 579684 410620 579694 410676
rect 247884 410172 263900 410228
rect 263956 410172 263966 410228
rect 19730 410060 19740 410116
rect 19796 410060 20104 410116
rect 61880 410060 74732 410116
rect 74788 410060 74798 410116
rect 82674 410060 82684 410116
rect 82740 410060 82750 410116
rect 123928 410060 126812 410116
rect 126868 410060 126878 410116
rect 142706 410060 142716 410116
rect 142772 410060 144088 410116
rect 247884 410088 247940 410172
rect 259746 410060 259756 410116
rect 259812 410060 268072 410116
rect 331912 410060 334348 410116
rect 334404 410060 334414 410116
rect 338594 410060 338604 410116
rect 338660 410060 352072 410116
rect 393960 410060 394828 410116
rect 394884 410060 394894 410116
rect 402322 410060 402332 410116
rect 402388 410060 414120 410116
rect 144274 409836 144284 409892
rect 144340 409836 144350 409892
rect 18386 409388 18396 409444
rect 18452 409388 20104 409444
rect 61880 409388 79772 409444
rect 79828 409388 79838 409444
rect 123928 409388 126252 409444
rect 126308 409388 126318 409444
rect 144284 409416 144340 409836
rect 249778 409500 249788 409556
rect 249844 409500 268072 409556
rect 331912 409500 334460 409556
rect 334516 409500 334526 409556
rect 455868 409444 455924 410088
rect 517944 410060 521052 410116
rect 521108 410060 521118 410116
rect 534258 410060 534268 410116
rect 534324 410060 538104 410116
rect 579628 410088 579684 410620
rect 203186 409388 203196 409444
rect 203252 409388 206136 409444
rect 347778 409388 347788 409444
rect 347844 409388 352072 409444
rect 455868 409388 456092 409444
rect 456148 409388 456158 409444
rect 533362 409388 533372 409444
rect 533428 409388 538104 409444
rect 579282 409388 579292 409444
rect 579348 409388 579358 409444
rect 334338 409052 334348 409108
rect 334404 409052 350364 409108
rect 350420 409052 350430 409108
rect 260306 408940 260316 408996
rect 260372 408940 268072 408996
rect 331912 408940 348572 408996
rect 348628 408940 348638 408996
rect 123928 408716 127260 408772
rect 127316 408716 127326 408772
rect 144284 408436 144340 408744
rect 206098 408716 206108 408772
rect 206164 408716 206174 408772
rect 455896 408716 458892 408772
rect 458948 408716 458958 408772
rect 467842 408716 467852 408772
rect 467908 408716 476056 408772
rect 535826 408716 535836 408772
rect 535892 408716 538104 408772
rect 144274 408380 144284 408436
rect 144340 408380 144350 408436
rect 256274 408380 256284 408436
rect 256340 408380 268072 408436
rect 331912 408380 335580 408436
rect 335636 408380 335646 408436
rect 18274 408044 18284 408100
rect 18340 408044 20104 408100
rect 20636 406756 20692 407400
rect 61880 407372 76412 407428
rect 76468 407372 76478 407428
rect 82348 407316 82404 408072
rect 144396 407316 144452 408072
rect 185864 408044 188972 408100
rect 189028 408044 189038 408100
rect 204866 408044 204876 408100
rect 204932 408044 206136 408100
rect 247912 408044 263340 408100
rect 263396 408044 263406 408100
rect 338482 408044 338492 408100
rect 338548 408044 352072 408100
rect 393960 408044 394940 408100
rect 394996 408044 395006 408100
rect 455896 408044 458780 408100
rect 458836 408044 458846 408100
rect 517944 408044 519148 408100
rect 519204 408044 519214 408100
rect 535042 408044 535052 408100
rect 535108 408044 538104 408100
rect 263106 407820 263116 407876
rect 263172 407820 268072 407876
rect 331912 407820 334460 407876
rect 334516 407820 334526 407876
rect 185864 407372 199836 407428
rect 199892 407372 199902 407428
rect 247912 407372 256172 407428
rect 256228 407372 256238 407428
rect 411170 407372 411180 407428
rect 411236 407372 414120 407428
rect 455522 407372 455532 407428
rect 455588 407372 455598 407428
rect 579880 407372 581308 407428
rect 581364 407372 581374 407428
rect 82338 407260 82348 407316
rect 82404 407260 82414 407316
rect 144386 407260 144396 407316
rect 144452 407260 144462 407316
rect 263778 407260 263788 407316
rect 263844 407260 268072 407316
rect 331912 407260 336924 407316
rect 336980 407260 336990 407316
rect 20626 406700 20636 406756
rect 20692 406700 20702 406756
rect 61880 406700 81452 406756
rect 81508 406700 81518 406756
rect 123928 406700 136108 406756
rect 136164 406700 136174 406756
rect 144284 406644 144340 406728
rect 247912 406700 259532 406756
rect 259588 406700 259598 406756
rect 260306 406700 260316 406756
rect 260372 406700 268072 406756
rect 331912 406700 338716 406756
rect 338772 406700 338782 406756
rect 411058 406700 411068 406756
rect 411124 406700 414120 406756
rect 455896 406700 457100 406756
rect 457156 406700 457166 406756
rect 579618 406700 579628 406756
rect 579684 406700 579694 406756
rect 144274 406588 144284 406644
rect 144340 406588 144350 406644
rect 579842 406476 579852 406532
rect 579908 406476 579918 406532
rect 262098 406140 262108 406196
rect 262164 406140 268072 406196
rect 331912 406140 342076 406196
rect 342132 406140 342142 406196
rect 61880 406028 64652 406084
rect 64708 406028 64718 406084
rect 123928 406028 127148 406084
rect 127204 406028 127214 406084
rect 185864 406028 191548 406084
rect 191604 406028 191614 406084
rect 247912 406028 253148 406084
rect 253204 406028 253214 406084
rect 341842 406028 341852 406084
rect 341908 406028 352072 406084
rect 393960 406028 395052 406084
rect 395108 406028 395118 406084
rect 406578 406028 406588 406084
rect 406644 406028 414120 406084
rect 455896 406028 458668 406084
rect 458724 406028 458734 406084
rect 472882 406028 472892 406084
rect 472948 406028 476056 406084
rect 579852 406056 579908 406476
rect 252914 405580 252924 405636
rect 252980 405580 268072 405636
rect 331912 405580 336028 405636
rect 336084 405580 336094 405636
rect 517916 405412 517972 406056
rect 61880 405356 73052 405412
rect 73108 405356 73118 405412
rect 185864 405356 204988 405412
rect 205044 405356 205054 405412
rect 455896 405356 456988 405412
rect 457044 405356 457054 405412
rect 517916 405356 519988 405412
rect 579880 405356 583100 405412
rect 583156 405356 583166 405412
rect 519932 405300 519988 405356
rect 519922 405244 519932 405300
rect 519988 405244 519998 405300
rect 263890 405020 263900 405076
rect 263956 405020 268072 405076
rect 331912 405020 352044 405076
rect 352100 405020 352110 405076
rect 61880 404684 81564 404740
rect 81620 404684 81630 404740
rect 185864 404684 189420 404740
rect 189476 404684 189486 404740
rect 393960 404684 396508 404740
rect 396564 404684 396574 404740
rect 411170 404684 411180 404740
rect 411236 404684 414120 404740
rect 455896 404684 459004 404740
rect 459060 404684 459070 404740
rect 263778 404460 263788 404516
rect 263844 404460 268072 404516
rect 331912 404460 340284 404516
rect 340340 404460 340350 404516
rect 123928 404012 126924 404068
rect 126980 404012 126990 404068
rect 185864 404012 189532 404068
rect 189588 404012 189598 404068
rect 455896 404012 457212 404068
rect 457268 404012 457278 404068
rect 461122 404012 461132 404068
rect 461188 404012 473116 404068
rect 473172 404012 473182 404068
rect -960 403732 480 403928
rect 263442 403900 263452 403956
rect 263508 403900 268072 403956
rect 331912 403900 334460 403956
rect 334516 403900 334526 403956
rect -960 403704 7532 403732
rect 392 403676 7532 403704
rect 7588 403676 7598 403732
rect 595560 403620 597000 403816
rect 580626 403564 580636 403620
rect 580692 403592 597000 403620
rect 580692 403564 595672 403592
rect 252802 403452 252812 403508
rect 252868 403452 268100 403508
rect 141026 403340 141036 403396
rect 141092 403340 144088 403396
rect 185864 403340 189308 403396
rect 189364 403340 189374 403396
rect 247912 403340 262892 403396
rect 262948 403340 262958 403396
rect 268044 403368 268100 403452
rect 331912 403340 350252 403396
rect 350308 403340 350318 403396
rect 393960 403340 396732 403396
rect 396788 403340 396798 403396
rect 455298 403340 455308 403396
rect 455364 403340 455374 403396
rect 472098 403340 472108 403396
rect 472164 403340 476056 403396
rect 340498 403228 340508 403284
rect 340564 403228 347788 403284
rect 347844 403228 347854 403284
rect 579730 403116 579740 403172
rect 579796 403116 579806 403172
rect 263778 402780 263788 402836
rect 263844 402780 268072 402836
rect 331912 402780 334460 402836
rect 334516 402780 334526 402836
rect 20066 402668 20076 402724
rect 20132 402668 20142 402724
rect 123928 402668 143612 402724
rect 143668 402668 143678 402724
rect 247912 402668 259644 402724
rect 259700 402668 259710 402724
rect 345202 402668 345212 402724
rect 345268 402668 352072 402724
rect 401202 402668 401212 402724
rect 401268 402668 414120 402724
rect 455410 402668 455420 402724
rect 455476 402668 455486 402724
rect 517944 402668 520940 402724
rect 520996 402668 521006 402724
rect 579740 402696 579796 403116
rect 579618 402556 579628 402612
rect 579684 402556 579694 402612
rect 398962 402332 398972 402388
rect 399028 402332 411180 402388
rect 411236 402332 411246 402388
rect 249666 402220 249676 402276
rect 249732 402220 268072 402276
rect 331912 402220 337708 402276
rect 337652 402052 337708 402220
rect 185864 401996 189532 402052
rect 189588 401996 189598 402052
rect 204754 401996 204764 402052
rect 204820 401996 206136 402052
rect 337652 401996 352044 402052
rect 352100 401996 352110 402052
rect 411170 401996 411180 402052
rect 411236 401996 414120 402052
rect 461122 401996 461132 402052
rect 461188 401996 476056 402052
rect 517458 401996 517468 402052
rect 517524 401996 517534 402052
rect 534258 401996 534268 402052
rect 534324 401996 538104 402052
rect 579628 402024 579684 402556
rect 263890 401660 263900 401716
rect 263956 401660 268072 401716
rect 331912 401660 350252 401716
rect 350308 401660 350318 401716
rect 18162 401324 18172 401380
rect 18228 401324 20104 401380
rect 61880 401324 64876 401380
rect 64932 401324 64942 401380
rect 82348 400708 82404 401352
rect 123928 401324 133532 401380
rect 133588 401324 133598 401380
rect 185864 401324 192332 401380
rect 192388 401324 192398 401380
rect 517234 401324 517244 401380
rect 517300 401324 517310 401380
rect 247762 401100 247772 401156
rect 247828 401100 268072 401156
rect 331912 401100 334348 401156
rect 334404 401100 334414 401156
rect 82338 400652 82348 400708
rect 82404 400652 82414 400708
rect 535602 400652 535612 400708
rect 535668 400652 538104 400708
rect 262098 400540 262108 400596
rect 262164 400540 268072 400596
rect 331912 400540 345436 400596
rect 345492 400540 345502 400596
rect 262210 399980 262220 400036
rect 262276 399980 268072 400036
rect 331912 399980 338492 400036
rect 338548 399980 338558 400036
rect 258178 399420 258188 399476
rect 258244 399420 268072 399476
rect 331912 399420 336252 399476
rect 336308 399420 336318 399476
rect 336802 398972 336812 399028
rect 336868 398972 348796 399028
rect 348852 398972 348862 399028
rect 264674 398860 264684 398916
rect 264740 398860 268072 398916
rect 331912 398860 334460 398916
rect 334516 398860 334526 398916
rect 533474 398524 533484 398580
rect 533540 398524 535612 398580
rect 535668 398524 535678 398580
rect 263778 398300 263788 398356
rect 263844 398300 268072 398356
rect 331912 398300 351036 398356
rect 351092 398300 351102 398356
rect 263778 397740 263788 397796
rect 263844 397740 268072 397796
rect 331912 397740 350364 397796
rect 350420 397740 350430 397796
rect 264898 397180 264908 397236
rect 264964 397180 268072 397236
rect 331912 397180 334460 397236
rect 334516 397180 334526 397236
rect 249442 396620 249452 396676
rect 249508 396620 268072 396676
rect 331912 396620 334348 396676
rect 334404 396620 334414 396676
rect 252802 396060 252812 396116
rect 252868 396060 268072 396116
rect 331912 396060 334460 396116
rect 334516 396060 334526 396116
rect 188962 395612 188972 395668
rect 189028 395612 205772 395668
rect 205828 395612 205838 395668
rect 263778 395500 263788 395556
rect 263844 395500 268072 395556
rect 331912 395500 334348 395556
rect 334404 395500 334414 395556
rect 61880 395276 74844 395332
rect 74900 395276 74910 395332
rect 263890 394940 263900 394996
rect 263956 394940 268072 394996
rect 331912 394940 345324 394996
rect 345380 394940 345390 394996
rect 249442 394380 249452 394436
rect 249508 394380 268072 394436
rect 331912 394380 334460 394436
rect 334516 394380 334526 394436
rect 249666 393820 249676 393876
rect 249732 393820 268072 393876
rect 331912 393820 334348 393876
rect 334404 393820 334414 393876
rect 256274 393260 256284 393316
rect 256340 393260 268072 393316
rect 331912 393260 341852 393316
rect 341908 393260 341918 393316
rect 263778 392700 263788 392756
rect 263844 392700 268072 392756
rect 331912 392700 334348 392756
rect 334404 392700 334414 392756
rect 257954 392140 257964 392196
rect 258020 392140 268072 392196
rect 331912 392140 334460 392196
rect 334516 392140 334526 392196
rect 256162 391580 256172 391636
rect 256228 391580 268072 391636
rect 331912 391580 352492 391636
rect 352548 391580 352558 391636
rect 263778 391020 263788 391076
rect 263844 391020 268072 391076
rect 331912 391020 347788 391076
rect 347844 391020 347854 391076
rect 579618 391020 579628 391076
rect 579684 391020 579694 391076
rect 579628 390600 579684 391020
rect 590594 390572 590604 390628
rect 590660 390600 595672 390628
rect 590660 390572 597000 390600
rect 263890 390460 263900 390516
rect 263956 390460 268072 390516
rect 331912 390460 350588 390516
rect 350644 390460 350654 390516
rect 455522 390460 455532 390516
rect 455588 390460 455598 390516
rect 263778 389900 263788 389956
rect 263844 389900 268072 389956
rect 331912 389900 341852 389956
rect 341908 389900 341918 389956
rect 455532 389928 455588 390460
rect 595560 390376 597000 390572
rect -960 389620 480 389816
rect -960 389592 15932 389620
rect 392 389564 15932 389592
rect 15988 389564 15998 389620
rect 264562 389340 264572 389396
rect 264628 389340 268072 389396
rect 331912 389340 352604 389396
rect 352660 389340 352670 389396
rect 253138 388892 253148 388948
rect 253204 388892 265020 388948
rect 265076 388892 265086 388948
rect 261314 388780 261324 388836
rect 261380 388780 268072 388836
rect 331912 388780 336028 388836
rect 336084 388780 336094 388836
rect 264786 388220 264796 388276
rect 264852 388220 268072 388276
rect 331912 388220 340508 388276
rect 340564 388220 340574 388276
rect 20066 387996 20076 388052
rect 20132 387996 263900 388052
rect 263956 387996 263966 388052
rect 81554 387884 81564 387940
rect 81620 387884 263788 387940
rect 263844 387884 263854 387940
rect 74722 387660 74732 387716
rect 74788 387660 268072 387716
rect 331912 387660 338604 387716
rect 338660 387660 338670 387716
rect 349458 387660 349468 387716
rect 349524 387660 396620 387716
rect 396676 387660 396686 387716
rect 335122 387548 335132 387604
rect 335188 387548 535948 387604
rect 536004 387548 536014 387604
rect 335570 387436 335580 387492
rect 335636 387436 537740 387492
rect 537796 387436 537806 387492
rect 335346 387324 335356 387380
rect 335412 387324 537628 387380
rect 537684 387324 537694 387380
rect 347778 387212 347788 387268
rect 347844 387212 583100 387268
rect 583156 387212 583166 387268
rect 73042 387100 73052 387156
rect 73108 387100 268072 387156
rect 331912 387100 351148 387156
rect 351204 387100 351214 387156
rect 19842 386540 19852 386596
rect 19908 386540 268072 386596
rect 331912 386540 336812 386596
rect 336868 386540 336878 386596
rect 259522 386316 259532 386372
rect 259588 386316 263788 386372
rect 263844 386316 263854 386372
rect 268044 385924 268100 386008
rect 69682 385868 69692 385924
rect 69748 385868 268100 385924
rect 331884 385924 331940 386008
rect 331884 385868 370860 385924
rect 370916 385868 370926 385924
rect 347778 385756 347788 385812
rect 347844 385756 374220 385812
rect 374276 385756 374286 385812
rect 503122 385756 503132 385812
rect 503188 385756 520940 385812
rect 520996 385756 521006 385812
rect 336018 385644 336028 385700
rect 336084 385644 370188 385700
rect 370244 385644 370254 385700
rect 371298 385644 371308 385700
rect 371364 385644 535052 385700
rect 535108 385644 535118 385700
rect 230850 385532 230860 385588
rect 230916 385532 261436 385588
rect 261492 385532 261502 385588
rect 331884 385532 395612 385588
rect 395668 385532 395678 385588
rect 400642 385532 400652 385588
rect 400708 385532 472892 385588
rect 472948 385532 472958 385588
rect 476242 385532 476252 385588
rect 476308 385532 521052 385588
rect 521108 385532 521118 385588
rect 81442 385420 81452 385476
rect 81508 385420 268072 385476
rect 331884 385448 331940 385532
rect 350242 385420 350252 385476
rect 350308 385420 495516 385476
rect 495572 385420 495582 385476
rect 168242 385308 168252 385364
rect 168308 385308 247772 385364
rect 247828 385308 247838 385364
rect 345426 385308 345436 385364
rect 345492 385308 367052 385364
rect 367108 385308 367118 385364
rect 372866 385308 372876 385364
rect 372932 385308 372942 385364
rect 384692 385308 499548 385364
rect 499604 385308 499614 385364
rect 372876 385252 372932 385308
rect 352482 385196 352492 385252
rect 352548 385196 372932 385252
rect 352594 385084 352604 385140
rect 352660 385084 369068 385140
rect 369124 385084 369134 385140
rect 384692 385028 384748 385308
rect 367042 384972 367052 385028
rect 367108 384972 384748 385028
rect 19954 384860 19964 384916
rect 20020 384860 268072 384916
rect 331912 384860 335916 384916
rect 335972 384860 335982 384916
rect 105522 384636 105532 384692
rect 105588 384636 256284 384692
rect 256340 384636 256350 384692
rect 370850 384636 370860 384692
rect 370916 384636 376908 384692
rect 376964 384636 376974 384692
rect 106194 384524 106204 384580
rect 106260 384524 249676 384580
rect 249732 384524 249742 384580
rect 331884 384524 349468 384580
rect 349524 384524 349534 384580
rect 352034 384524 352044 384580
rect 352100 384524 498876 384580
rect 498932 384524 498942 384580
rect 222786 384412 222796 384468
rect 222852 384412 258076 384468
rect 258132 384412 258142 384468
rect 74834 384300 74844 384356
rect 74900 384300 268072 384356
rect 331884 384328 331940 384524
rect 350354 384412 350364 384468
rect 350420 384412 430780 384468
rect 430836 384412 430846 384468
rect 350578 384300 350588 384356
rect 350644 384300 375564 384356
rect 375620 384300 375630 384356
rect 341842 384188 341852 384244
rect 341908 384188 368844 384244
rect 368900 384188 368910 384244
rect 351138 384076 351148 384132
rect 351204 384076 374892 384132
rect 374948 384076 374958 384132
rect 348562 383964 348572 384020
rect 348628 383964 559580 384020
rect 559636 383964 559646 384020
rect 335906 383852 335916 383908
rect 335972 383852 352716 383908
rect 352772 383852 352782 383908
rect 203186 383740 203196 383796
rect 203252 383740 268072 383796
rect 331912 383740 581308 383796
rect 581364 383740 581374 383796
rect 259634 383180 259644 383236
rect 259700 383180 268072 383236
rect 331912 383180 347788 383236
rect 347844 383180 347854 383236
rect 257842 383068 257852 383124
rect 257908 383068 263788 383124
rect 263844 383068 263854 383124
rect 352706 382956 352716 383012
rect 352772 382956 373548 383012
rect 373604 382956 373614 383012
rect 537618 382956 537628 383012
rect 537684 382956 558908 383012
rect 558964 382956 558974 383012
rect 535938 382844 535948 382900
rect 536004 382844 554204 382900
rect 554260 382844 554270 382900
rect 537730 382732 537740 382788
rect 537796 382732 553532 382788
rect 553588 382732 553598 382788
rect 263778 382620 263788 382676
rect 263844 382620 268072 382676
rect 331912 382620 467852 382676
rect 467908 382620 467918 382676
rect 265010 382060 265020 382116
rect 265076 382060 268072 382116
rect 331912 382060 399196 382116
rect 399252 382060 399262 382116
rect 206098 381500 206108 381556
rect 206164 381500 268072 381556
rect 331912 381500 371308 381556
rect 371364 381500 371374 381556
rect 392242 381276 392252 381332
rect 392308 381276 396732 381332
rect 396788 381276 396798 381332
rect 262994 380940 263004 380996
rect 263060 380940 268072 380996
rect 331912 380940 579628 380996
rect 579684 380940 579694 380996
rect 133522 380716 133532 380772
rect 133588 380716 264908 380772
rect 264964 380716 264974 380772
rect 42242 380604 42252 380660
rect 42308 380604 247772 380660
rect 247828 380604 247838 380660
rect 42914 380492 42924 380548
rect 42980 380492 261436 380548
rect 261492 380492 261502 380548
rect 335234 380492 335244 380548
rect 335300 380492 455420 380548
rect 455476 380492 455486 380548
rect 204866 380380 204876 380436
rect 204932 380380 268072 380436
rect 331912 380380 474684 380436
rect 474740 380380 474750 380436
rect 261202 379820 261212 379876
rect 261268 379820 268072 379876
rect 331912 379820 533372 379876
rect 533428 379820 533438 379876
rect 259522 379260 259532 379316
rect 259588 379260 268072 379316
rect 331912 379260 530012 379316
rect 530068 379260 530078 379316
rect 79762 379036 79772 379092
rect 79828 379036 264796 379092
rect 264852 379036 264862 379092
rect 18162 378924 18172 378980
rect 18228 378924 257852 378980
rect 257908 378924 257918 378980
rect 19730 378812 19740 378868
rect 19796 378812 264572 378868
rect 264628 378812 264638 378868
rect 335122 378812 335132 378868
rect 335188 378812 395052 378868
rect 395108 378812 395118 378868
rect 256162 378700 256172 378756
rect 256228 378700 268072 378756
rect 331912 378700 560252 378756
rect 560308 378700 560318 378756
rect 263778 378140 263788 378196
rect 263844 378140 268072 378196
rect 331912 378140 462812 378196
rect 462868 378140 462878 378196
rect 229506 377580 229516 377636
rect 229572 377580 268072 377636
rect 331912 377580 533484 377636
rect 533540 377580 533550 377636
rect 69682 377132 69692 377188
rect 69748 377132 264684 377188
rect 264740 377132 264750 377188
rect 595560 377160 597000 377384
rect 141026 377020 141036 377076
rect 141092 377020 268072 377076
rect 331912 377020 476252 377076
rect 476308 377020 476318 377076
rect 167570 376460 167580 376516
rect 167636 376460 268072 376516
rect 331912 376460 519148 376516
rect 519204 376460 519214 376516
rect 189074 375900 189084 375956
rect 189140 375900 268072 375956
rect 331912 375900 519932 375956
rect 519988 375900 519998 375956
rect -960 375480 480 375704
rect 336130 375452 336140 375508
rect 336196 375452 458780 375508
rect 458836 375452 458846 375508
rect 197362 375340 197372 375396
rect 197428 375340 268072 375396
rect 331912 375340 461132 375396
rect 461188 375340 461198 375396
rect 192322 374780 192332 374836
rect 192388 374780 268072 374836
rect 331912 374780 400652 374836
rect 400708 374780 400718 374836
rect 142706 374220 142716 374276
rect 142772 374220 268072 374276
rect 331912 374220 493500 374276
rect 493556 374220 493566 374276
rect 130162 373772 130172 373828
rect 130228 373772 263788 373828
rect 263844 373772 263854 373828
rect 188962 373660 188972 373716
rect 189028 373660 268072 373716
rect 331912 373660 517468 373716
rect 517524 373660 517534 373716
rect 187394 373100 187404 373156
rect 187460 373100 268072 373156
rect 331912 373100 498204 373156
rect 498260 373100 498270 373156
rect 195682 372540 195692 372596
rect 195748 372540 268072 372596
rect 331912 372540 467852 372596
rect 467908 372540 467918 372596
rect 76402 372092 76412 372148
rect 76468 372092 263788 372148
rect 263844 372092 263854 372148
rect 192322 371980 192332 372036
rect 192388 371980 268072 372036
rect 331912 371980 464492 372036
rect 464548 371980 464558 372036
rect 205762 371420 205772 371476
rect 205828 371420 268072 371476
rect 331912 371420 503132 371476
rect 503188 371420 503198 371476
rect 187282 370860 187292 370916
rect 187348 370860 268072 370916
rect 331912 370860 407372 370916
rect 407428 370860 407438 370916
rect 264898 370300 264908 370356
rect 264964 370300 268072 370356
rect 331912 370300 336140 370356
rect 336196 370300 336206 370356
rect 263778 369740 263788 369796
rect 263844 369740 268072 369796
rect 331912 369740 335244 369796
rect 335300 369740 335310 369796
rect 127026 369180 127036 369236
rect 127092 369180 268072 369236
rect 331912 369180 457212 369236
rect 457268 369180 457278 369236
rect 334562 368732 334572 368788
rect 334628 368732 394940 368788
rect 394996 368732 395006 368788
rect 103506 368620 103516 368676
rect 103572 368620 268072 368676
rect 331912 368620 455308 368676
rect 455364 368620 455374 368676
rect 127250 368060 127260 368116
rect 127316 368060 268072 368116
rect 331912 368060 404012 368116
rect 404068 368060 404078 368116
rect 100818 367500 100828 367556
rect 100884 367500 268072 367556
rect 331912 367500 457324 367556
rect 457380 367500 457390 367556
rect 334338 367052 334348 367108
rect 334404 367052 402332 367108
rect 402388 367052 402398 367108
rect 107538 366940 107548 366996
rect 107604 366940 268072 366996
rect 331912 366940 398972 366996
rect 399028 366940 399038 366996
rect 126914 366380 126924 366436
rect 126980 366380 268072 366436
rect 331912 366380 457100 366436
rect 457156 366380 457166 366436
rect 100146 365820 100156 365876
rect 100212 365820 268072 365876
rect 331912 365820 412412 365876
rect 412468 365820 412478 365876
rect 334450 365484 334460 365540
rect 334516 365484 396508 365540
rect 396564 365484 396574 365540
rect 393138 365372 393148 365428
rect 393204 365372 459004 365428
rect 459060 365372 459070 365428
rect 126802 365260 126812 365316
rect 126868 365260 268072 365316
rect 331912 365260 456092 365316
rect 456148 365260 456158 365316
rect 127138 364700 127148 364756
rect 127204 364700 268072 364756
rect 331912 364700 334348 364756
rect 334404 364700 334414 364756
rect 143602 364140 143612 364196
rect 143668 364140 268072 364196
rect 331912 364140 393148 364196
rect 393204 364140 393214 364196
rect 595560 363972 597000 364168
rect 393922 363916 393932 363972
rect 393988 363944 597000 363972
rect 393988 363916 595672 363944
rect 257842 363580 257852 363636
rect 257908 363580 268072 363636
rect 331912 363580 335132 363636
rect 335188 363580 335198 363636
rect 263778 363020 263788 363076
rect 263844 363020 268072 363076
rect 331912 363020 334460 363076
rect 334516 363020 334526 363076
rect 18274 362460 18284 362516
rect 18340 362460 268072 362516
rect 331912 362460 334572 362516
rect 334628 362460 334638 362516
rect 335906 362124 335916 362180
rect 335972 362124 351932 362180
rect 351988 362124 351998 362180
rect 335906 362012 335916 362068
rect 335972 362012 394828 362068
rect 394884 362012 394894 362068
rect 18050 361900 18060 361956
rect 18116 361900 268072 361956
rect 331912 361900 392252 361956
rect 392308 361900 392318 361956
rect -960 361396 480 361592
rect -960 361368 8428 361396
rect 392 361340 8428 361368
rect 264674 361340 264684 361396
rect 264740 361340 268072 361396
rect 331912 361340 345212 361396
rect 345268 361340 345278 361396
rect 8372 361284 8428 361340
rect 8372 361228 266364 361284
rect 266420 361228 266430 361284
rect 73042 360780 73052 360836
rect 73108 360780 268072 360836
rect 331912 360780 345212 360836
rect 345268 360780 345278 360836
rect 342626 360332 342636 360388
rect 342692 360332 377580 360388
rect 377636 360332 377646 360388
rect 64866 360220 64876 360276
rect 64932 360220 268072 360276
rect 331912 360220 341852 360276
rect 341908 360220 341918 360276
rect 64642 359660 64652 359716
rect 64708 359660 268072 359716
rect 331912 359660 372204 359716
rect 372260 359660 372270 359716
rect 247762 359100 247772 359156
rect 247828 359100 268072 359156
rect 331912 359100 335916 359156
rect 335972 359100 335982 359156
rect 339266 358652 339276 358708
rect 339332 358652 558908 358708
rect 558964 358652 558974 358708
rect 264786 358540 264796 358596
rect 264852 358540 268072 358596
rect 331912 358540 342636 358596
rect 342692 358540 342702 358596
rect 402322 358428 402332 358484
rect 402388 358428 439516 358484
rect 439572 358428 439582 358484
rect 229506 358316 229516 358372
rect 229572 358316 249452 358372
rect 249508 358316 249518 358372
rect 340274 358316 340284 358372
rect 340340 358316 370860 358372
rect 370916 358316 370926 358372
rect 393138 358316 393148 358372
rect 393204 358316 498204 358372
rect 498260 358316 498270 358372
rect 45602 358204 45612 358260
rect 45668 358204 62188 358260
rect 62244 358204 62254 358260
rect 158834 358204 158844 358260
rect 158900 358204 186396 358260
rect 186452 358204 186462 358260
rect 225474 358204 225484 358260
rect 225540 358204 248556 358260
rect 248612 358204 248622 358260
rect 350242 358204 350252 358260
rect 350308 358204 493500 358260
rect 493556 358204 493566 358260
rect 539186 358204 539196 358260
rect 539252 358204 566972 358260
rect 567028 358204 567038 358260
rect 36194 358092 36204 358148
rect 36260 358092 61292 358148
rect 61348 358092 61358 358148
rect 97458 358092 97468 358148
rect 97524 358092 122668 358148
rect 122724 358092 122734 358148
rect 163538 358092 163548 358148
rect 163604 358092 199052 358148
rect 199108 358092 199118 358148
rect 224802 358092 224812 358148
rect 224868 358092 257964 358148
rect 258020 358092 258030 358148
rect 352706 358092 352716 358148
rect 352772 358092 562940 358148
rect 562996 358092 563006 358148
rect 35522 357980 35532 358036
rect 35588 357980 62972 358036
rect 63028 357980 63038 358036
rect 100818 357980 100828 358036
rect 100884 357980 138572 358036
rect 138628 357980 138638 358036
rect 166226 357980 166236 358036
rect 166292 357980 247996 358036
rect 248052 357980 248062 358036
rect 261426 357980 261436 358036
rect 261492 357980 268072 358036
rect 331912 357980 338492 358036
rect 338548 357980 338558 358036
rect 341842 357980 341852 358036
rect 341908 357980 557564 358036
rect 557620 357980 557630 358036
rect 38882 357868 38892 357924
rect 38948 357868 74732 357924
rect 74788 357868 74798 357924
rect 104178 357868 104188 357924
rect 104244 357868 261660 357924
rect 261716 357868 261726 357924
rect 348674 357868 348684 357924
rect 348740 357868 369516 357924
rect 369572 357868 369582 357924
rect 410722 357868 410732 357924
rect 410788 357868 435484 357924
rect 435540 357868 435550 357924
rect 475458 357868 475468 357924
rect 475524 357868 494844 357924
rect 494900 357868 494910 357924
rect 264562 357420 264572 357476
rect 264628 357420 268072 357476
rect 331912 357420 335916 357476
rect 335972 357420 335982 357476
rect 337138 357084 337148 357140
rect 337204 357084 500220 357140
rect 500276 357084 500286 357140
rect 205650 356860 205660 356916
rect 205716 356860 268072 356916
rect 331912 356860 352716 356916
rect 352772 356860 352782 356916
rect 336914 356748 336924 356804
rect 336980 356748 372876 356804
rect 372932 356748 372942 356804
rect 398962 356748 398972 356804
rect 399028 356748 432124 356804
rect 432180 356748 432190 356804
rect 166898 356636 166908 356692
rect 166964 356636 187292 356692
rect 187348 356636 187358 356692
rect 228162 356636 228172 356692
rect 228228 356636 263788 356692
rect 263844 356636 263854 356692
rect 341954 356636 341964 356692
rect 342020 356636 378252 356692
rect 378308 356636 378318 356692
rect 400642 356636 400652 356692
rect 400708 356636 436156 356692
rect 436212 356636 436222 356692
rect 158162 356524 158172 356580
rect 158228 356524 247772 356580
rect 247828 356524 247838 356580
rect 352370 356524 352380 356580
rect 352436 356524 500892 356580
rect 500948 356524 500958 356580
rect 108210 356412 108220 356468
rect 108276 356412 258076 356468
rect 258132 356412 258142 356468
rect 345426 356412 345436 356468
rect 345492 356412 497532 356468
rect 497588 356412 497598 356468
rect 40898 356300 40908 356356
rect 40964 356300 81452 356356
rect 81508 356300 81518 356356
rect 99474 356300 99484 356356
rect 99540 356300 252924 356356
rect 252980 356300 252990 356356
rect 259522 356300 259532 356356
rect 259588 356300 268072 356356
rect 331912 356300 581308 356356
rect 581364 356300 581374 356356
rect 44258 356188 44268 356244
rect 44324 356188 261324 356244
rect 261380 356188 261390 356244
rect 334338 356188 334348 356244
rect 334404 356188 339276 356244
rect 339332 356188 339342 356244
rect 352146 356188 352156 356244
rect 352212 356188 374220 356244
rect 374276 356188 374286 356244
rect 412402 356188 412412 356244
rect 412468 356188 430780 356244
rect 430836 356188 430846 356244
rect 232194 356076 232204 356132
rect 232260 356076 249564 356132
rect 249620 356076 249630 356132
rect 223346 355964 223356 356020
rect 223412 355964 252812 356020
rect 252868 355964 252878 356020
rect 351922 355964 351932 356020
rect 351988 355964 495628 356020
rect 495684 355964 495694 356020
rect 168914 355852 168924 355908
rect 168980 355852 248332 355908
rect 248388 355852 248398 355908
rect 349234 355852 349244 355908
rect 349300 355852 581420 355908
rect 581476 355852 581486 355908
rect 161522 355740 161532 355796
rect 161588 355740 187516 355796
rect 187572 355740 187582 355796
rect 206658 355740 206668 355796
rect 206724 355740 268072 355796
rect 331912 355740 583100 355796
rect 583156 355740 583166 355796
rect 107538 355628 107548 355684
rect 107604 355628 249788 355684
rect 249844 355628 249854 355684
rect 335122 355628 335132 355684
rect 335188 355628 501116 355684
rect 501172 355628 501182 355684
rect 34850 355516 34860 355572
rect 34916 355516 264572 355572
rect 264628 355516 264638 355572
rect 338594 355516 338604 355572
rect 338660 355516 499548 355572
rect 499604 355516 499614 355572
rect 104850 355404 104860 355460
rect 104916 355404 259644 355460
rect 259700 355404 259710 355460
rect 331884 355404 518252 355460
rect 518308 355404 518318 355460
rect 40226 355292 40236 355348
rect 40292 355292 256284 355348
rect 256340 355292 256350 355348
rect 264786 355180 264796 355236
rect 264852 355180 268072 355236
rect 331884 355208 331940 355404
rect 345314 355292 345324 355348
rect 345380 355292 374892 355348
rect 374948 355292 374958 355348
rect 349234 355180 349244 355236
rect 349300 355180 349310 355236
rect 349244 355012 349300 355180
rect 331884 354956 349300 355012
rect 331884 354648 331940 354956
rect 268044 354564 268100 354648
rect 263788 354508 268100 354564
rect 263788 354228 263844 354508
rect 206210 354172 206220 354228
rect 206276 354172 263844 354228
rect 204754 354060 204764 354116
rect 204820 354060 268072 354116
rect 331912 354060 580412 354116
rect 580468 354060 580478 354116
rect 186386 353948 186396 354004
rect 186452 353948 264460 354004
rect 264516 353948 264526 354004
rect 122658 353836 122668 353892
rect 122724 353836 265356 353892
rect 265412 353836 265422 353892
rect 335234 353836 335244 353892
rect 335300 353836 393148 353892
rect 393204 353836 393214 353892
rect 62178 353724 62188 353780
rect 62244 353724 264908 353780
rect 264964 353724 264974 353780
rect 335458 353724 335468 353780
rect 335524 353724 475468 353780
rect 475524 353724 475534 353780
rect 61282 353612 61292 353668
rect 61348 353612 264684 353668
rect 264740 353612 264750 353668
rect 334450 353612 334460 353668
rect 334516 353612 539196 353668
rect 539252 353612 539262 353668
rect 263778 353500 263788 353556
rect 263844 353500 268072 353556
rect 331912 353500 334348 353556
rect 334404 353500 334414 353556
rect 351026 353052 351036 353108
rect 351092 353052 535164 353108
rect 535220 353052 535230 353108
rect 265122 352940 265132 352996
rect 265188 352940 268072 352996
rect 331912 352940 579628 352996
rect 579684 352940 579694 352996
rect 352594 352828 352604 352884
rect 352660 352828 583212 352884
rect 583268 352828 583278 352884
rect 202962 352604 202972 352660
rect 203028 352604 206668 352660
rect 206724 352604 206734 352660
rect 264562 352380 264572 352436
rect 264628 352380 268072 352436
rect 331912 352380 351036 352436
rect 351092 352380 351102 352436
rect 263330 351820 263340 351876
rect 263396 351820 268072 351876
rect 331912 351820 338492 351876
rect 338548 351820 338558 351876
rect 261202 351260 261212 351316
rect 261268 351260 268072 351316
rect 331912 351260 352604 351316
rect 352660 351260 352670 351316
rect 202850 351036 202860 351092
rect 202916 351036 205660 351092
rect 205716 351036 205726 351092
rect 590482 350924 590492 350980
rect 590548 350952 595672 350980
rect 590548 350924 597000 350952
rect 268044 350308 268100 350728
rect 331912 350700 334460 350756
rect 334516 350700 334526 350756
rect 595560 350728 597000 350924
rect 247884 350252 268100 350308
rect 247884 349720 247940 350252
rect 263778 350140 263788 350196
rect 263844 350140 268072 350196
rect 331912 350140 335356 350196
rect 335412 350140 335422 350196
rect 393372 349972 393428 350392
rect 393362 349916 393372 349972
rect 393428 349916 393438 349972
rect 473218 349692 473228 349748
rect 473284 349692 476056 349748
rect 248546 349580 248556 349636
rect 248612 349580 268072 349636
rect 331912 349580 334460 349636
rect 334516 349580 334526 349636
rect 248322 349020 248332 349076
rect 248388 349020 268072 349076
rect 331912 349020 351932 349076
rect 351988 349020 351998 349076
rect 247986 348572 247996 348628
rect 248052 348572 263788 348628
rect 263844 348572 263854 348628
rect 262882 348460 262892 348516
rect 262948 348460 268072 348516
rect 331912 348460 335468 348516
rect 335524 348460 335534 348516
rect 263778 347900 263788 347956
rect 263844 347900 268072 347956
rect 331912 347900 350364 347956
rect 350420 347900 350430 347956
rect 392 347480 7644 347508
rect -960 347452 7644 347480
rect 7700 347452 7710 347508
rect -960 347256 480 347452
rect 260082 347340 260092 347396
rect 260148 347340 268072 347396
rect 331912 347340 345212 347396
rect 345268 347340 345278 347396
rect 257842 346780 257852 346836
rect 257908 346780 268072 346836
rect 331912 346780 351932 346836
rect 351988 346780 351998 346836
rect 262098 346220 262108 346276
rect 262164 346220 268072 346276
rect 331912 346220 335132 346276
rect 335188 346220 335198 346276
rect 263778 345660 263788 345716
rect 263844 345660 268072 345716
rect 331912 345660 334460 345716
rect 334516 345660 334526 345716
rect 263890 345100 263900 345156
rect 263956 345100 268072 345156
rect 331912 345100 334348 345156
rect 334404 345100 334414 345156
rect 247762 344540 247772 344596
rect 247828 344540 268072 344596
rect 331912 344540 345436 344596
rect 345492 344540 345502 344596
rect 263778 343980 263788 344036
rect 263844 343980 268072 344036
rect 331912 343980 338604 344036
rect 338660 343980 338670 344036
rect 264450 343420 264460 343476
rect 264516 343420 268072 343476
rect 331912 343420 334460 343476
rect 334516 343420 334526 343476
rect 261426 342860 261436 342916
rect 261492 342860 268072 342916
rect 331912 342860 352044 342916
rect 352100 342860 352110 342916
rect 263778 342300 263788 342356
rect 263844 342300 268072 342356
rect 331912 342300 334348 342356
rect 334404 342300 334414 342356
rect 263778 341740 263788 341796
rect 263844 341740 268072 341796
rect 331912 341740 352380 341796
rect 352436 341740 352446 341796
rect 580402 341740 580412 341796
rect 580468 341740 580478 341796
rect 580412 341684 580468 341740
rect 18386 341628 18396 341684
rect 18452 341628 20076 341684
rect 20132 341628 20142 341684
rect 82674 341628 82684 341684
rect 82740 341628 82750 341684
rect 141026 341628 141036 341684
rect 141092 341628 144060 341684
rect 144116 341628 144126 341684
rect 349346 341628 349356 341684
rect 349412 341656 352632 341684
rect 349412 341628 352660 341656
rect 473666 341628 473676 341684
rect 473732 341628 476028 341684
rect 476084 341628 476094 341684
rect 534258 341628 534268 341684
rect 534324 341628 535836 341684
rect 535892 341628 538104 341684
rect 579852 341628 580468 341684
rect 352604 341236 352660 341628
rect 263778 341180 263788 341236
rect 263844 341180 268072 341236
rect 331912 341180 334460 341236
rect 334516 341180 334526 341236
rect 352594 341180 352604 341236
rect 352660 341180 352670 341236
rect 201282 340956 201292 341012
rect 201348 340956 206136 341012
rect 263890 340620 263900 340676
rect 263956 340620 268072 340676
rect 331912 340620 334348 340676
rect 334404 340620 334414 340676
rect 393932 340452 393988 340984
rect 414642 340956 414652 341012
rect 414708 340956 414718 341012
rect 579852 340984 579908 341628
rect 455420 340452 455476 340984
rect 393932 340396 394044 340452
rect 394100 340396 394110 340452
rect 455410 340396 455420 340452
rect 455476 340396 455486 340452
rect 82450 340284 82460 340340
rect 82516 340284 82526 340340
rect 123928 340284 127484 340340
rect 127540 340284 127550 340340
rect 141026 340284 141036 340340
rect 141092 340284 144088 340340
rect 185864 340284 189532 340340
rect 189588 340284 189598 340340
rect 247912 340284 264572 340340
rect 264628 340284 264638 340340
rect 61880 339612 65212 339668
rect 65268 339612 65278 339668
rect 82460 339640 82516 340284
rect 256162 340060 256172 340116
rect 256228 340060 268072 340116
rect 331912 340060 334460 340116
rect 334516 340060 334526 340116
rect 393372 339780 393428 340312
rect 455868 339780 455924 340312
rect 518242 340284 518252 340340
rect 518308 340284 538104 340340
rect 579880 340284 581420 340340
rect 581476 340284 581486 340340
rect 393362 339724 393372 339780
rect 393428 339724 393438 339780
rect 455868 339724 457828 339780
rect 185864 339612 200956 339668
rect 201012 339612 201022 339668
rect 345202 339612 345212 339668
rect 345268 339612 352072 339668
rect 455522 339612 455532 339668
rect 455588 339612 455598 339668
rect 457772 339556 457828 339724
rect 473218 339612 473228 339668
rect 473284 339612 476056 339668
rect 263778 339500 263788 339556
rect 263844 339500 268072 339556
rect 331912 339500 348572 339556
rect 348628 339500 348638 339556
rect 457762 339500 457772 339556
rect 457828 339500 457838 339556
rect 126130 339276 126140 339332
rect 126196 339276 130060 339332
rect 130116 339276 130126 339332
rect 18050 338940 18060 338996
rect 18116 338940 20104 338996
rect 261650 338940 261660 338996
rect 261716 338940 268072 338996
rect 331912 338940 334348 338996
rect 334404 338940 334414 338996
rect 341842 338940 341852 338996
rect 341908 338940 352072 338996
rect 472882 338940 472892 338996
rect 472948 338940 476056 338996
rect 517458 338716 517468 338772
rect 517524 338716 517534 338772
rect 127474 338492 127484 338548
rect 127540 338492 143612 338548
rect 143668 338492 143678 338548
rect 189522 338492 189532 338548
rect 189588 338492 204092 338548
rect 204148 338492 204158 338548
rect 335122 338492 335132 338548
rect 335188 338492 348684 338548
rect 348740 338492 348750 338548
rect 259634 338380 259644 338436
rect 259700 338380 268072 338436
rect 331912 338380 337708 338436
rect 337764 338380 337774 338436
rect 123928 338268 127596 338324
rect 127652 338268 127662 338324
rect 206098 338268 206108 338324
rect 206164 338268 206174 338324
rect 517468 338296 517524 338716
rect 455308 337876 455364 338296
rect 265346 337820 265356 337876
rect 265412 337820 268072 337876
rect 331912 337820 334460 337876
rect 334516 337820 334526 337876
rect 455298 337820 455308 337876
rect 455364 337820 455374 337876
rect 82226 337596 82236 337652
rect 82292 337596 82302 337652
rect 123928 337596 126028 337652
rect 140914 337596 140924 337652
rect 140980 337596 144088 337652
rect 185864 337596 192444 337652
rect 192500 337596 192510 337652
rect 247912 337596 261212 337652
rect 261268 337596 261278 337652
rect 125972 337428 126028 337596
rect 125972 337372 141932 337428
rect 141988 337372 141998 337428
rect 252914 337260 252924 337316
rect 252980 337260 268072 337316
rect 331912 337260 334348 337316
rect 334404 337260 334414 337316
rect 393484 337092 393540 337624
rect 517458 337596 517468 337652
rect 517524 337596 517534 337652
rect 579880 337596 583100 337652
rect 583156 337596 583166 337652
rect 595560 337512 597000 337736
rect 393474 337036 393484 337092
rect 393540 337036 393550 337092
rect 20636 336420 20692 336952
rect 61880 336924 64092 336980
rect 64148 336924 64158 336980
rect 82012 336420 82068 336952
rect 123928 336924 127596 336980
rect 127652 336924 127662 336980
rect 185864 336924 188972 336980
rect 189028 336924 189038 336980
rect 247912 336924 265132 336980
rect 265188 336924 265198 336980
rect 264562 336700 264572 336756
rect 264628 336700 268072 336756
rect 331912 336700 334460 336756
rect 334516 336700 334526 336756
rect 393932 336532 393988 336952
rect 517944 336924 520828 336980
rect 520884 336924 520894 336980
rect 579880 336924 581308 336980
rect 581364 336924 581374 336980
rect 455298 336812 455308 336868
rect 455364 336812 455374 336868
rect 393932 336476 396508 336532
rect 20626 336364 20636 336420
rect 20692 336364 20702 336420
rect 80546 336364 80556 336420
rect 80612 336364 82068 336420
rect 396452 336364 396508 336476
rect 396564 336364 396574 336420
rect 18274 336252 18284 336308
rect 18340 336252 20104 336308
rect 61880 336252 64204 336308
rect 64260 336252 64270 336308
rect 185864 336252 195804 336308
rect 195860 336252 195870 336308
rect 204866 336252 204876 336308
rect 204932 336252 206136 336308
rect 247912 336252 264796 336308
rect 264852 336252 264862 336308
rect 455308 336280 455364 336812
rect 249778 336140 249788 336196
rect 249844 336140 268072 336196
rect 331912 336140 334460 336196
rect 334516 336140 334526 336196
rect 393932 336084 393988 336280
rect 393932 336028 394828 336084
rect 394884 336028 394894 336084
rect 61880 335580 64764 335636
rect 64820 335580 64830 335636
rect 185864 335580 195692 335636
rect 195748 335580 195758 335636
rect 264002 335580 264012 335636
rect 264068 335580 268072 335636
rect 331912 335580 351148 335636
rect 351204 335580 351214 335636
rect 455522 335580 455532 335636
rect 455588 335580 455598 335636
rect 517944 335580 519148 335636
rect 519204 335580 519214 335636
rect 260306 335020 260316 335076
rect 260372 335020 268072 335076
rect 331912 335020 334460 335076
rect 334516 335020 334526 335076
rect 18386 334908 18396 334964
rect 18452 334908 20104 334964
rect 258066 334460 258076 334516
rect 258132 334460 268072 334516
rect 331912 334460 334460 334516
rect 334516 334460 334526 334516
rect 393932 334404 393988 334936
rect 461122 334908 461132 334964
rect 461188 334908 476056 334964
rect 579880 334908 582988 334964
rect 583044 334908 583054 334964
rect 393932 334348 394996 334404
rect 394940 334292 394996 334348
rect 206210 334236 206220 334292
rect 206276 334236 206286 334292
rect 247912 334236 251020 334292
rect 251076 334236 251086 334292
rect 264898 333900 264908 333956
rect 264964 333900 268072 333956
rect 331912 333900 340396 333956
rect 340452 333900 340462 333956
rect 393372 333732 393428 334264
rect 394930 334236 394940 334292
rect 394996 334236 395006 334292
rect 399746 334236 399756 334292
rect 399812 334236 414120 334292
rect 535154 334236 535164 334292
rect 535220 334236 538104 334292
rect 393362 333676 393372 333732
rect 393428 333676 393438 333732
rect 123928 333564 126140 333620
rect 126196 333564 126206 333620
rect 185864 333564 189084 333620
rect 189140 333564 189150 333620
rect 202962 333564 202972 333620
rect 203028 333564 206136 333620
rect 455634 333564 455644 333620
rect 455700 333564 455710 333620
rect 473106 333564 473116 333620
rect 473172 333564 476056 333620
rect 534258 333564 534268 333620
rect 534324 333564 538104 333620
rect 579618 333564 579628 333620
rect 579684 333564 579694 333620
rect -960 333144 480 333368
rect 264674 333340 264684 333396
rect 264740 333340 268072 333396
rect 331912 333340 334460 333396
rect 334516 333340 334526 333396
rect 20066 332892 20076 332948
rect 20132 332892 20142 332948
rect 61880 332892 64652 332948
rect 64708 332892 64718 332948
rect 123928 332892 127596 332948
rect 127652 332892 127662 332948
rect 185864 332892 192332 332948
rect 192388 332892 192398 332948
rect 204754 332892 204764 332948
rect 204820 332892 206136 332948
rect 455644 332920 455700 333564
rect 456082 333452 456092 333508
rect 456148 333452 473228 333508
rect 473284 333452 473294 333508
rect 263778 332780 263788 332836
rect 263844 332780 268072 332836
rect 331912 332780 352268 332836
rect 352324 332780 352334 332836
rect 393932 332724 393988 332920
rect 517944 332892 521052 332948
rect 521108 332892 521118 332948
rect 523282 332892 523292 332948
rect 523348 332892 538104 332948
rect 393932 332668 396844 332724
rect 396900 332668 396910 332724
rect 18162 332220 18172 332276
rect 18228 332220 20104 332276
rect 61880 332220 69692 332276
rect 69748 332220 69758 332276
rect 185864 332220 205772 332276
rect 205828 332220 205838 332276
rect 247912 332220 261324 332276
rect 261380 332220 261390 332276
rect 264898 332220 264908 332276
rect 264964 332220 268072 332276
rect 331912 332220 352156 332276
rect 352212 332220 352222 332276
rect 393922 332220 393932 332276
rect 393988 332220 414120 332276
rect 455298 332220 455308 332276
rect 455364 332220 455374 332276
rect 517944 332220 520940 332276
rect 520996 332220 521006 332276
rect 523282 332220 523292 332276
rect 523348 332220 538104 332276
rect 579628 331716 579684 332248
rect 263890 331660 263900 331716
rect 263956 331660 268072 331716
rect 331912 331660 334460 331716
rect 334516 331660 334526 331716
rect 579618 331660 579628 331716
rect 579684 331660 579694 331716
rect 61880 331548 64204 331604
rect 64260 331548 64270 331604
rect 185864 331548 189420 331604
rect 189476 331548 189486 331604
rect 80546 331436 80556 331492
rect 80612 331436 81452 331492
rect 81508 331436 81518 331492
rect 455308 331268 455364 331576
rect 455298 331212 455308 331268
rect 455364 331212 455374 331268
rect 263778 331100 263788 331156
rect 263844 331100 268072 331156
rect 331912 331100 345324 331156
rect 345380 331100 345390 331156
rect 203074 330876 203084 330932
rect 203140 330876 206136 330932
rect 395602 330876 395612 330932
rect 395668 330876 396508 330932
rect 396564 330876 396574 330932
rect 535042 330876 535052 330932
rect 535108 330876 538104 330932
rect 205986 330652 205996 330708
rect 206052 330652 206164 330708
rect 82012 329700 82068 330232
rect 123928 330204 126812 330260
rect 126868 330204 126878 330260
rect 206108 330232 206164 330652
rect 263778 330540 263788 330596
rect 263844 330540 268072 330596
rect 331912 330540 341964 330596
rect 342020 330540 342030 330596
rect 247912 330204 251916 330260
rect 251972 330204 251982 330260
rect 338482 330204 338492 330260
rect 338548 330204 352072 330260
rect 256274 329980 256284 330036
rect 256340 329980 268072 330036
rect 331912 329980 334460 330036
rect 334516 329980 334526 330036
rect 80434 329644 80444 329700
rect 80500 329644 82068 329700
rect 393932 329700 393988 330232
rect 407362 330204 407372 330260
rect 407428 330204 414120 330260
rect 393932 329644 394828 329700
rect 394884 329644 394894 329700
rect 82012 329364 82068 329560
rect 123928 329532 127596 329588
rect 127652 329532 127662 329588
rect 202850 329532 202860 329588
rect 202916 329532 206136 329588
rect 247912 329532 259532 329588
rect 259588 329532 259598 329588
rect 393250 329532 393260 329588
rect 393316 329532 393326 329588
rect 261314 329420 261324 329476
rect 261380 329420 268072 329476
rect 331912 329420 344428 329476
rect 344484 329420 344494 329476
rect 80546 329308 80556 329364
rect 80612 329308 82068 329364
rect 185864 328860 197372 328916
rect 197428 328860 197438 328916
rect 263890 328860 263900 328916
rect 263956 328860 268072 328916
rect 331912 328860 338604 328916
rect 338660 328860 338670 328916
rect 455522 328860 455532 328916
rect 455588 328860 455598 328916
rect 455410 328636 455420 328692
rect 455476 328636 455486 328692
rect 264674 328300 264684 328356
rect 264740 328300 268072 328356
rect 331912 328300 350588 328356
rect 350644 328300 350654 328356
rect 455420 328216 455476 328636
rect 263778 327740 263788 327796
rect 263844 327740 268072 327796
rect 331912 327740 334460 327796
rect 334516 327740 334526 327796
rect 258066 327180 258076 327236
rect 258132 327180 268072 327236
rect 331912 327180 334460 327236
rect 334516 327180 334526 327236
rect 264562 326620 264572 326676
rect 264628 326620 268072 326676
rect 331912 326620 350252 326676
rect 350308 326620 350318 326676
rect 261314 326060 261324 326116
rect 261380 326060 268072 326116
rect 331912 326060 334348 326116
rect 334404 326060 334414 326116
rect 263778 325500 263788 325556
rect 263844 325500 268072 325556
rect 331912 325500 334460 325556
rect 334516 325500 334526 325556
rect 579880 325500 583212 325556
rect 583268 325500 583278 325556
rect 251010 324940 251020 324996
rect 251076 324940 268072 324996
rect 331912 324940 341852 324996
rect 341908 324940 341918 324996
rect 587234 324492 587244 324548
rect 587300 324520 595672 324548
rect 587300 324492 597000 324520
rect 249554 324380 249564 324436
rect 249620 324380 268072 324436
rect 331912 324380 334460 324436
rect 334516 324380 334526 324436
rect 595560 324296 597000 324492
rect 263778 323820 263788 323876
rect 263844 323820 268072 323876
rect 331912 323820 334460 323876
rect 334516 323820 334526 323876
rect 257954 323260 257964 323316
rect 258020 323260 268072 323316
rect 331912 323260 345324 323316
rect 345380 323260 345390 323316
rect 259522 322700 259532 322756
rect 259588 322700 268072 322756
rect 331912 322700 334348 322756
rect 334404 322700 334414 322756
rect 261202 322140 261212 322196
rect 261268 322140 268072 322196
rect 331912 322140 348684 322196
rect 348740 322140 348750 322196
rect 251906 321580 251916 321636
rect 251972 321580 268072 321636
rect 331912 321580 334460 321636
rect 334516 321580 334526 321636
rect 252802 321020 252812 321076
rect 252868 321020 268072 321076
rect 331912 321020 335468 321076
rect 335524 321020 335534 321076
rect 261314 320460 261324 320516
rect 261380 320460 268072 320516
rect 331912 320460 351932 320516
rect 351988 320460 351998 320516
rect 247762 319900 247772 319956
rect 247828 319900 268072 319956
rect 331912 319900 334460 319956
rect 334516 319900 334526 319956
rect 249442 319340 249452 319396
rect 249508 319340 268072 319396
rect 331912 319340 350476 319396
rect 350532 319340 350542 319396
rect -960 319060 480 319256
rect 140914 319116 140924 319172
rect 140980 319116 142828 319172
rect 142884 319116 142894 319172
rect -960 319032 15932 319060
rect 392 319004 15932 319032
rect 15988 319004 15998 319060
rect 249442 318780 249452 318836
rect 249508 318780 268072 318836
rect 331912 318780 334460 318836
rect 334516 318780 334526 318836
rect 456866 318444 456876 318500
rect 456932 318444 473116 318500
rect 473172 318444 473182 318500
rect 188962 318332 188972 318388
rect 189028 318332 204988 318388
rect 205044 318332 205054 318388
rect 335682 318332 335692 318388
rect 335748 318332 350252 318388
rect 350308 318332 350318 318388
rect 456194 318332 456204 318388
rect 456260 318332 472892 318388
rect 472948 318332 472958 318388
rect 247986 318220 247996 318276
rect 248052 318220 268072 318276
rect 331912 318220 341852 318276
rect 341908 318220 341918 318276
rect 248546 317660 248556 317716
rect 248612 317660 268072 317716
rect 331912 317660 352156 317716
rect 352212 317660 352222 317716
rect 517580 317548 520828 317604
rect 520884 317548 520894 317604
rect 268044 317044 268100 317128
rect 204978 316988 204988 317044
rect 205044 316988 268100 317044
rect 331884 317044 331940 317128
rect 517580 317044 517636 317548
rect 331884 316988 517636 317044
rect 142818 316540 142828 316596
rect 142884 316540 268072 316596
rect 331912 316540 519148 316596
rect 519204 316540 519214 316596
rect 204082 315980 204092 316036
rect 204148 315980 268072 316036
rect 331912 315980 335244 316036
rect 335300 315980 335310 316036
rect 187282 315420 187292 315476
rect 187348 315420 268072 315476
rect 331912 315420 456876 315476
rect 456932 315420 456942 315476
rect 80434 314636 80444 314692
rect 80500 314636 161308 314692
rect 161364 314636 161374 314692
rect 166226 314636 166236 314692
rect 166292 314636 262892 314692
rect 262948 314636 262958 314692
rect 163538 314524 163548 314580
rect 163604 314524 248556 314580
rect 248612 314524 248622 314580
rect 260988 314524 261436 314580
rect 261492 314524 261502 314580
rect 225474 314412 225484 314468
rect 225540 314412 259532 314468
rect 259588 314412 259598 314468
rect 260988 314356 261044 314524
rect 268044 314468 268100 314888
rect 331912 314860 456092 314916
rect 456148 314860 456158 314916
rect 335346 314636 335356 314692
rect 335412 314636 561036 314692
rect 561092 314636 561102 314692
rect 351922 314524 351932 314580
rect 351988 314524 500892 314580
rect 500948 314524 500958 314580
rect 141026 314300 141036 314356
rect 141092 314300 261044 314356
rect 261100 314412 268100 314468
rect 345202 314412 345212 314468
rect 345268 314412 493500 314468
rect 493556 314412 493566 314468
rect 261100 314244 261156 314412
rect 261426 314300 261436 314356
rect 261492 314300 268072 314356
rect 331912 314300 517468 314356
rect 517524 314300 517534 314356
rect 187506 314188 187516 314244
rect 187572 314188 261156 314244
rect 334450 314188 334460 314244
rect 334516 314188 404796 314244
rect 404852 314188 404862 314244
rect 44258 314076 44268 314132
rect 44324 314076 258076 314132
rect 258132 314076 258142 314132
rect 350578 314076 350588 314132
rect 350644 314076 359436 314132
rect 359492 314076 359502 314132
rect 562902 314076 562940 314132
rect 562996 314076 563006 314132
rect 56354 313964 56364 314020
rect 56420 313964 261324 314020
rect 261380 313964 261390 314020
rect 350354 313964 350364 314020
rect 350420 313964 499772 314020
rect 499828 313964 499838 314020
rect 100146 313852 100156 313908
rect 100212 313852 256172 313908
rect 256228 313852 256238 313908
rect 352034 313852 352044 313908
rect 352100 313852 496188 313908
rect 496244 313852 496254 313908
rect 160178 313740 160188 313796
rect 160244 313740 249452 313796
rect 249508 313740 249518 313796
rect 268044 313684 268100 313768
rect 331912 313740 337148 313796
rect 337204 313740 337214 313796
rect 340386 313740 340396 313796
rect 340452 313740 444220 313796
rect 444276 313740 444286 313796
rect 205762 313628 205772 313684
rect 205828 313628 268100 313684
rect 348562 313628 348572 313684
rect 348628 313628 434812 313684
rect 434868 313628 434878 313684
rect 341842 313516 341852 313572
rect 341908 313516 499548 313572
rect 499604 313516 499614 313572
rect 352258 313404 352268 313460
rect 352324 313404 374220 313460
rect 374276 313404 374286 313460
rect 126802 313292 126812 313348
rect 126868 313292 198156 313348
rect 198212 313292 198222 313348
rect 335458 313292 335468 313348
rect 335524 313292 558124 313348
rect 558180 313292 558190 313348
rect 199042 313180 199052 313236
rect 199108 313180 268072 313236
rect 331912 313180 456204 313236
rect 456260 313180 456270 313236
rect 200946 312620 200956 312676
rect 201012 312620 268072 312676
rect 331912 312620 335692 312676
rect 335748 312620 335758 312676
rect 167570 312396 167580 312452
rect 167636 312396 261436 312452
rect 261492 312396 261502 312452
rect 164210 312284 164220 312340
rect 164276 312284 257852 312340
rect 257908 312284 257918 312340
rect 345314 312284 345324 312340
rect 345380 312284 557788 312340
rect 557844 312284 557854 312340
rect 168914 312172 168924 312228
rect 168980 312172 247996 312228
rect 248052 312172 248062 312228
rect 350466 312172 350476 312228
rect 350532 312172 562268 312228
rect 562324 312172 562334 312228
rect 80546 312060 80556 312116
rect 80612 312060 268072 312116
rect 331912 312060 436156 312116
rect 436212 312060 436222 312116
rect 221442 311948 221452 312004
rect 221508 311948 261212 312004
rect 261268 311948 261278 312004
rect 348674 311948 348684 312004
rect 348740 311948 553532 312004
rect 553588 311948 553598 312004
rect 224130 311836 224140 311892
rect 224196 311836 247772 311892
rect 247828 311836 247838 311892
rect 404786 311836 404796 311892
rect 404852 311836 554876 311892
rect 554932 311836 554942 311892
rect 352146 311724 352156 311780
rect 352212 311724 496860 311780
rect 496916 311724 496926 311780
rect 104850 311612 104860 311668
rect 104916 311612 166236 311668
rect 166292 311612 166302 311668
rect 338482 311612 338492 311668
rect 338548 311612 560924 311668
rect 560980 311612 560990 311668
rect 161298 311500 161308 311556
rect 161364 311500 268072 311556
rect 331912 311500 437500 311556
rect 437556 311500 437566 311556
rect 595560 311108 597000 311304
rect 474562 311052 474572 311108
rect 474628 311080 597000 311108
rect 474628 311052 595672 311080
rect 138562 310940 138572 310996
rect 138628 310940 268072 310996
rect 331912 310940 398972 310996
rect 399028 310940 399038 310996
rect 143602 310380 143612 310436
rect 143668 310380 268072 310436
rect 331912 310380 400652 310436
rect 400708 310380 400718 310436
rect 166226 309820 166236 309876
rect 166292 309820 268072 309876
rect 331912 309820 402332 309876
rect 402388 309820 402398 309876
rect 198146 309260 198156 309316
rect 198212 309260 268072 309316
rect 331912 309260 430108 309316
rect 430164 309260 430174 309316
rect 104178 308700 104188 308756
rect 104244 308700 268072 308756
rect 331912 308700 433468 308756
rect 433524 308700 433534 308756
rect 69682 308252 69692 308308
rect 69748 308252 263788 308308
rect 263844 308252 263854 308308
rect 81442 308140 81452 308196
rect 81508 308140 268072 308196
rect 331912 308140 410732 308196
rect 410788 308140 410798 308196
rect 141922 307580 141932 307636
rect 141988 307580 268072 307636
rect 331912 307580 393932 307636
rect 393988 307580 393998 307636
rect 101490 307020 101500 307076
rect 101556 307020 268072 307076
rect 331912 307020 412412 307076
rect 412468 307020 412478 307076
rect 99474 306460 99484 306516
rect 99540 306460 268072 306516
rect 331912 306460 430780 306516
rect 430836 306460 430846 306516
rect 106194 305900 106204 305956
rect 106260 305900 268072 305956
rect 331912 305900 457772 305956
rect 457828 305900 457838 305956
rect 38882 305340 38892 305396
rect 38948 305340 268072 305396
rect 331912 305340 345212 305396
rect 345268 305340 345278 305396
rect -960 304948 480 305144
rect -960 304920 266588 304948
rect 392 304892 266588 304920
rect 266644 304892 266654 304948
rect 64754 304780 64764 304836
rect 64820 304780 268072 304836
rect 331912 304780 336924 304836
rect 336980 304780 336990 304836
rect 263778 304220 263788 304276
rect 263844 304220 268072 304276
rect 331912 304220 376236 304276
rect 376292 304220 376302 304276
rect 64642 303660 64652 303716
rect 64708 303660 268072 303716
rect 331912 303660 373548 303716
rect 373604 303660 373614 303716
rect 81442 303100 81452 303156
rect 81508 303100 268072 303156
rect 331912 303100 370188 303156
rect 370244 303100 370254 303156
rect 43586 302540 43596 302596
rect 43652 302540 268072 302596
rect 331912 302540 396844 302596
rect 396900 302540 396910 302596
rect 18274 301980 18284 302036
rect 18340 301980 268072 302036
rect 331912 301980 372204 302036
rect 372260 301980 372270 302036
rect 62962 301420 62972 301476
rect 63028 301420 268072 301476
rect 331912 301420 340284 301476
rect 340340 301420 340350 301476
rect 36866 300860 36876 300916
rect 36932 300860 268072 300916
rect 331912 300860 341852 300916
rect 341908 300860 341918 300916
rect 74722 300300 74732 300356
rect 74788 300300 268072 300356
rect 331912 300300 335132 300356
rect 335188 300300 335198 300356
rect 18162 299740 18172 299796
rect 18228 299740 268072 299796
rect 331912 299740 338492 299796
rect 338548 299740 338558 299796
rect 18386 299180 18396 299236
rect 18452 299180 268072 299236
rect 331912 299180 395612 299236
rect 395668 299180 395678 299236
rect 264562 298620 264572 298676
rect 264628 298620 268072 298676
rect 331912 298620 400652 298676
rect 400708 298620 400718 298676
rect 263890 298060 263900 298116
rect 263956 298060 268072 298116
rect 331912 298060 334460 298116
rect 334516 298060 334526 298116
rect 595560 297864 597000 298088
rect 263778 297500 263788 297556
rect 263844 297500 268072 297556
rect 331912 297500 334348 297556
rect 334404 297500 334414 297556
rect 257842 296940 257852 296996
rect 257908 296940 268072 296996
rect 331912 296940 563724 296996
rect 563780 296940 563790 296996
rect 225922 296604 225932 296660
rect 225988 296604 263788 296660
rect 263844 296604 263854 296660
rect 4498 296492 4508 296548
rect 4564 296492 267932 296548
rect 267988 296492 267998 296548
rect 334450 296492 334460 296548
rect 334516 296492 504812 296548
rect 504868 296492 504878 296548
rect 228834 296380 228844 296436
rect 228900 296380 268072 296436
rect 331912 296380 518252 296436
rect 518308 296380 518318 296436
rect 202962 295820 202972 295876
rect 203028 295820 268072 295876
rect 331912 295820 560364 295876
rect 560420 295820 560430 295876
rect 224802 295260 224812 295316
rect 224868 295260 268072 295316
rect 331912 295260 583548 295316
rect 583604 295260 583614 295316
rect 230850 294812 230860 294868
rect 230916 294812 263900 294868
rect 263956 294812 263966 294868
rect 334338 294812 334348 294868
rect 334404 294812 499772 294868
rect 499828 294812 499838 294868
rect 203074 294700 203084 294756
rect 203140 294700 268072 294756
rect 331912 294700 582092 294756
rect 582148 294700 582158 294756
rect 224130 294140 224140 294196
rect 224196 294140 268072 294196
rect 331912 294140 580412 294196
rect 580468 294140 580478 294196
rect 204754 293580 204764 293636
rect 204820 293580 268072 293636
rect 331912 293580 581308 293636
rect 581364 293580 581374 293636
rect 206098 293020 206108 293076
rect 206164 293020 268072 293076
rect 331912 293020 523292 293076
rect 523348 293020 523358 293076
rect 252802 292460 252812 292516
rect 252868 292460 268072 292516
rect 331912 292460 580524 292516
rect 580580 292460 580590 292516
rect 232866 291900 232876 291956
rect 232932 291900 268072 291956
rect 331912 291900 430108 291956
rect 430164 291900 430174 291956
rect 204866 291340 204876 291396
rect 204932 291340 268072 291396
rect 331912 291340 502348 291396
rect 502404 291340 502414 291396
rect -960 290808 480 291032
rect 263778 290780 263788 290836
rect 263844 290780 268072 290836
rect 331912 290780 335916 290836
rect 335972 290780 335982 290836
rect 189186 290220 189196 290276
rect 189252 290220 268072 290276
rect 331912 290220 449372 290276
rect 449428 290220 449438 290276
rect 140914 289772 140924 289828
rect 140980 289772 263788 289828
rect 263844 289772 263854 289828
rect 335906 289772 335916 289828
rect 335972 289772 517468 289828
rect 517524 289772 517534 289828
rect 518242 289772 518252 289828
rect 518308 289772 559468 289828
rect 559524 289772 559534 289828
rect 187282 289660 187292 289716
rect 187348 289660 268072 289716
rect 331912 289660 517580 289716
rect 517636 289660 517646 289716
rect 188962 289100 188972 289156
rect 189028 289100 268072 289156
rect 331912 289100 519148 289156
rect 519204 289100 519214 289156
rect 249666 288540 249676 288596
rect 249732 288540 268072 288596
rect 331912 288540 340284 288596
rect 340340 288540 340350 288596
rect 45042 288204 45052 288260
rect 45108 288204 259532 288260
rect 259588 288204 259598 288260
rect 504802 288204 504812 288260
rect 504868 288204 556108 288260
rect 556164 288204 556174 288260
rect 334450 288092 334460 288148
rect 334516 288092 351932 288148
rect 351988 288092 351998 288148
rect 499762 288092 499772 288148
rect 499828 288092 561708 288148
rect 561764 288092 561774 288148
rect 200722 287980 200732 288036
rect 200788 287980 268072 288036
rect 331912 287980 498876 288036
rect 498932 287980 498942 288036
rect 166898 287868 166908 287924
rect 166964 287868 247772 287924
rect 247828 287868 247838 287924
rect 334450 287868 334460 287924
rect 334516 287868 334526 287924
rect 334460 287812 334516 287868
rect 98802 287756 98812 287812
rect 98868 287756 122668 287812
rect 122724 287756 122734 287812
rect 162866 287756 162876 287812
rect 162932 287756 248108 287812
rect 248164 287756 248174 287812
rect 331884 287756 334516 287812
rect 341842 287756 341852 287812
rect 341908 287756 376236 287812
rect 376292 287756 376302 287812
rect 105522 287644 105532 287700
rect 105588 287644 258636 287700
rect 258692 287644 258702 287700
rect 98130 287532 98140 287588
rect 98196 287532 256172 287588
rect 256228 287532 256238 287588
rect 40226 287420 40236 287476
rect 40292 287420 143612 287476
rect 143668 287420 143678 287476
rect 169586 287420 169596 287476
rect 169652 287420 268072 287476
rect 331884 287448 331940 287756
rect 350242 287644 350252 287700
rect 350308 287644 436828 287700
rect 436884 287644 436894 287700
rect 342066 287532 342076 287588
rect 342132 287532 438732 287588
rect 438788 287532 438798 287588
rect 477138 287532 477148 287588
rect 477204 287532 501564 287588
rect 501620 287532 501630 287588
rect 350466 287420 350476 287476
rect 350532 287420 498204 287476
rect 498260 287420 498270 287476
rect 223458 287308 223468 287364
rect 223524 287308 225932 287364
rect 225988 287308 225998 287364
rect 228162 287308 228172 287364
rect 228228 287308 252924 287364
rect 252980 287308 252990 287364
rect 338594 287308 338604 287364
rect 338660 287308 554428 287364
rect 554484 287308 554494 287364
rect 170930 286860 170940 286916
rect 170996 286860 268072 286916
rect 331912 286860 352716 286916
rect 352772 286860 352782 286916
rect 335122 286412 335132 286468
rect 335188 286412 477148 286468
rect 477204 286412 477214 286468
rect 502338 286412 502348 286468
rect 502404 286412 583100 286468
rect 583156 286412 583166 286468
rect 168914 286300 168924 286356
rect 168980 286300 268072 286356
rect 331912 286300 500220 286356
rect 500276 286300 500286 286356
rect 164210 286076 164220 286132
rect 164276 286076 258076 286132
rect 258132 286076 258142 286132
rect 106194 285964 106204 286020
rect 106260 285964 249452 286020
rect 249508 285964 249518 286020
rect 258188 285964 261212 286020
rect 261268 285964 261278 286020
rect 352258 285964 352268 286020
rect 352324 285964 375564 286020
rect 375620 285964 375630 286020
rect 102162 285852 102172 285908
rect 102228 285852 256284 285908
rect 256340 285852 256350 285908
rect 258188 285796 258244 285964
rect 41906 285740 41916 285796
rect 41972 285740 258244 285796
rect 258412 285852 261492 285908
rect 348674 285852 348684 285908
rect 348740 285852 433468 285908
rect 433524 285852 433534 285908
rect 258412 285684 258468 285852
rect 261436 285796 261492 285852
rect 261426 285740 261436 285796
rect 261492 285740 261502 285796
rect 263778 285740 263788 285796
rect 263844 285740 268072 285796
rect 331912 285740 464492 285796
rect 464548 285740 464558 285796
rect 475458 285740 475468 285796
rect 475524 285740 500892 285796
rect 500948 285740 500958 285796
rect 41346 285628 41356 285684
rect 41412 285628 258468 285684
rect 259522 285628 259532 285684
rect 259588 285628 264572 285684
rect 264628 285628 264638 285684
rect 338706 285628 338716 285684
rect 338772 285628 368844 285684
rect 368900 285628 368910 285684
rect 369628 285628 499548 285684
rect 499604 285628 499614 285684
rect 369628 285236 369684 285628
rect 197362 285180 197372 285236
rect 197428 285180 268072 285236
rect 331912 285180 369684 285236
rect 144050 284844 144060 284900
rect 144116 284844 261212 284900
rect 261268 284844 261278 284900
rect 449362 284844 449372 284900
rect 449428 284844 521052 284900
rect 521108 284844 521118 284900
rect 160850 284732 160860 284788
rect 160916 284732 262892 284788
rect 262948 284732 262958 284788
rect 263116 284732 268100 284788
rect 430098 284732 430108 284788
rect 430164 284732 535164 284788
rect 535220 284732 535230 284788
rect 263116 284676 263172 284732
rect 205762 284620 205772 284676
rect 205828 284620 263172 284676
rect 268044 284648 268100 284732
rect 595560 284676 597000 284872
rect 331884 284564 331940 284648
rect 333554 284620 333564 284676
rect 333620 284648 597000 284676
rect 333620 284620 595672 284648
rect 102834 284508 102844 284564
rect 102900 284508 249564 284564
rect 249620 284508 249630 284564
rect 331884 284508 473116 284564
rect 473172 284508 473182 284564
rect 101490 284396 101500 284452
rect 101556 284396 252812 284452
rect 252868 284396 252878 284452
rect 261202 284396 261212 284452
rect 261268 284396 268100 284452
rect 352146 284396 352156 284452
rect 352212 284396 376908 284452
rect 376964 284396 376974 284452
rect 37538 284284 37548 284340
rect 37604 284284 192332 284340
rect 192388 284284 192398 284340
rect 42242 284172 42252 284228
rect 42308 284172 264908 284228
rect 264964 284172 264974 284228
rect 268044 284088 268100 284396
rect 345314 284284 345324 284340
rect 345380 284284 434812 284340
rect 434868 284284 434878 284340
rect 336018 284172 336028 284228
rect 336084 284172 432796 284228
rect 432852 284172 432862 284228
rect 331912 284060 342636 284116
rect 342692 284060 342702 284116
rect 204082 283500 204092 283556
rect 204148 283500 268072 283556
rect 331912 283500 475468 283556
rect 475524 283500 475534 283556
rect 143602 283276 143612 283332
rect 143668 283276 265020 283332
rect 265076 283276 265086 283332
rect 142706 283164 142716 283220
rect 142772 283164 263788 283220
rect 263844 283164 263854 283220
rect 342626 283164 342636 283220
rect 342692 283164 472892 283220
rect 472948 283164 472958 283220
rect 473106 283164 473116 283220
rect 473172 283164 520828 283220
rect 520884 283164 520894 283220
rect 122658 283052 122668 283108
rect 122724 283052 264572 283108
rect 264628 283052 264638 283108
rect 352706 283052 352716 283108
rect 352772 283052 520940 283108
rect 520996 283052 521006 283108
rect 523282 283052 523292 283108
rect 523348 283052 583212 283108
rect 583268 283052 583278 283108
rect 138562 282940 138572 282996
rect 138628 282940 268072 282996
rect 331912 282940 456988 282996
rect 457044 282940 457054 282996
rect 80322 282380 80332 282436
rect 80388 282380 268072 282436
rect 331912 282380 455308 282436
rect 455364 282380 455374 282436
rect 136882 281820 136892 281876
rect 136948 281820 268072 281876
rect 331912 281820 456092 281876
rect 456148 281820 456158 281876
rect 130274 281596 130284 281652
rect 130340 281596 268100 281652
rect 334450 281596 334460 281652
rect 334516 281596 458780 281652
rect 458836 281596 458846 281652
rect 82002 281484 82012 281540
rect 82068 281484 255388 281540
rect 255332 281092 255388 281484
rect 268044 281288 268100 281596
rect 349412 281484 457772 281540
rect 457828 281484 457838 281540
rect 331912 281260 345212 281316
rect 345268 281260 345278 281316
rect 349412 281092 349468 281484
rect 255332 281036 268100 281092
rect 268044 280728 268100 281036
rect 331884 281036 349468 281092
rect 331884 280728 331940 281036
rect 258626 280140 258636 280196
rect 258692 280140 268072 280196
rect 331912 280140 348572 280196
rect 348628 280140 348638 280196
rect 263778 279580 263788 279636
rect 263844 279580 268072 279636
rect 331912 279580 334460 279636
rect 334516 279580 334526 279636
rect 455420 279412 455476 279832
rect 455410 279356 455420 279412
rect 455476 279356 455486 279412
rect 204754 279132 204764 279188
rect 204820 279132 206136 279188
rect 263330 279020 263340 279076
rect 263396 279020 268072 279076
rect 331912 279020 336028 279076
rect 336084 279020 336094 279076
rect 257954 278460 257964 278516
rect 258020 278460 268072 278516
rect 331912 278460 334460 278516
rect 334516 278460 334526 278516
rect 517944 278460 520828 278516
rect 520884 278460 520894 278516
rect 256274 277900 256284 277956
rect 256340 277900 268072 277956
rect 331912 277900 348684 277956
rect 348740 277900 348750 277956
rect 262098 277340 262108 277396
rect 262164 277340 268072 277396
rect 331912 277340 342188 277396
rect 342244 277340 342254 277396
rect 61880 277116 64204 277172
rect 64260 277116 64270 277172
rect 455298 277116 455308 277172
rect 455364 277116 455374 277172
rect -960 276724 480 276920
rect 263778 276780 263788 276836
rect 263844 276780 268072 276836
rect 331912 276780 334460 276836
rect 334516 276780 334526 276836
rect -960 276696 19292 276724
rect 392 276668 19292 276696
rect 19348 276668 19358 276724
rect 249554 276220 249564 276276
rect 249620 276220 268072 276276
rect 331912 276220 345324 276276
rect 345380 276220 345390 276276
rect 262210 275660 262220 275716
rect 262276 275660 268072 275716
rect 331912 275660 334348 275716
rect 334404 275660 334414 275716
rect 249442 275100 249452 275156
rect 249508 275100 268072 275156
rect 331912 275100 336924 275156
rect 336980 275100 336990 275156
rect 262882 274540 262892 274596
rect 262948 274540 268072 274596
rect 331912 274540 334572 274596
rect 334628 274540 334638 274596
rect 263788 273980 268072 274036
rect 331912 273980 334460 274036
rect 334516 273980 334526 274036
rect 263788 273812 263844 273980
rect 256274 273756 256284 273812
rect 256340 273756 263844 273812
rect 261314 273420 261324 273476
rect 261380 273420 268072 273476
rect 331912 273420 334348 273476
rect 334404 273420 334414 273476
rect 262098 272860 262108 272916
rect 262164 272860 268072 272916
rect 331912 272860 351036 272916
rect 351092 272860 351102 272916
rect 263778 272300 263788 272356
rect 263844 272300 268072 272356
rect 331912 272300 334460 272356
rect 334516 272300 334526 272356
rect 263890 271740 263900 271796
rect 263956 271740 268072 271796
rect 331912 271740 338492 271796
rect 338548 271740 338558 271796
rect 595560 271460 597000 271656
rect 582082 271404 582092 271460
rect 582148 271432 597000 271460
rect 582148 271404 595672 271432
rect 464482 271292 464492 271348
rect 464548 271292 473004 271348
rect 473060 271292 473070 271348
rect 264674 271180 264684 271236
rect 264740 271180 268072 271236
rect 331912 271180 352044 271236
rect 352100 271180 352110 271236
rect 141026 271068 141036 271124
rect 141092 271068 144060 271124
rect 144116 271068 144126 271124
rect 201618 271068 201628 271124
rect 201684 271068 206136 271124
rect 265010 270620 265020 270676
rect 265076 270620 268072 270676
rect 331912 270620 352268 270676
rect 352324 270620 352334 270676
rect 18386 270396 18396 270452
rect 18452 270396 20076 270452
rect 20132 270396 20142 270452
rect 82450 270396 82460 270452
rect 82516 270396 82526 270452
rect 123928 270396 127596 270452
rect 127652 270396 127662 270452
rect 534258 270396 534268 270452
rect 534324 270396 538104 270452
rect 61880 269724 64204 269780
rect 64260 269724 64270 269780
rect 82460 269752 82516 270396
rect 264786 270060 264796 270116
rect 264852 270060 268072 270116
rect 331912 270060 334460 270116
rect 334516 270060 334526 270116
rect 123928 269724 130172 269780
rect 130228 269724 130238 269780
rect 414652 269556 414708 269752
rect 455896 269724 457212 269780
rect 457268 269724 457278 269780
rect 473666 269724 473676 269780
rect 473732 269724 476056 269780
rect 263778 269500 263788 269556
rect 263844 269500 268072 269556
rect 331912 269500 352156 269556
rect 352212 269500 352222 269556
rect 414642 269500 414652 269556
rect 414708 269500 414718 269556
rect 61880 269052 64092 269108
rect 64148 269052 64158 269108
rect 123928 269052 127484 269108
rect 127540 269052 127550 269108
rect 404002 269052 404012 269108
rect 404068 269052 414120 269108
rect 455896 269052 458892 269108
rect 458948 269052 458958 269108
rect 472098 269052 472108 269108
rect 472164 269052 476056 269108
rect 579880 269052 583212 269108
rect 583268 269052 583278 269108
rect 261426 268940 261436 268996
rect 261492 268940 268072 268996
rect 331912 268940 335692 268996
rect 335748 268940 335758 268996
rect 457762 268716 457772 268772
rect 457828 268716 458668 268772
rect 458724 268716 458734 268772
rect 18386 268380 18396 268436
rect 18452 268380 20104 268436
rect 141026 268380 141036 268436
rect 141092 268380 144088 268436
rect 185864 268380 189532 268436
rect 189588 268380 189598 268436
rect 20066 267708 20076 267764
rect 20132 267708 20142 267764
rect 61880 267708 64204 267764
rect 64260 267708 64270 267764
rect 185864 267708 205772 267764
rect 205828 267708 205838 267764
rect 206444 267652 206500 268408
rect 264898 268380 264908 268436
rect 264964 268380 268072 268436
rect 331912 268380 334348 268436
rect 334404 268380 334414 268436
rect 349346 268380 349356 268436
rect 349412 268380 352716 268436
rect 352772 268380 352782 268436
rect 410722 268380 410732 268436
rect 410788 268380 414120 268436
rect 455522 268380 455532 268436
rect 455588 268380 455598 268436
rect 472098 268380 472108 268436
rect 472164 268380 476056 268436
rect 534258 268380 534268 268436
rect 534324 268380 538104 268436
rect 248098 267932 248108 267988
rect 248164 267932 265132 267988
rect 265188 267932 265198 267988
rect 263778 267820 263788 267876
rect 263844 267820 268072 267876
rect 331912 267820 338716 267876
rect 338772 267820 338782 267876
rect 338482 267708 338492 267764
rect 338548 267708 352072 267764
rect 206434 267596 206444 267652
rect 206500 267596 206510 267652
rect 517468 267316 517524 267736
rect 579880 267708 583100 267764
rect 583156 267708 583166 267764
rect 248098 267260 248108 267316
rect 248164 267260 268072 267316
rect 331912 267260 334460 267316
rect 334516 267260 334526 267316
rect 517458 267260 517468 267316
rect 517524 267260 517534 267316
rect 203074 267036 203084 267092
rect 203140 267036 206136 267092
rect 247912 267036 262444 267092
rect 262500 267036 262510 267092
rect 345202 267036 345212 267092
rect 345268 267036 352072 267092
rect 393960 267036 395052 267092
rect 395108 267036 395118 267092
rect 579282 267036 579292 267092
rect 579348 267036 579358 267092
rect 82450 266924 82460 266980
rect 82516 266924 82526 266980
rect 82460 266392 82516 266924
rect 263778 266700 263788 266756
rect 263844 266700 268072 266756
rect 331912 266700 335244 266756
rect 335300 266700 335310 266756
rect 189522 266588 189532 266644
rect 189588 266588 199836 266644
rect 199892 266588 199902 266644
rect 123928 266364 130284 266420
rect 130340 266364 130350 266420
rect 142594 266364 142604 266420
rect 142660 266364 144088 266420
rect 185864 266364 189532 266420
rect 189588 266364 189598 266420
rect 204866 266364 204876 266420
rect 204932 266364 206136 266420
rect 247912 266364 259532 266420
rect 259588 266364 259598 266420
rect 407362 266364 407372 266420
rect 407428 266364 414120 266420
rect 472098 266364 472108 266420
rect 472164 266364 476056 266420
rect 579880 266364 583548 266420
rect 583604 266364 583614 266420
rect 335682 266252 335692 266308
rect 335748 266252 347788 266308
rect 347844 266252 347854 266308
rect 393362 266252 393372 266308
rect 393428 266252 393438 266308
rect 206322 266140 206332 266196
rect 206388 266140 206398 266196
rect 263778 266140 263788 266196
rect 263844 266140 268072 266196
rect 331912 266140 334460 266196
rect 334516 266140 334526 266196
rect 61880 265692 64652 265748
rect 64708 265692 64718 265748
rect 80434 265692 80444 265748
rect 80500 265692 82040 265748
rect 123928 265692 126812 265748
rect 126868 265692 126878 265748
rect 206332 265720 206388 266140
rect 247912 265692 262220 265748
rect 262276 265692 262286 265748
rect 336802 265692 336812 265748
rect 336868 265692 352072 265748
rect 393372 265720 393428 266252
rect 579852 266140 582092 266196
rect 582148 266140 582158 266196
rect 455896 265692 456988 265748
rect 457044 265692 457054 265748
rect 461122 265692 461132 265748
rect 461188 265692 476056 265748
rect 517794 265692 517804 265748
rect 517860 265692 517870 265748
rect 579852 265720 579908 266140
rect 260306 265580 260316 265636
rect 260372 265580 268072 265636
rect 331912 265580 335468 265636
rect 335524 265580 335534 265636
rect 61880 265020 69692 265076
rect 69748 265020 69758 265076
rect 127586 265020 127596 265076
rect 127652 265020 133532 265076
rect 133588 265020 133598 265076
rect 140914 265020 140924 265076
rect 140980 265020 144088 265076
rect 206098 265020 206108 265076
rect 206164 265020 206174 265076
rect 249554 265020 249564 265076
rect 249620 265020 268072 265076
rect 331912 265020 338604 265076
rect 338660 265020 338670 265076
rect 393960 265020 394940 265076
rect 394996 265020 395006 265076
rect 402322 265020 402332 265076
rect 402388 265020 414120 265076
rect 455896 265020 458668 265076
rect 458724 265020 458734 265076
rect 393362 264796 393372 264852
rect 393428 264796 393438 264852
rect 264002 264460 264012 264516
rect 264068 264460 268072 264516
rect 331912 264460 334460 264516
rect 334516 264460 334526 264516
rect 123928 264348 136892 264404
rect 136948 264348 136958 264404
rect 202962 264348 202972 264404
rect 203028 264348 206136 264404
rect 348562 264348 348572 264404
rect 348628 264348 352072 264404
rect 393372 264376 393428 264796
rect 464482 264572 464492 264628
rect 464548 264572 472108 264628
rect 472164 264572 472174 264628
rect 472994 264348 473004 264404
rect 473060 264348 476056 264404
rect 517944 264348 520940 264404
rect 520996 264348 521006 264404
rect 579282 264348 579292 264404
rect 579348 264348 579358 264404
rect 252914 263900 252924 263956
rect 252980 263900 268072 263956
rect 331912 263900 334460 263956
rect 334516 263900 334526 263956
rect 580402 263788 580412 263844
rect 580468 263788 580478 263844
rect 61880 263676 64204 263732
rect 64260 263676 64270 263732
rect 123928 263676 126812 263732
rect 126868 263676 126878 263732
rect 61880 263004 64204 263060
rect 64260 263004 64270 263060
rect 80322 263004 80332 263060
rect 80388 263004 82040 263060
rect 123928 263004 127596 263060
rect 127652 263004 127662 263060
rect 144284 262836 144340 263704
rect 185864 263676 189196 263732
rect 189252 263676 189262 263732
rect 393960 263676 396620 263732
rect 396676 263676 396686 263732
rect 472882 263676 472892 263732
rect 472948 263676 476056 263732
rect 262322 263340 262332 263396
rect 262388 263340 268072 263396
rect 331912 263340 335356 263396
rect 335412 263340 335422 263396
rect 579628 263284 579684 263704
rect 580412 263508 580468 263788
rect 579852 263452 580468 263508
rect 579618 263228 579628 263284
rect 579684 263228 579694 263284
rect 185864 263004 204092 263060
rect 204148 263004 204158 263060
rect 392 262808 4396 262836
rect -960 262780 4396 262808
rect 4452 262780 4462 262836
rect 144274 262780 144284 262836
rect 144340 262780 144350 262836
rect -960 262584 480 262780
rect 247884 262612 247940 263032
rect 393960 263004 394828 263060
rect 394884 263004 394894 263060
rect 534258 263004 534268 263060
rect 534324 263004 538104 263060
rect 579852 263032 579908 263452
rect 262098 262780 262108 262836
rect 262164 262780 268072 262836
rect 331912 262780 334460 262836
rect 334516 262780 334526 262836
rect 247884 262556 268100 262612
rect 82674 262332 82684 262388
rect 82740 262332 82750 262388
rect 185836 262164 185892 262360
rect 268044 262248 268100 262556
rect 393960 262332 396956 262388
rect 397012 262332 397022 262388
rect 331912 262220 340396 262276
rect 340452 262220 340462 262276
rect 476028 262164 476084 262360
rect 517944 262332 521052 262388
rect 521108 262332 521118 262388
rect 579880 262332 582988 262388
rect 583044 262332 583054 262388
rect 185836 262108 188244 262164
rect 188188 262052 188244 262108
rect 472108 262108 476084 262164
rect 472108 262052 472164 262108
rect 188188 261996 194908 262052
rect 194964 261996 194974 262052
rect 468626 261996 468636 262052
rect 468692 261996 472164 262052
rect 579852 261996 580524 262052
rect 580580 261996 580590 262052
rect 61880 261660 64764 261716
rect 64820 261660 64830 261716
rect 262210 261660 262220 261716
rect 262276 261660 268072 261716
rect 331912 261660 334460 261716
rect 334516 261660 334526 261716
rect 393960 261660 396844 261716
rect 396900 261660 396910 261716
rect 398962 261660 398972 261716
rect 399028 261660 414120 261716
rect 455896 261660 457100 261716
rect 457156 261660 457166 261716
rect 579852 261688 579908 261996
rect 206434 261548 206444 261604
rect 206500 261548 206510 261604
rect 64194 261212 64204 261268
rect 64260 261212 81452 261268
rect 81508 261212 81518 261268
rect 123928 260988 135212 261044
rect 135268 260988 135278 261044
rect 142706 260988 142716 261044
rect 142772 260988 144088 261044
rect 206444 261016 206500 261548
rect 393474 261436 393484 261492
rect 393540 261436 393550 261492
rect 262434 261100 262444 261156
rect 262500 261100 268072 261156
rect 247912 260988 262108 261044
rect 262164 260988 262174 261044
rect 331884 260708 331940 261128
rect 348786 260988 348796 261044
rect 348852 260988 352072 261044
rect 393484 261016 393540 261436
rect 455896 260988 458780 261044
rect 458836 260988 458846 261044
rect 472210 260988 472220 261044
rect 472276 260988 476056 261044
rect 579282 260988 579292 261044
rect 579348 260988 579358 261044
rect 331884 260652 334516 260708
rect 334460 260596 334516 260652
rect 261538 260540 261548 260596
rect 261604 260540 268072 260596
rect 331884 260484 331940 260568
rect 334450 260540 334460 260596
rect 334516 260540 334526 260596
rect 331884 260428 336924 260484
rect 336980 260428 336990 260484
rect 61880 260316 64652 260372
rect 64708 260316 64718 260372
rect 82002 260316 82012 260372
rect 82068 260316 82078 260372
rect 123928 260316 138572 260372
rect 138628 260316 138638 260372
rect 144050 260316 144060 260372
rect 144116 260316 144126 260372
rect 185864 260316 200732 260372
rect 200788 260316 200798 260372
rect 393250 260316 393260 260372
rect 393316 260316 393326 260372
rect 472098 260316 472108 260372
rect 472164 260316 476056 260372
rect 517944 260316 519148 260372
rect 519204 260316 519214 260372
rect 263778 259980 263788 260036
rect 263844 259980 268072 260036
rect 331912 259980 334460 260036
rect 334516 259980 334526 260036
rect 123928 259644 133532 259700
rect 133588 259644 133598 259700
rect 346882 259644 346892 259700
rect 346948 259644 352072 259700
rect 393960 259644 396620 259700
rect 396676 259644 396686 259700
rect 579880 259644 581308 259700
rect 581364 259644 581374 259700
rect 395602 259532 395612 259588
rect 395668 259532 395678 259588
rect 456866 259532 456876 259588
rect 456932 259532 472220 259588
rect 472276 259532 472286 259588
rect 395612 259476 395668 259532
rect 263890 259420 263900 259476
rect 263956 259420 268072 259476
rect 331912 259420 350476 259476
rect 350532 259420 350542 259476
rect 393932 259420 395668 259476
rect 185864 258972 188972 259028
rect 189028 258972 189038 259028
rect 247912 258972 262332 259028
rect 262388 258972 262398 259028
rect 393932 259000 393988 259420
rect 252914 258860 252924 258916
rect 252980 258860 268072 258916
rect 331912 258860 334460 258916
rect 334516 258860 334526 258916
rect 455868 258636 456092 258692
rect 456148 258636 456158 258692
rect 61880 258300 81564 258356
rect 81620 258300 81630 258356
rect 247912 258300 252812 258356
rect 252868 258300 252878 258356
rect 263778 258300 263788 258356
rect 263844 258300 268072 258356
rect 331912 258300 334460 258356
rect 334516 258300 334526 258356
rect 455868 258328 455924 258636
rect 517682 258300 517692 258356
rect 517748 258300 517758 258356
rect 535154 258300 535164 258356
rect 535220 258300 538104 258356
rect 595560 258216 597000 258440
rect 517458 258076 517468 258132
rect 517524 258076 517534 258132
rect 263890 257740 263900 257796
rect 263956 257740 268072 257796
rect 331912 257740 334348 257796
rect 334404 257740 334414 257796
rect 247912 257628 264012 257684
rect 264068 257628 264078 257684
rect 455298 257628 455308 257684
rect 455364 257628 455374 257684
rect 517468 257656 517524 258076
rect 259970 257180 259980 257236
rect 260036 257180 268072 257236
rect 331912 257180 335132 257236
rect 335188 257180 335198 257236
rect 262546 256620 262556 256676
rect 262612 256620 268072 256676
rect 331912 256620 351932 256676
rect 351988 256620 351998 256676
rect 247762 256060 247772 256116
rect 247828 256060 268072 256116
rect 331912 256060 351036 256116
rect 351092 256060 351102 256116
rect 265122 255500 265132 255556
rect 265188 255500 268072 255556
rect 331912 255500 334572 255556
rect 334628 255500 334638 255556
rect 258066 254940 258076 254996
rect 258132 254940 268072 254996
rect 331912 254940 334460 254996
rect 334516 254940 334526 254996
rect 262994 254380 263004 254436
rect 263060 254380 268072 254436
rect 331912 254380 334684 254436
rect 334740 254380 334750 254436
rect 263778 253820 263788 253876
rect 263844 253820 268072 253876
rect 331912 253820 334348 253876
rect 334404 253820 334414 253876
rect 263778 253260 263788 253316
rect 263844 253260 268072 253316
rect 331912 253260 350364 253316
rect 350420 253260 350430 253316
rect 64754 252812 64764 252868
rect 64820 252812 80556 252868
rect 80612 252812 80622 252868
rect 263890 252700 263900 252756
rect 263956 252700 268072 252756
rect 331912 252700 334460 252756
rect 334516 252700 334526 252756
rect 256162 252140 256172 252196
rect 256228 252140 268072 252196
rect 331912 252140 352156 252196
rect 352212 252140 352222 252196
rect 264562 251580 264572 251636
rect 264628 251580 268072 251636
rect 331912 251580 334460 251636
rect 334516 251580 334526 251636
rect 263778 251020 263788 251076
rect 263844 251020 268072 251076
rect 331912 251020 351036 251076
rect 351092 251020 351102 251076
rect 263778 250460 263788 250516
rect 263844 250460 268072 250516
rect 331912 250460 334348 250516
rect 334404 250460 334414 250516
rect 249442 249900 249452 249956
rect 249508 249900 268072 249956
rect 331912 249900 342076 249956
rect 342132 249900 342142 249956
rect 249778 249340 249788 249396
rect 249844 249340 268072 249396
rect 331912 249340 350252 249396
rect 350308 249340 350318 249396
rect 260306 248780 260316 248836
rect 260372 248780 268072 248836
rect 331912 248780 334460 248836
rect 334516 248780 334526 248836
rect -960 248472 480 248696
rect 252802 248220 252812 248276
rect 252868 248220 268072 248276
rect 331912 248220 334460 248276
rect 334516 248220 334526 248276
rect 253026 247660 253036 247716
rect 253092 247660 268072 247716
rect 331912 247660 351036 247716
rect 351092 247660 351102 247716
rect 263778 247100 263788 247156
rect 263844 247100 268072 247156
rect 331912 247100 338492 247156
rect 338548 247100 338558 247156
rect 248546 246540 248556 246596
rect 248612 246540 268072 246596
rect 331912 246540 346892 246596
rect 346948 246540 346958 246596
rect 336018 246204 336028 246260
rect 336084 246204 348572 246260
rect 348628 246204 348638 246260
rect 248434 246092 248444 246148
rect 248500 246092 263788 246148
rect 263844 246092 263854 246148
rect 335346 246092 335356 246148
rect 335412 246092 347788 246148
rect 347844 246092 347854 246148
rect 259522 245980 259532 246036
rect 259588 245980 268072 246036
rect 331912 245980 348796 246036
rect 348852 245980 348862 246036
rect 351026 245756 351036 245812
rect 351092 245756 410732 245812
rect 410788 245756 410798 245812
rect 255332 245420 268072 245476
rect 331912 245420 349468 245476
rect 349524 245420 349534 245476
rect 255332 245364 255388 245420
rect 18386 245308 18396 245364
rect 18452 245308 20972 245364
rect 21028 245308 21038 245364
rect 247996 245308 255388 245364
rect 247996 245252 248052 245308
rect 64642 245196 64652 245252
rect 64708 245196 248052 245252
rect 595560 245028 597000 245224
rect 333442 244972 333452 245028
rect 333508 245000 597000 245028
rect 333508 244972 595672 245000
rect 80546 244860 80556 244916
rect 80612 244860 268072 244916
rect 331912 244860 345212 244916
rect 345268 244860 345278 244916
rect 345986 244412 345996 244468
rect 346052 244412 396620 244468
rect 396676 244412 396686 244468
rect 81554 244300 81564 244356
rect 81620 244300 268072 244356
rect 331912 244300 336812 244356
rect 336868 244300 336878 244356
rect 261202 243740 261212 243796
rect 261268 243740 268072 243796
rect 331912 243740 336028 243796
rect 336084 243740 336094 243796
rect 338482 243292 338492 243348
rect 338548 243292 374892 243348
rect 374948 243292 374958 243348
rect 69682 243180 69692 243236
rect 69748 243180 268072 243236
rect 331912 243180 341852 243236
rect 341908 243180 341918 243236
rect 352146 243180 352156 243236
rect 352212 243180 438844 243236
rect 438900 243180 438910 243236
rect 222114 243068 222124 243124
rect 222180 243068 249564 243124
rect 249620 243068 249630 243124
rect 348562 243068 348572 243124
rect 348628 243068 436828 243124
rect 436884 243068 436894 243124
rect 108882 242956 108892 243012
rect 108948 242956 249788 243012
rect 249844 242956 249854 243012
rect 342178 242956 342188 243012
rect 342244 242956 448924 243012
rect 448980 242956 448990 243012
rect 94098 242844 94108 242900
rect 94164 242844 257964 242900
rect 258020 242844 258030 242900
rect 351922 242844 351932 242900
rect 351988 242844 493500 242900
rect 493556 242844 493566 242900
rect 167122 242732 167132 242788
rect 167188 242732 264684 242788
rect 264740 242732 264750 242788
rect 81442 242620 81452 242676
rect 81508 242620 268072 242676
rect 331912 242620 395052 242676
rect 395108 242620 395118 242676
rect 20962 242060 20972 242116
rect 21028 242060 268072 242116
rect 331912 242060 359548 242116
rect 359604 242060 359614 242116
rect 44258 241836 44268 241892
rect 44324 241836 261324 241892
rect 261380 241836 261390 241892
rect 349458 241836 349468 241892
rect 349524 241836 370188 241892
rect 370244 241836 370254 241892
rect 400642 241836 400652 241892
rect 400708 241836 562268 241892
rect 562324 241836 562334 241892
rect 38210 241724 38220 241780
rect 38276 241724 248556 241780
rect 248612 241724 248622 241780
rect 340274 241724 340284 241780
rect 340340 241724 494172 241780
rect 494228 241724 494238 241780
rect 106194 241612 106204 241668
rect 106260 241612 253036 241668
rect 253092 241612 253102 241668
rect 345202 241612 345212 241668
rect 345268 241612 432124 241668
rect 432180 241612 432190 241668
rect 192322 241500 192332 241556
rect 192388 241500 268072 241556
rect 331912 241500 394940 241556
rect 394996 241500 395006 241556
rect 166226 241388 166236 241444
rect 166292 241388 261548 241444
rect 261604 241388 261614 241444
rect 350354 241388 350364 241444
rect 350420 241388 434812 241444
rect 434868 241388 434878 241444
rect 352034 241276 352044 241332
rect 352100 241276 375564 241332
rect 375620 241276 375630 241332
rect 48626 241052 48636 241108
rect 48692 241052 264796 241108
rect 264852 241052 264862 241108
rect 20066 240940 20076 240996
rect 20132 240940 268072 240996
rect 331912 240940 345996 240996
rect 346052 240940 346062 240996
rect 263778 240380 263788 240436
rect 263844 240380 268072 240436
rect 331912 240380 503132 240436
rect 503188 240380 503198 240436
rect 26786 240156 26796 240212
rect 26852 240156 48636 240212
rect 48692 240156 48702 240212
rect 170258 240156 170268 240212
rect 170324 240156 187292 240212
rect 187348 240156 187358 240212
rect 222786 240156 222796 240212
rect 222852 240156 247884 240212
rect 247940 240156 247950 240212
rect 359538 240156 359548 240212
rect 359604 240156 372876 240212
rect 372932 240156 372942 240212
rect 37538 240044 37548 240100
rect 37604 240044 256284 240100
rect 256340 240044 256350 240100
rect 335458 240044 335468 240100
rect 335524 240044 555548 240100
rect 555604 240044 555614 240100
rect 46274 239932 46284 239988
rect 46340 239932 248444 239988
rect 248500 239932 248510 239988
rect 340386 239932 340396 239988
rect 340452 239932 560252 239988
rect 560308 239932 560318 239988
rect 42914 239820 42924 239876
rect 42980 239820 167132 239876
rect 167188 239820 167198 239876
rect 248546 239820 248556 239876
rect 248612 239820 268072 239876
rect 331912 239820 335916 239876
rect 335972 239820 335982 239876
rect 347778 239820 347788 239876
rect 347844 239820 553532 239876
rect 553588 239820 553598 239876
rect 163538 239708 163548 239764
rect 163604 239708 252924 239764
rect 252980 239708 252990 239764
rect 336914 239708 336924 239764
rect 336980 239708 496188 239764
rect 496244 239708 496254 239764
rect 162194 239596 162204 239652
rect 162260 239596 197372 239652
rect 197428 239596 197438 239652
rect 230850 239596 230860 239652
rect 230916 239596 257852 239652
rect 257908 239596 257918 239652
rect 335234 239596 335244 239652
rect 335300 239596 557564 239652
rect 557620 239596 557630 239652
rect 40226 239484 40236 239540
rect 40292 239484 262892 239540
rect 262948 239484 262958 239540
rect 249442 239372 249452 239428
rect 249508 239372 263788 239428
rect 263844 239372 263854 239428
rect 165554 239260 165564 239316
rect 165620 239260 249676 239316
rect 249732 239260 249742 239316
rect 263778 239260 263788 239316
rect 263844 239260 268072 239316
rect 331912 239260 334348 239316
rect 334404 239260 334414 239316
rect 263890 238700 263900 238756
rect 263956 238700 268072 238756
rect 331912 238700 335692 238756
rect 335748 238700 335758 238756
rect 262882 238140 262892 238196
rect 262948 238140 268072 238196
rect 331912 238140 334460 238196
rect 334516 238140 334526 238196
rect 261202 237580 261212 237636
rect 261268 237580 268072 237636
rect 331912 237580 338492 237636
rect 338548 237580 338558 237636
rect 259522 237020 259532 237076
rect 259588 237020 268072 237076
rect 331912 237020 335132 237076
rect 335188 237020 335198 237076
rect 203186 236460 203196 236516
rect 203252 236460 268072 236516
rect 331912 236460 400652 236516
rect 400708 236460 400718 236516
rect 204866 236012 204876 236068
rect 204932 236012 263788 236068
rect 263844 236012 263854 236068
rect 334450 236012 334460 236068
rect 334516 236012 536732 236068
rect 536788 236012 536798 236068
rect 264898 235900 264908 235956
rect 264964 235900 268072 235956
rect 331912 235900 560364 235956
rect 560420 235900 560430 235956
rect 257842 235340 257852 235396
rect 257908 235340 263900 235396
rect 263956 235340 263966 235396
rect 268044 235284 268100 235368
rect 331912 235340 581308 235396
rect 581364 235340 581374 235396
rect 263788 235228 268100 235284
rect 263788 235172 263844 235228
rect 262882 235116 262892 235172
rect 262948 235116 263844 235172
rect 261202 234780 261212 234836
rect 261268 234780 268072 234836
rect 331912 234780 523292 234836
rect 523348 234780 523358 234836
rect -960 234388 480 234584
rect 203074 234556 203084 234612
rect 203140 234556 248556 234612
rect 248612 234556 248622 234612
rect 4386 234444 4396 234500
rect 4452 234444 266476 234500
rect 266532 234444 266542 234500
rect -960 234360 264572 234388
rect 392 234332 264572 234360
rect 264628 234332 264638 234388
rect 256162 234220 256172 234276
rect 256228 234220 268072 234276
rect 331912 234220 459452 234276
rect 459508 234220 459518 234276
rect 263788 233660 268072 233716
rect 331912 233660 583436 233716
rect 583492 233660 583502 233716
rect 263788 233492 263844 233660
rect 257954 233436 257964 233492
rect 258020 233436 263844 233492
rect 225474 233100 225484 233156
rect 225540 233100 268072 233156
rect 331912 233100 350252 233156
rect 350308 233100 350318 233156
rect 334338 232652 334348 232708
rect 334404 232652 533484 232708
rect 533540 232652 533550 232708
rect 140578 232540 140588 232596
rect 140644 232540 268072 232596
rect 331912 232540 437612 232596
rect 437668 232540 437678 232596
rect 199042 231980 199052 232036
rect 199108 231980 268072 232036
rect 331912 231980 462812 232036
rect 462868 231980 462878 232036
rect 595560 231924 597000 232008
rect 336802 231868 336812 231924
rect 336868 231868 597000 231924
rect 595560 231784 597000 231868
rect 140690 231420 140700 231476
rect 140756 231420 268072 231476
rect 331912 231420 518364 231476
rect 518420 231420 518430 231476
rect 335906 230972 335916 231028
rect 335972 230972 583100 231028
rect 583156 230972 583166 231028
rect 195682 230860 195692 230916
rect 195748 230860 268072 230916
rect 331912 230860 473116 230916
rect 473172 230860 473182 230916
rect 140802 230300 140812 230356
rect 140868 230300 268072 230356
rect 331912 230300 440972 230356
rect 441028 230300 441038 230356
rect 140914 229740 140924 229796
rect 140980 229740 268072 229796
rect 331912 229740 519932 229796
rect 519988 229740 519998 229796
rect 166226 229180 166236 229236
rect 166292 229180 268072 229236
rect 331912 229180 418348 229236
rect 418404 229180 418414 229236
rect 163538 228620 163548 228676
rect 163604 228620 268072 228676
rect 331912 228620 520156 228676
rect 520212 228620 520222 228676
rect 189186 228060 189196 228116
rect 189252 228060 268072 228116
rect 331912 228060 396172 228116
rect 396228 228060 396238 228116
rect 338482 227612 338492 227668
rect 338548 227612 560252 227668
rect 560308 227612 560318 227668
rect 188962 227500 188972 227556
rect 189028 227500 268072 227556
rect 331912 227500 474684 227556
rect 474740 227500 474750 227556
rect 158834 226940 158844 226996
rect 158900 226940 268072 226996
rect 331912 226940 518252 226996
rect 518308 226940 518318 226996
rect 197362 226380 197372 226436
rect 197428 226380 268072 226436
rect 331912 226380 464492 226436
rect 464548 226380 464558 226436
rect 263890 225820 263900 225876
rect 263956 225820 268072 225876
rect 331912 225820 461132 225876
rect 461188 225820 461198 225876
rect 263778 225260 263788 225316
rect 263844 225260 268072 225316
rect 331912 225260 338492 225316
rect 338548 225260 338558 225316
rect 80322 224700 80332 224756
rect 80388 224700 268072 224756
rect 331912 224700 427532 224756
rect 427588 224700 427598 224756
rect 418338 224364 418348 224420
rect 418404 224364 520940 224420
rect 520996 224364 521006 224420
rect 144050 224252 144060 224308
rect 144116 224252 263788 224308
rect 263844 224252 263854 224308
rect 335122 224252 335132 224308
rect 335188 224252 581420 224308
rect 581476 224252 581486 224308
rect 133522 224140 133532 224196
rect 133588 224140 268072 224196
rect 331912 224140 414092 224196
rect 414148 224140 414158 224196
rect 126802 223580 126812 223636
rect 126868 223580 268072 223636
rect 331912 223580 419132 223636
rect 419188 223580 419198 223636
rect 80098 223020 80108 223076
rect 80164 223020 268072 223076
rect 331912 223020 406588 223076
rect 406644 223020 406654 223076
rect 192322 222572 192332 222628
rect 192388 222572 263900 222628
rect 263956 222572 263966 222628
rect 350242 222572 350252 222628
rect 350308 222572 564284 222628
rect 564340 222572 564350 222628
rect 80434 222460 80444 222516
rect 80500 222460 268072 222516
rect 331912 222460 455308 222516
rect 455364 222460 455374 222516
rect 126914 221900 126924 221956
rect 126980 221900 268072 221956
rect 331912 221900 429212 221956
rect 429268 221900 429278 221956
rect 83122 221340 83132 221396
rect 83188 221340 268072 221396
rect 331912 221340 351932 221396
rect 351988 221340 351998 221396
rect 130162 220780 130172 220836
rect 130228 220780 268072 220836
rect 331912 220780 335916 220836
rect 335972 220780 335982 220836
rect 392 220472 4284 220500
rect -960 220444 4284 220472
rect 4340 220444 4350 220500
rect -960 220248 480 220444
rect 263778 220220 263788 220276
rect 263844 220220 268072 220276
rect 331912 220220 398972 220276
rect 399028 220220 399038 220276
rect 105522 219660 105532 219716
rect 105588 219660 268072 219716
rect 331912 219660 407372 219716
rect 407428 219660 407438 219716
rect 406578 219324 406588 219380
rect 406644 219324 434140 219380
rect 434196 219324 434206 219380
rect 82002 219212 82012 219268
rect 82068 219212 263788 219268
rect 263844 219212 263854 219268
rect 335682 219212 335692 219268
rect 335748 219212 579628 219268
rect 579684 219212 579694 219268
rect 102162 219100 102172 219156
rect 102228 219100 268072 219156
rect 331912 219100 339276 219156
rect 339332 219100 339342 219156
rect 263778 218540 263788 218596
rect 263844 218540 268072 218596
rect 331912 218540 412412 218596
rect 412468 218540 412478 218596
rect 595560 218568 597000 218792
rect 427522 218092 427532 218148
rect 427588 218092 433468 218148
rect 433524 218092 433534 218148
rect 106194 217980 106204 218036
rect 106260 217980 268072 218036
rect 331912 217980 356188 218036
rect 356244 217980 356254 218036
rect 429202 217756 429212 217812
rect 429268 217756 439516 217812
rect 439572 217756 439582 217812
rect 440962 217756 440972 217812
rect 441028 217756 501564 217812
rect 501620 217756 501630 217812
rect 437602 217644 437612 217700
rect 437668 217644 500892 217700
rect 500948 217644 500958 217700
rect 82226 217532 82236 217588
rect 82292 217532 263788 217588
rect 263844 217532 263854 217588
rect 335906 217532 335916 217588
rect 335972 217532 456988 217588
rect 457044 217532 457054 217588
rect 503122 217532 503132 217588
rect 503188 217532 555548 217588
rect 555604 217532 555614 217588
rect 104178 217420 104188 217476
rect 104244 217420 268072 217476
rect 331912 217420 436156 217476
rect 436212 217420 436222 217476
rect 141922 216860 141932 216916
rect 141988 216860 268072 216916
rect 331912 216860 372876 216916
rect 372932 216860 372942 216916
rect 560354 216636 560364 216692
rect 560420 216636 562268 216692
rect 562324 216636 562334 216692
rect 263778 216300 263788 216356
rect 263844 216300 268072 216356
rect 331912 216300 336028 216356
rect 336084 216300 336094 216356
rect 41570 215964 41580 216020
rect 41636 215964 256284 216020
rect 256340 215964 256350 216020
rect 101490 215852 101500 215908
rect 101556 215852 228508 215908
rect 228564 215852 228574 215908
rect 252802 215852 252812 215908
rect 252868 215852 264908 215908
rect 264964 215852 264974 215908
rect 222786 215740 222796 215796
rect 222852 215740 249676 215796
rect 249732 215740 249742 215796
rect 263890 215740 263900 215796
rect 263956 215740 268072 215796
rect 331912 215740 336812 215796
rect 336868 215740 336878 215796
rect 164210 215628 164220 215684
rect 164276 215628 253036 215684
rect 253092 215628 253102 215684
rect 335234 215628 335244 215684
rect 335300 215628 562940 215684
rect 562996 215628 563006 215684
rect 223458 215516 223468 215572
rect 223524 215516 256508 215572
rect 256564 215516 256574 215572
rect 338482 215516 338492 215572
rect 338548 215516 437500 215572
rect 437556 215516 437566 215572
rect 475458 215516 475468 215572
rect 475524 215516 496860 215572
rect 496916 215516 496926 215572
rect 40898 215404 40908 215460
rect 40964 215404 61292 215460
rect 61348 215404 61358 215460
rect 106866 215404 106876 215460
rect 106932 215404 259756 215460
rect 259812 215404 259822 215460
rect 352146 215404 352156 215460
rect 352212 215404 495516 215460
rect 495572 215404 495582 215460
rect 35522 215292 35532 215348
rect 35588 215292 83804 215348
rect 83860 215292 83870 215348
rect 103506 215292 103516 215348
rect 103572 215292 258188 215348
rect 258244 215292 258254 215348
rect 348562 215292 348572 215348
rect 348628 215292 492156 215348
rect 492212 215292 492222 215348
rect 539186 215292 539196 215348
rect 539252 215292 558908 215348
rect 558964 215292 558974 215348
rect 98130 215180 98140 215236
rect 98196 215180 261548 215236
rect 261604 215180 261614 215236
rect 264674 215180 264684 215236
rect 264740 215180 268072 215236
rect 331912 215180 337036 215236
rect 337092 215180 337102 215236
rect 340274 215180 340284 215236
rect 340340 215180 563612 215236
rect 563668 215180 563678 215236
rect 44930 215068 44940 215124
rect 44996 215068 99484 215124
rect 99540 215068 99550 215124
rect 159506 215068 159516 215124
rect 159572 215068 186396 215124
rect 186452 215068 186462 215124
rect 228834 215068 228844 215124
rect 228900 215068 247996 215124
rect 248052 215068 248062 215124
rect 350354 215068 350364 215124
rect 350420 215068 368172 215124
rect 368228 215068 368238 215124
rect 74722 214620 74732 214676
rect 74788 214620 268072 214676
rect 331912 214620 340396 214676
rect 340452 214620 340462 214676
rect 356178 214396 356188 214452
rect 356244 214396 410732 214452
rect 410788 214396 410798 214452
rect 228498 214284 228508 214340
rect 228564 214284 264908 214340
rect 264964 214284 264974 214340
rect 336018 214284 336028 214340
rect 336084 214284 396732 214340
rect 396788 214284 396798 214340
rect 419122 214284 419132 214340
rect 419188 214284 458892 214340
rect 458948 214284 458958 214340
rect 459442 214284 459452 214340
rect 459508 214284 535276 214340
rect 535332 214284 535342 214340
rect 81442 214172 81452 214228
rect 81508 214172 263788 214228
rect 263844 214172 263854 214228
rect 338482 214172 338492 214228
rect 338548 214172 472108 214228
rect 472164 214172 472174 214228
rect 206658 214060 206668 214116
rect 206724 214060 268072 214116
rect 331912 214060 340620 214116
rect 340676 214060 340686 214116
rect 166898 213836 166908 213892
rect 166964 213836 254492 213892
rect 254548 213836 254558 213892
rect 98802 213724 98812 213780
rect 98868 213724 249788 213780
rect 249844 213724 249854 213780
rect 351922 213724 351932 213780
rect 351988 213724 376236 213780
rect 376292 213724 376302 213780
rect 46946 213612 46956 213668
rect 47012 213612 248556 213668
rect 248612 213612 248622 213668
rect 339266 213612 339276 213668
rect 339332 213612 366716 213668
rect 366772 213612 366782 213668
rect 45602 213500 45612 213556
rect 45668 213500 249564 213556
rect 249620 213500 249630 213556
rect 263778 213500 263788 213556
rect 263844 213500 268072 213556
rect 331912 213500 340172 213556
rect 340228 213500 340238 213556
rect 345538 213500 345548 213556
rect 345604 213500 430780 213556
rect 430836 213500 430846 213556
rect 40226 213388 40236 213444
rect 40292 213388 263116 213444
rect 263172 213388 263182 213444
rect 350466 213388 350476 213444
rect 350532 213388 496188 213444
rect 496244 213388 496254 213444
rect 73042 213276 73052 213332
rect 73108 213276 263900 213332
rect 263956 213276 263966 213332
rect 352034 213276 352044 213332
rect 352100 213276 436828 213332
rect 436884 213276 436894 213332
rect 99474 213164 99484 213220
rect 99540 213164 261100 213220
rect 261156 213164 261166 213220
rect 339266 213164 339276 213220
rect 339332 213164 458780 213220
rect 458836 213164 458846 213220
rect 69682 213052 69692 213108
rect 69748 213052 268100 213108
rect 44258 212940 44268 212996
rect 44324 212940 261436 212996
rect 261492 212940 261502 212996
rect 268044 212968 268100 213052
rect 337652 213052 395836 213108
rect 395892 213052 395902 213108
rect 396162 213052 396172 213108
rect 396228 213052 521164 213108
rect 521220 213052 521230 213108
rect 331884 212884 331940 212968
rect 102834 212828 102844 212884
rect 102900 212828 114268 212884
rect 160150 212828 160188 212884
rect 160244 212828 160254 212884
rect 226818 212828 226828 212884
rect 226884 212828 226894 212884
rect 231494 212828 231532 212884
rect 231588 212828 231598 212884
rect 331884 212828 334460 212884
rect 334516 212828 334526 212884
rect 114212 212660 114268 212828
rect 226828 212772 226884 212828
rect 337652 212772 337708 213052
rect 342066 212940 342076 212996
rect 342132 212940 557564 212996
rect 557620 212940 557630 212996
rect 370822 212828 370860 212884
rect 370916 212828 370926 212884
rect 375778 212828 375788 212884
rect 375844 212828 378252 212884
rect 378308 212828 378318 212884
rect 156212 212716 168028 212772
rect 226828 212716 231756 212772
rect 231812 212716 231822 212772
rect 331996 212716 337708 212772
rect 372988 212716 384748 212772
rect 156212 212660 156268 212716
rect 167972 212660 168028 212716
rect 114212 212604 156268 212660
rect 160178 212604 160188 212660
rect 160244 212604 160254 212660
rect 167972 212604 252812 212660
rect 252868 212604 252878 212660
rect 160188 212548 160244 212604
rect 331996 212548 332052 212716
rect 372988 212660 373044 212716
rect 384692 212660 384748 212716
rect 334450 212604 334460 212660
rect 334516 212604 373044 212660
rect 375778 212604 375788 212660
rect 375844 212604 375854 212660
rect 384692 212604 396620 212660
rect 396676 212604 396686 212660
rect 375788 212548 375844 212604
rect 160188 212492 247884 212548
rect 247940 212492 247950 212548
rect 331884 212492 332052 212548
rect 350242 212492 350252 212548
rect 350308 212492 375844 212548
rect 231522 212380 231532 212436
rect 231588 212380 231598 212436
rect 231746 212380 231756 212436
rect 231812 212380 248108 212436
rect 248164 212380 248174 212436
rect 259634 212380 259644 212436
rect 259700 212380 268072 212436
rect 331884 212408 331940 212492
rect 341842 212380 341852 212436
rect 341908 212380 370860 212436
rect 370916 212380 370926 212436
rect 231532 212324 231588 212380
rect 231532 212268 249900 212324
rect 249956 212268 249966 212324
rect 261090 212156 261100 212212
rect 261156 212156 268100 212212
rect 74834 212044 74844 212100
rect 74900 212044 263788 212100
rect 263844 212044 263854 212100
rect 268044 211848 268100 212156
rect 331912 211820 338492 211876
rect 338548 211820 338558 211876
rect 79986 211596 79996 211652
rect 80052 211596 83132 211652
rect 83188 211596 83198 211652
rect 125122 211260 125132 211316
rect 125188 211260 268072 211316
rect 331912 211260 396396 211316
rect 396452 211260 396462 211316
rect 80210 211148 80220 211204
rect 80276 211148 130172 211204
rect 130228 211148 130238 211204
rect 186386 211148 186396 211204
rect 186452 211148 263788 211204
rect 263844 211148 263854 211204
rect 351922 211148 351932 211204
rect 351988 211148 410844 211204
rect 410900 211148 410910 211204
rect 462802 211148 462812 211204
rect 462868 211148 521052 211204
rect 521108 211148 521118 211204
rect 64642 211036 64652 211092
rect 64708 211036 206668 211092
rect 206724 211036 206734 211092
rect 335346 211036 335356 211092
rect 335412 211036 475468 211092
rect 475524 211036 475534 211092
rect 83794 210924 83804 210980
rect 83860 210924 265020 210980
rect 265076 210924 265086 210980
rect 400642 210924 400652 210980
rect 400708 210924 583324 210980
rect 583380 210924 583390 210980
rect 61282 210812 61292 210868
rect 61348 210812 264796 210868
rect 264852 210812 264862 210868
rect 335906 210812 335916 210868
rect 335972 210812 539196 210868
rect 539252 210812 539262 210868
rect 81666 210700 81676 210756
rect 81732 210700 268072 210756
rect 331912 210700 396844 210756
rect 396900 210700 396910 210756
rect 351138 210588 351148 210644
rect 351204 210588 535164 210644
rect 535220 210588 535230 210644
rect 345986 210476 345996 210532
rect 346052 210476 535500 210532
rect 535556 210476 535566 210532
rect 20066 210364 20076 210420
rect 20132 210364 263788 210420
rect 263844 210364 263854 210420
rect 351026 210364 351036 210420
rect 351092 210364 583212 210420
rect 583268 210364 583278 210420
rect 248546 210140 248556 210196
rect 248612 210140 268072 210196
rect 331912 210140 340284 210196
rect 340340 210140 340350 210196
rect 263778 209580 263788 209636
rect 263844 209580 268072 209636
rect 331912 209580 339276 209636
rect 339332 209580 339342 209636
rect 251906 209020 251916 209076
rect 251972 209020 268072 209076
rect 331912 209020 351036 209076
rect 351092 209020 351102 209076
rect 144050 208572 144060 208628
rect 144116 208572 144126 208628
rect 472098 208572 472108 208628
rect 472164 208572 476056 208628
rect 252914 208460 252924 208516
rect 252980 208460 268072 208516
rect 331912 208460 335132 208516
rect 335188 208460 335198 208516
rect 247762 207900 247772 207956
rect 247828 207900 268072 207956
rect 331912 207900 351148 207956
rect 351204 207900 351214 207956
rect 247986 207340 247996 207396
rect 248052 207340 268072 207396
rect 331912 207340 335244 207396
rect 335300 207340 335310 207396
rect 262098 206780 262108 206836
rect 262164 206780 268072 206836
rect 331912 206780 340284 206836
rect 340340 206780 340350 206836
rect -960 206136 480 206360
rect 258066 206220 258076 206276
rect 258132 206220 268072 206276
rect 331912 206220 334460 206276
rect 334516 206220 334526 206276
rect 247912 205884 261212 205940
rect 261268 205884 261278 205940
rect 264786 205660 264796 205716
rect 264852 205660 268072 205716
rect 331912 205660 335916 205716
rect 335972 205660 335982 205716
rect 595560 205352 597000 205576
rect 264562 205100 264572 205156
rect 264628 205100 268072 205156
rect 331912 205100 340284 205156
rect 340340 205100 340350 205156
rect 256498 204540 256508 204596
rect 256564 204540 268072 204596
rect 331912 204540 334460 204596
rect 334516 204540 334526 204596
rect 248098 203980 248108 204036
rect 248164 203980 268072 204036
rect 331912 203980 342076 204036
rect 342132 203980 342142 204036
rect 249890 203420 249900 203476
rect 249956 203420 268072 203476
rect 331912 203420 345996 203476
rect 346052 203420 346062 203476
rect 249666 202860 249676 202916
rect 249732 202860 268072 202916
rect 331912 202860 335244 202916
rect 335300 202860 335310 202916
rect 256162 202300 256172 202356
rect 256228 202300 268072 202356
rect 331912 202300 334460 202356
rect 334516 202300 334526 202356
rect 262994 201740 263004 201796
rect 263060 201740 268072 201796
rect 331912 201740 341852 201796
rect 341908 201740 341918 201796
rect 254482 201180 254492 201236
rect 254548 201180 268072 201236
rect 331912 201180 352156 201236
rect 352212 201180 352222 201236
rect 263778 200620 263788 200676
rect 263844 200620 268072 200676
rect 331912 200620 334460 200676
rect 334516 200620 334526 200676
rect 247874 200060 247884 200116
rect 247940 200060 268072 200116
rect 331912 200060 348572 200116
rect 348628 200060 348638 200116
rect 141026 199836 141036 199892
rect 141092 199836 144088 199892
rect 201618 199836 201628 199892
rect 201684 199836 206136 199892
rect 253026 199500 253036 199556
rect 253092 199500 268072 199556
rect 331912 199500 345212 199556
rect 345268 199500 345278 199556
rect 393960 199164 396508 199220
rect 396564 199164 396574 199220
rect 414652 199108 414708 199864
rect 534258 199164 534268 199220
rect 534324 199164 538104 199220
rect 414642 199052 414652 199108
rect 414708 199052 414718 199108
rect 18358 198940 18396 198996
rect 18452 198940 18462 198996
rect 263778 198940 263788 198996
rect 263844 198940 268072 198996
rect 331912 198940 334460 198996
rect 334516 198940 334526 198996
rect 82674 198492 82684 198548
rect 82740 198492 82750 198548
rect 140690 198492 140700 198548
rect 140756 198492 144088 198548
rect 349346 198492 349356 198548
rect 349412 198492 352716 198548
rect 352772 198492 352782 198548
rect 455298 198492 455308 198548
rect 455364 198492 455374 198548
rect 261314 198380 261324 198436
rect 261380 198380 268072 198436
rect 331912 198380 335356 198436
rect 335412 198380 335422 198436
rect 18386 197820 18396 197876
rect 18452 197820 20104 197876
rect 80322 197820 80332 197876
rect 80388 197820 82040 197876
rect 263890 197820 263900 197876
rect 263956 197820 268072 197876
rect 331912 197820 334348 197876
rect 334404 197820 334414 197876
rect 473666 197820 473676 197876
rect 473732 197820 476056 197876
rect 263778 197260 263788 197316
rect 263844 197260 268072 197316
rect 331912 197260 334460 197316
rect 334516 197260 334526 197316
rect 61880 197148 64204 197204
rect 64260 197148 64270 197204
rect 185864 197148 197372 197204
rect 197428 197148 197438 197204
rect 579618 197148 579628 197204
rect 579684 197148 579694 197204
rect 248546 196700 248556 196756
rect 248612 196700 268072 196756
rect 331912 196700 350476 196756
rect 350532 196700 350542 196756
rect 455308 196700 455420 196756
rect 455476 196700 455486 196756
rect 395826 196588 395836 196644
rect 395892 196588 396508 196644
rect 396564 196588 396574 196644
rect 20636 196084 20692 196504
rect 185864 196476 196588 196532
rect 196644 196476 196654 196532
rect 337026 196476 337036 196532
rect 337092 196476 352072 196532
rect 393960 196476 394828 196532
rect 394884 196476 394894 196532
rect 410834 196476 410844 196532
rect 410900 196476 414120 196532
rect 455308 196504 455364 196700
rect 467842 196476 467852 196532
rect 467908 196476 476056 196532
rect 517944 196476 520940 196532
rect 520996 196476 521006 196532
rect 524962 196476 524972 196532
rect 525028 196476 538104 196532
rect 579880 196476 583324 196532
rect 583380 196476 583390 196532
rect 520146 196364 520156 196420
rect 520212 196364 520222 196420
rect 520156 196308 520212 196364
rect 517916 196252 520212 196308
rect 263778 196140 263788 196196
rect 263844 196140 268072 196196
rect 331912 196140 334460 196196
rect 334516 196140 334526 196196
rect 20626 196028 20636 196084
rect 20692 196028 20702 196084
rect 20300 194964 20356 195832
rect 185864 195804 189532 195860
rect 189588 195804 189598 195860
rect 340610 195804 340620 195860
rect 340676 195804 352072 195860
rect 517916 195832 517972 196252
rect 535490 195804 535500 195860
rect 535556 195804 538104 195860
rect 579880 195804 581420 195860
rect 581476 195804 581486 195860
rect 261538 195580 261548 195636
rect 261604 195580 268072 195636
rect 331912 195580 338492 195636
rect 338548 195580 338558 195636
rect 331884 195356 351932 195412
rect 351988 195356 351998 195412
rect 61880 195132 64204 195188
rect 64260 195132 64270 195188
rect 80434 195132 80444 195188
rect 80500 195132 82040 195188
rect 123928 195132 127484 195188
rect 127540 195132 127550 195188
rect 185864 195132 189196 195188
rect 189252 195132 189262 195188
rect 202962 195132 202972 195188
rect 203028 195132 206136 195188
rect 247912 195132 262892 195188
rect 262948 195132 262958 195188
rect 249778 195020 249788 195076
rect 249844 195020 268072 195076
rect 331884 195048 331940 195356
rect 340386 195132 340396 195188
rect 340452 195132 352072 195188
rect 393960 195132 396732 195188
rect 396788 195132 396798 195188
rect 411170 195132 411180 195188
rect 411236 195132 414120 195188
rect 535266 195132 535276 195188
rect 535332 195132 538104 195188
rect 20290 194908 20300 194964
rect 20356 194908 20366 194964
rect 61740 194684 67228 194740
rect 20066 194460 20076 194516
rect 20132 194460 20142 194516
rect 61740 194488 61796 194684
rect 67172 194628 67228 194684
rect 67172 194572 81676 194628
rect 81732 194572 81742 194628
rect 79986 194460 79996 194516
rect 80052 194460 82040 194516
rect 123928 194460 127596 194516
rect 127652 194460 127662 194516
rect 247912 194460 257964 194516
rect 258020 194460 258030 194516
rect 258178 194460 258188 194516
rect 258244 194460 268072 194516
rect 331912 194460 334460 194516
rect 334516 194460 334526 194516
rect 340162 194460 340172 194516
rect 340228 194460 352072 194516
rect 411282 194460 411292 194516
rect 411348 194460 414120 194516
rect 455308 194068 455364 194488
rect 61740 194012 67228 194068
rect 455298 194012 455308 194068
rect 455364 194012 455374 194068
rect 61740 193816 61796 194012
rect 67172 193956 67228 194012
rect 67172 193900 81452 193956
rect 81508 193900 81518 193956
rect 252802 193900 252812 193956
rect 252868 193900 268072 193956
rect 331912 193900 334348 193956
rect 334404 193900 334414 193956
rect 80210 193788 80220 193844
rect 80276 193788 82040 193844
rect 185864 193788 192332 193844
rect 192388 193788 192398 193844
rect 247912 193788 264796 193844
rect 264852 193788 264862 193844
rect 455896 193788 456988 193844
rect 457044 193788 457054 193844
rect 472098 193788 472108 193844
rect 472164 193788 476056 193844
rect 264002 193340 264012 193396
rect 264068 193340 268072 193396
rect 331912 193340 334460 193396
rect 334516 193340 334526 193396
rect 519922 193228 519932 193284
rect 519988 193228 519998 193284
rect 519932 193172 519988 193228
rect 185864 193116 188972 193172
rect 189028 193116 189038 193172
rect 393960 193116 396508 193172
rect 396564 193116 396574 193172
rect 517944 193116 519988 193172
rect 535154 193116 535164 193172
rect 535220 193116 538104 193172
rect 579880 193116 583100 193172
rect 583156 193116 583166 193172
rect 264898 192780 264908 192836
rect 264964 192780 268072 192836
rect 331912 192780 345324 192836
rect 345380 192780 345390 192836
rect 334338 192668 334348 192724
rect 334404 192668 351820 192724
rect 351876 192668 351886 192724
rect 61880 192444 74844 192500
rect 74900 192444 74910 192500
rect 123928 192444 126924 192500
rect 126980 192444 126990 192500
rect 140802 192444 140812 192500
rect 140868 192444 144088 192500
rect 340274 192444 340284 192500
rect 340340 192444 352072 192500
rect 411170 192444 411180 192500
rect 411236 192444 414120 192500
rect 517944 192444 521052 192500
rect 521108 192444 521118 192500
rect 189522 192332 189532 192388
rect 189588 192332 204988 192388
rect 205044 192332 205054 192388
rect 463586 192332 463596 192388
rect 463652 192332 472108 192388
rect 472164 192332 472174 192388
rect -960 192052 480 192248
rect 249666 192220 249676 192276
rect 249732 192220 268072 192276
rect 331912 192220 334460 192276
rect 334516 192220 334526 192276
rect 595560 192164 597000 192360
rect 580402 192108 580412 192164
rect 580468 192136 597000 192164
rect 580468 192108 595672 192136
rect -960 192024 4620 192052
rect 392 191996 4620 192024
rect 4676 191996 4686 192052
rect 185864 191772 205660 191828
rect 205716 191772 205726 191828
rect 247912 191772 256172 191828
rect 256228 191772 256238 191828
rect 393960 191772 396732 191828
rect 396788 191772 396798 191828
rect 410722 191772 410732 191828
rect 410788 191772 414120 191828
rect 455896 191772 458892 191828
rect 458948 191772 458958 191828
rect 263778 191660 263788 191716
rect 263844 191660 268072 191716
rect 331912 191660 345548 191716
rect 345604 191660 345614 191716
rect 518354 191436 518364 191492
rect 518420 191436 518430 191492
rect 247772 191324 255388 191380
rect 123928 191100 127596 191156
rect 127652 191100 127662 191156
rect 247772 191128 247828 191324
rect 255332 191268 255388 191324
rect 255332 191212 264572 191268
rect 264628 191212 264638 191268
rect 518364 191156 518420 191436
rect 258402 191100 258412 191156
rect 258468 191100 268072 191156
rect 331884 191044 331940 191128
rect 338482 191100 338492 191156
rect 338548 191100 352072 191156
rect 407362 191100 407372 191156
rect 407428 191100 414120 191156
rect 455896 191100 458780 191156
rect 458836 191100 458846 191156
rect 472098 191100 472108 191156
rect 472164 191100 476056 191156
rect 517916 191100 518420 191156
rect 331884 190988 341964 191044
rect 342020 190988 342030 191044
rect 259746 190540 259756 190596
rect 259812 190540 268072 190596
rect 331912 190540 334348 190596
rect 334404 190540 334414 190596
rect 80098 190428 80108 190484
rect 80164 190428 82040 190484
rect 247912 190428 252812 190484
rect 252868 190428 252878 190484
rect 517916 190456 517972 191100
rect 579730 190988 579740 191044
rect 579796 190988 579806 191044
rect 579740 190456 579796 190988
rect 262098 189980 262108 190036
rect 262164 189980 268072 190036
rect 331912 189980 336028 190036
rect 336084 189980 336094 190036
rect 61880 189756 73052 189812
rect 73108 189756 73118 189812
rect 185864 189756 189532 189812
rect 189588 189756 189598 189812
rect 247912 189756 257852 189812
rect 257908 189756 257918 189812
rect 472098 189756 472108 189812
rect 472164 189756 476056 189812
rect 517944 189756 519148 189812
rect 519204 189756 519214 189812
rect 579880 189756 583436 189812
rect 583492 189756 583502 189812
rect 263778 189420 263788 189476
rect 263844 189420 268072 189476
rect 331912 189420 347788 189476
rect 347844 189420 347854 189476
rect 123928 189084 126812 189140
rect 126868 189084 126878 189140
rect 204866 189084 204876 189140
rect 204932 189084 206136 189140
rect 247912 189084 258076 189140
rect 258132 189084 258142 189140
rect 393960 189084 396620 189140
rect 396676 189084 396686 189140
rect 579880 189084 581308 189140
rect 581364 189084 581374 189140
rect 455410 188972 455420 189028
rect 455476 188972 455486 189028
rect 263218 188860 263228 188916
rect 263284 188860 268072 188916
rect 331912 188860 350364 188916
rect 350420 188860 350430 188916
rect 20076 188244 20132 188440
rect 61880 188412 74732 188468
rect 74788 188412 74798 188468
rect 123928 188412 134428 188468
rect 134484 188412 134494 188468
rect 140914 188412 140924 188468
rect 140980 188412 144088 188468
rect 346098 188412 346108 188468
rect 346164 188412 352072 188468
rect 393960 188412 396844 188468
rect 396900 188412 396910 188468
rect 455420 188440 455476 188972
rect 263890 188300 263900 188356
rect 263956 188300 268072 188356
rect 331912 188300 338492 188356
rect 338548 188300 338558 188356
rect 20066 188188 20076 188244
rect 20132 188188 20142 188244
rect 82114 187740 82124 187796
rect 82180 187740 82190 187796
rect 140578 187740 140588 187796
rect 140644 187740 144088 187796
rect 185864 187740 197484 187796
rect 197540 187740 197550 187796
rect 203074 187740 203084 187796
rect 203140 187740 206136 187796
rect 256274 187740 256284 187796
rect 256340 187740 268072 187796
rect 331912 187740 352044 187796
rect 352100 187740 352110 187796
rect 263106 187180 263116 187236
rect 263172 187180 268072 187236
rect 331912 187180 350588 187236
rect 350644 187180 350654 187236
rect 61880 187068 64652 187124
rect 64708 187068 64718 187124
rect 82226 187068 82236 187124
rect 82292 187068 82302 187124
rect 203186 187068 203196 187124
rect 203252 187068 206136 187124
rect 247912 187068 251916 187124
rect 251972 187068 251982 187124
rect 472098 187068 472108 187124
rect 472164 187068 476056 187124
rect 579880 187068 583212 187124
rect 583268 187068 583278 187124
rect 258626 186620 258636 186676
rect 258692 186620 268072 186676
rect 331912 186620 342636 186676
rect 342692 186620 342702 186676
rect 82674 186396 82684 186452
rect 82740 186396 82750 186452
rect 393250 186396 393260 186452
rect 393316 186396 393326 186452
rect 455298 186396 455308 186452
rect 455364 186396 455374 186452
rect 467012 186396 476056 186452
rect 467012 186340 467068 186396
rect 456082 186284 456092 186340
rect 456148 186284 467068 186340
rect 265010 186060 265020 186116
rect 265076 186060 268072 186116
rect 331912 186060 341852 186116
rect 341908 186060 341918 186116
rect 263778 185500 263788 185556
rect 263844 185500 268072 185556
rect 331912 185500 346108 185556
rect 346164 185500 346174 185556
rect 248546 184940 248556 184996
rect 248612 184940 268072 184996
rect 331912 184940 351820 184996
rect 351876 184940 351886 184996
rect 249554 184380 249564 184436
rect 249620 184380 268072 184436
rect 331912 184380 336140 184436
rect 336196 184380 336206 184436
rect 263890 183820 263900 183876
rect 263956 183820 268072 183876
rect 331912 183820 350252 183876
rect 350308 183820 350318 183876
rect 261426 183260 261436 183316
rect 261492 183260 268072 183316
rect 331912 183260 335132 183316
rect 335188 183260 335198 183316
rect 264786 182700 264796 182756
rect 264852 182700 268072 182756
rect 331912 182700 352156 182756
rect 352212 182700 352222 182756
rect 261426 182140 261436 182196
rect 261492 182140 268072 182196
rect 331912 182140 340396 182196
rect 340452 182140 340462 182196
rect 517944 181692 521164 181748
rect 521220 181692 521230 181748
rect 264562 181580 264572 181636
rect 264628 181580 268072 181636
rect 331912 181580 348572 181636
rect 348628 181580 348638 181636
rect 259746 181020 259756 181076
rect 259812 181020 268072 181076
rect 331912 181020 338492 181076
rect 338548 181020 338558 181076
rect 257842 180460 257852 180516
rect 257908 180460 268072 180516
rect 331912 180460 350252 180516
rect 350308 180460 350318 180516
rect 252802 179900 252812 179956
rect 252868 179900 268072 179956
rect 331912 179900 345212 179956
rect 345268 179900 345278 179956
rect 262882 179340 262892 179396
rect 262948 179340 268072 179396
rect 331912 179340 335356 179396
rect 335412 179340 335422 179396
rect 595560 178920 597000 179144
rect 257842 178780 257852 178836
rect 257908 178780 268072 178836
rect 331912 178780 351932 178836
rect 351988 178780 351998 178836
rect 256386 178220 256396 178276
rect 256452 178220 268072 178276
rect 331912 178220 341852 178276
rect 341908 178220 341918 178276
rect -960 178052 480 178136
rect -960 177996 4396 178052
rect 4452 177996 4462 178052
rect 335122 177996 335132 178052
rect 335188 177996 338716 178052
rect 338772 177996 338782 178052
rect -960 177912 480 177996
rect 264674 177660 264684 177716
rect 264740 177660 268072 177716
rect 331912 177660 335356 177716
rect 335412 177660 335422 177716
rect 252802 177100 252812 177156
rect 252868 177100 268072 177156
rect 331912 177100 350252 177156
rect 350308 177100 350318 177156
rect 257954 176540 257964 176596
rect 258020 176540 268072 176596
rect 331912 176540 334460 176596
rect 334516 176540 334526 176596
rect 517944 176316 518252 176372
rect 518308 176316 518318 176372
rect 263778 175980 263788 176036
rect 263844 175980 268072 176036
rect 331912 175980 348572 176036
rect 348628 175980 348638 176036
rect 249554 175420 249564 175476
rect 249620 175420 268072 175476
rect 331912 175420 341852 175476
rect 341908 175420 341918 175476
rect 256274 174860 256284 174916
rect 256340 174860 268072 174916
rect 331912 174860 351932 174916
rect 351988 174860 351998 174916
rect 186498 174300 186508 174356
rect 186564 174300 268072 174356
rect 331912 174300 474572 174356
rect 474628 174300 474638 174356
rect 206098 173964 206108 174020
rect 206164 173964 263788 174020
rect 263844 173964 263854 174020
rect 335234 173964 335244 174020
rect 335300 173964 393932 174020
rect 393988 173964 393998 174020
rect 62066 173852 62076 173908
rect 62132 173852 264684 173908
rect 264740 173852 264750 173908
rect 334450 173852 334460 173908
rect 334516 173852 579628 173908
rect 579684 173852 579694 173908
rect 140802 173740 140812 173796
rect 140868 173740 268072 173796
rect 331912 173740 462812 173796
rect 462868 173740 462878 173796
rect 185602 173180 185612 173236
rect 185668 173180 268072 173236
rect 331912 173180 517468 173236
rect 517524 173180 517534 173236
rect 246418 172620 246428 172676
rect 246484 172620 268072 172676
rect 331912 172620 350364 172676
rect 350420 172620 350430 172676
rect 204866 172172 204876 172228
rect 204932 172172 264684 172228
rect 264740 172172 264750 172228
rect 335346 172172 335356 172228
rect 335412 172172 533372 172228
rect 533428 172172 533438 172228
rect 261426 172060 261436 172116
rect 261492 172060 268072 172116
rect 331912 172060 345436 172116
rect 345492 172060 345502 172116
rect 164882 171724 164892 171780
rect 164948 171724 199052 171780
rect 199108 171724 199118 171780
rect 230850 171724 230860 171780
rect 230916 171724 261212 171780
rect 261268 171724 261278 171780
rect 352146 171724 352156 171780
rect 352212 171724 368844 171780
rect 368900 171724 368910 171780
rect 102834 171612 102844 171668
rect 102900 171612 249676 171668
rect 249732 171612 249742 171668
rect 350578 171612 350588 171668
rect 350644 171612 375564 171668
rect 375620 171612 375630 171668
rect 414082 171612 414092 171668
rect 414148 171612 432124 171668
rect 432180 171612 432190 171668
rect 263778 171500 263788 171556
rect 263844 171500 268072 171556
rect 331912 171500 336028 171556
rect 336084 171500 336094 171556
rect 44930 171276 44940 171332
rect 44996 171276 141932 171332
rect 141988 171276 141998 171332
rect 166898 171276 166908 171332
rect 166964 171276 195692 171332
rect 195748 171276 195758 171332
rect 223458 171276 223468 171332
rect 223524 171276 259532 171332
rect 259588 171276 259598 171332
rect 345202 171276 345212 171332
rect 345268 171276 493500 171332
rect 493556 171276 493566 171332
rect 523282 171276 523292 171332
rect 523348 171276 571676 171332
rect 571732 171276 571742 171332
rect 41570 171164 41580 171220
rect 41636 171164 69692 171220
rect 69748 171164 69758 171220
rect 100146 171164 100156 171220
rect 100212 171164 133532 171220
rect 133588 171164 133598 171220
rect 229506 171164 229516 171220
rect 229572 171164 262892 171220
rect 262948 171164 262958 171220
rect 336802 171164 336812 171220
rect 336868 171164 376908 171220
rect 376964 171164 376974 171220
rect 398962 171164 398972 171220
rect 399028 171164 438508 171220
rect 438564 171164 438574 171220
rect 461122 171164 461132 171220
rect 461188 171164 496188 171220
rect 496244 171164 496254 171220
rect 228162 171052 228172 171108
rect 228228 171052 247772 171108
rect 247828 171052 247838 171108
rect 412402 171052 412412 171108
rect 412468 171052 440300 171108
rect 440356 171052 440366 171108
rect 464482 171052 464492 171108
rect 464548 171052 495516 171108
rect 495572 171052 495582 171108
rect 200722 170940 200732 170996
rect 200788 170940 268072 170996
rect 331912 170940 380492 170996
rect 380548 170940 380558 170996
rect 473106 170940 473116 170996
rect 473172 170940 494172 170996
rect 494228 170940 494238 170996
rect 474674 170828 474684 170884
rect 474740 170828 494844 170884
rect 494900 170828 494910 170884
rect 168354 170604 168364 170660
rect 168420 170604 186508 170660
rect 186564 170604 186574 170660
rect 167570 170492 167580 170548
rect 167636 170492 263788 170548
rect 263844 170492 263854 170548
rect 336018 170492 336028 170548
rect 336084 170492 520828 170548
rect 520884 170492 520894 170548
rect 187282 170380 187292 170436
rect 187348 170380 268072 170436
rect 331912 170380 461356 170436
rect 461412 170380 461422 170436
rect 188962 169820 188972 169876
rect 189028 169820 268072 169876
rect 331912 169820 472892 169876
rect 472948 169820 472958 169876
rect 226146 169596 226156 169652
rect 226212 169596 249452 169652
rect 249508 169596 249518 169652
rect 340274 169596 340284 169652
rect 340340 169596 562828 169652
rect 562884 169596 562894 169652
rect 35186 169484 35196 169540
rect 35252 169484 259644 169540
rect 259700 169484 259710 169540
rect 338706 169484 338716 169540
rect 338772 169484 556108 169540
rect 556164 169484 556174 169540
rect 39554 169372 39564 169428
rect 39620 169372 125132 169428
rect 125188 169372 125198 169428
rect 162866 169372 162876 169428
rect 162932 169372 261324 169428
rect 261380 169372 261390 169428
rect 338482 169372 338492 169428
rect 338548 169372 373548 169428
rect 373604 169372 373614 169428
rect 393922 169372 393932 169428
rect 393988 169372 559580 169428
rect 559636 169372 559646 169428
rect 43474 169260 43484 169316
rect 43540 169260 62076 169316
rect 62132 169260 62142 169316
rect 168242 169260 168252 169316
rect 168308 169260 263004 169316
rect 263060 169260 263070 169316
rect 263778 169260 263788 169316
rect 263844 169260 268072 169316
rect 331912 169260 338940 169316
rect 338996 169260 339006 169316
rect 345314 169260 345324 169316
rect 345380 169260 439068 169316
rect 439124 169260 439134 169316
rect 533474 169260 533484 169316
rect 533540 169260 558236 169316
rect 558292 169260 558302 169316
rect 162194 169148 162204 169204
rect 162260 169148 256172 169204
rect 256228 169148 256238 169204
rect 341954 169148 341964 169204
rect 342020 169148 432348 169204
rect 432404 169148 432414 169204
rect 536722 169148 536732 169204
rect 536788 169148 554876 169204
rect 554932 169148 554942 169204
rect 225474 169036 225484 169092
rect 225540 169036 252924 169092
rect 252980 169036 252990 169092
rect 352034 169036 352044 169092
rect 352100 169036 377580 169092
rect 377636 169036 377646 169092
rect 38546 168924 38556 168980
rect 38612 168924 263228 168980
rect 263284 168924 263294 168980
rect 263890 168700 263900 168756
rect 263956 168700 268072 168756
rect 331912 168700 334460 168756
rect 334516 168700 334526 168756
rect 263778 168140 263788 168196
rect 263844 168140 268072 168196
rect 331912 168140 336924 168196
rect 336980 168140 336990 168196
rect 197362 167580 197372 167636
rect 197428 167580 268072 167636
rect 331912 167580 519148 167636
rect 519204 167580 519214 167636
rect 334450 167132 334460 167188
rect 334516 167132 493500 167188
rect 493556 167132 493566 167188
rect 199042 167020 199052 167076
rect 199108 167020 268072 167076
rect 331912 167020 341964 167076
rect 342020 167020 342030 167076
rect 125122 166460 125132 166516
rect 125188 166460 268072 166516
rect 331912 166460 356972 166516
rect 357028 166460 357038 166516
rect 130162 165900 130172 165956
rect 130228 165900 268072 165956
rect 331912 165900 414092 165956
rect 414148 165900 414158 165956
rect 595560 165704 597000 165928
rect 204194 165452 204204 165508
rect 204260 165452 263788 165508
rect 263844 165452 263854 165508
rect 261538 165340 261548 165396
rect 261604 165340 268072 165396
rect 331912 165340 455308 165396
rect 455364 165340 455374 165396
rect 262994 164780 263004 164836
rect 263060 164780 268072 164836
rect 331912 164780 338604 164836
rect 338660 164780 338670 164836
rect 127138 164220 127148 164276
rect 127204 164220 268072 164276
rect 331912 164220 398972 164276
rect 399028 164220 399038 164276
rect -960 163800 480 164024
rect 195682 163772 195692 163828
rect 195748 163772 263788 163828
rect 263844 163772 263854 163828
rect 341842 163772 341852 163828
rect 341908 163772 582988 163828
rect 583044 163772 583054 163828
rect 126914 163660 126924 163716
rect 126980 163660 268072 163716
rect 331912 163660 410732 163716
rect 410788 163660 410798 163716
rect 127362 163100 127372 163156
rect 127428 163100 268072 163156
rect 331912 163100 452732 163156
rect 452788 163100 452798 163156
rect 127250 162540 127260 162596
rect 127316 162540 268072 162596
rect 331912 162540 457772 162596
rect 457828 162540 457838 162596
rect 192322 162092 192332 162148
rect 192388 162092 263900 162148
rect 263956 162092 263966 162148
rect 341842 162092 341852 162148
rect 341908 162092 556892 162148
rect 556948 162092 556958 162148
rect 135202 161980 135212 162036
rect 135268 161980 268072 162036
rect 331912 161980 456092 162036
rect 456148 161980 456158 162036
rect 126802 161420 126812 161476
rect 126868 161420 268072 161476
rect 331912 161420 412412 161476
rect 412468 161420 412478 161476
rect 127474 160860 127484 160916
rect 127540 160860 268072 160916
rect 331912 160860 407372 160916
rect 407428 160860 407438 160916
rect 338930 160524 338940 160580
rect 338996 160524 520940 160580
rect 520996 160524 521006 160580
rect 230178 160412 230188 160468
rect 230244 160412 256284 160468
rect 256340 160412 256350 160468
rect 340386 160412 340396 160468
rect 340452 160412 557564 160468
rect 557620 160412 557630 160468
rect 125234 160300 125244 160356
rect 125300 160300 268072 160356
rect 331912 160300 390572 160356
rect 390628 160300 390638 160356
rect 127026 159740 127036 159796
rect 127092 159740 268072 159796
rect 331912 159740 414204 159796
rect 414260 159740 414270 159796
rect 88050 159180 88060 159236
rect 88116 159180 268072 159236
rect 331912 159180 410844 159236
rect 410900 159180 410910 159236
rect 341954 158844 341964 158900
rect 342020 158844 494172 158900
rect 494228 158844 494238 158900
rect 228162 158732 228172 158788
rect 228228 158732 257964 158788
rect 258020 158732 258030 158788
rect 335346 158732 335356 158788
rect 335412 158732 581308 158788
rect 581364 158732 581374 158788
rect 64866 158620 64876 158676
rect 64932 158620 268072 158676
rect 331912 158620 352044 158676
rect 352100 158620 352110 158676
rect 81442 158060 81452 158116
rect 81508 158060 268072 158116
rect 331912 158060 395612 158116
rect 395668 158060 395678 158116
rect 64978 157500 64988 157556
rect 65044 157500 268072 157556
rect 331912 157500 390460 157556
rect 390516 157500 390526 157556
rect 390562 157276 390572 157332
rect 390628 157276 459004 157332
rect 459060 157276 459070 157332
rect 338594 157164 338604 157220
rect 338660 157164 410844 157220
rect 410900 157164 410910 157220
rect 228834 157052 228844 157108
rect 228900 157052 259756 157108
rect 259812 157052 259822 157108
rect 348562 157052 348572 157108
rect 348628 157052 583212 157108
rect 583268 157052 583278 157108
rect 64754 156940 64764 156996
rect 64820 156940 268072 156996
rect 331912 156940 395724 156996
rect 395780 156940 395790 156996
rect 18162 156380 18172 156436
rect 18228 156380 268072 156436
rect 331912 156380 341852 156436
rect 341908 156380 341918 156436
rect 69682 155820 69692 155876
rect 69748 155820 268072 155876
rect 331912 155820 357196 155876
rect 357252 155820 357262 155876
rect 356962 155596 356972 155652
rect 357028 155596 458780 155652
rect 458836 155596 458846 155652
rect 338482 155484 338492 155540
rect 338548 155484 535052 155540
rect 535108 155484 535118 155540
rect 351922 155372 351932 155428
rect 351988 155372 583100 155428
rect 583156 155372 583166 155428
rect 74722 155260 74732 155316
rect 74788 155260 268072 155316
rect 331912 155260 395836 155316
rect 395892 155260 395902 155316
rect 64642 154700 64652 154756
rect 64708 154700 268072 154756
rect 331912 154700 392252 154756
rect 392308 154700 392318 154756
rect 133522 154140 133532 154196
rect 133588 154140 268072 154196
rect 331912 154140 336028 154196
rect 336084 154140 336094 154196
rect 263778 153580 263788 153636
rect 263844 153580 268072 153636
rect 331912 153580 340284 153636
rect 340340 153580 340350 153636
rect 264674 153020 264684 153076
rect 264740 153020 268072 153076
rect 331912 153020 339276 153076
rect 339332 153020 339342 153076
rect 595560 152516 597000 152712
rect 42242 152460 42252 152516
rect 42308 152460 268072 152516
rect 331884 152404 331940 152488
rect 340162 152460 340172 152516
rect 340228 152488 597000 152516
rect 340228 152460 595672 152488
rect 331884 152348 372652 152404
rect 372708 152348 372718 152404
rect 339266 152124 339276 152180
rect 339332 152124 376908 152180
rect 376964 152124 376974 152180
rect 380482 152124 380492 152180
rect 380548 152124 473004 152180
rect 473060 152124 473070 152180
rect 73042 152012 73052 152068
rect 73108 152012 263788 152068
rect 263844 152012 263854 152068
rect 351922 152012 351932 152068
rect 351988 152012 556220 152068
rect 556276 152012 556286 152068
rect 62962 151900 62972 151956
rect 63028 151900 268072 151956
rect 331912 151900 338492 151956
rect 338548 151900 338558 151956
rect 263778 151340 263788 151396
rect 263844 151340 268072 151396
rect 331912 151340 396508 151396
rect 396564 151340 396574 151396
rect 261314 150780 261324 150836
rect 261380 150780 268072 150836
rect 331912 150780 536732 150836
rect 536788 150780 536798 150836
rect 162866 150668 162876 150724
rect 162932 150668 246428 150724
rect 246484 150668 246494 150724
rect 105522 150556 105532 150612
rect 105588 150556 261548 150612
rect 261604 150556 261614 150612
rect 81442 150444 81452 150500
rect 81508 150444 263788 150500
rect 263844 150444 263854 150500
rect 4610 150332 4620 150388
rect 4676 150332 205772 150388
rect 205828 150332 205838 150388
rect 336018 150332 336028 150388
rect 336084 150332 372876 150388
rect 372932 150332 372942 150388
rect 259970 150220 259980 150276
rect 260036 150220 268072 150276
rect 331912 150220 526652 150276
rect 526708 150220 526718 150276
rect -960 149716 480 149912
rect -960 149688 4396 149716
rect 392 149660 4396 149688
rect 4452 149660 4462 149716
rect 259746 149660 259756 149716
rect 259812 149660 268072 149716
rect 331912 149660 524972 149716
rect 525028 149660 525038 149716
rect 237682 149100 237692 149156
rect 237748 149100 268072 149156
rect 331912 149100 523292 149156
rect 523348 149100 523358 149156
rect 226146 148540 226156 148596
rect 226212 148540 268072 148596
rect 331912 148540 449372 148596
rect 449428 148540 449438 148596
rect 268044 147924 268100 148008
rect 331912 147980 334460 148036
rect 334516 147980 334526 148036
rect 265132 147868 268100 147924
rect 265132 147812 265188 147868
rect 263106 147756 263116 147812
rect 263172 147756 265188 147812
rect 203074 147420 203084 147476
rect 203140 147420 268072 147476
rect 331912 147420 581532 147476
rect 581588 147420 581598 147476
rect 164210 147196 164220 147252
rect 164276 147196 185612 147252
rect 185668 147196 185678 147252
rect 229506 147196 229516 147252
rect 229572 147196 237692 147252
rect 237748 147196 237758 147252
rect 161522 147084 161532 147140
rect 161588 147084 261436 147140
rect 261492 147084 261502 147140
rect 372642 147084 372652 147140
rect 372708 147084 374220 147140
rect 374276 147084 374286 147140
rect 69682 146972 69692 147028
rect 69748 146972 264684 147028
rect 264740 146972 264750 147028
rect 334450 146972 334460 147028
rect 334516 146972 437612 147028
rect 437668 146972 437678 147028
rect 261202 146860 261212 146916
rect 261268 146860 268072 146916
rect 331912 146860 579740 146916
rect 579796 146860 579806 146916
rect 268044 146244 268100 146328
rect 331912 146300 581420 146356
rect 581476 146300 581486 146356
rect 263788 146188 268100 146244
rect 263788 146132 263844 146188
rect 259634 146076 259644 146132
rect 259700 146076 263844 146132
rect 224802 145740 224812 145796
rect 224868 145740 268072 145796
rect 331912 145740 561596 145796
rect 561652 145740 561662 145796
rect 437602 145292 437612 145348
rect 437668 145292 560252 145348
rect 560308 145292 560318 145348
rect 203186 145180 203196 145236
rect 203252 145180 268072 145236
rect 331912 145180 581644 145236
rect 581700 145180 581710 145236
rect 38210 144956 38220 145012
rect 38276 144956 247772 145012
rect 247828 144956 247838 145012
rect 413970 144956 413980 145012
rect 414036 144956 435484 145012
rect 435540 144956 435550 145012
rect 106866 144844 106876 144900
rect 106932 144844 248108 144900
rect 248164 144844 248174 144900
rect 352706 144844 352716 144900
rect 352772 144844 434812 144900
rect 434868 144844 434878 144900
rect 204082 144732 204092 144788
rect 204148 144732 268100 144788
rect 348674 144732 348684 144788
rect 348740 144732 432796 144788
rect 432852 144732 432862 144788
rect 42914 144620 42924 144676
rect 42980 144620 249452 144676
rect 249508 144620 249518 144676
rect 268044 144648 268100 144732
rect 331912 144620 580412 144676
rect 580468 144620 580478 144676
rect 338594 144508 338604 144564
rect 338660 144508 437500 144564
rect 437556 144508 437566 144564
rect 475458 144508 475468 144564
rect 475524 144508 497532 144564
rect 497588 144508 497598 144564
rect 142818 144060 142828 144116
rect 142884 144060 268072 144116
rect 331912 144060 519260 144116
rect 519316 144060 519326 144116
rect 335234 143724 335244 143780
rect 335300 143724 352716 143780
rect 352772 143724 352782 143780
rect 357186 143724 357196 143780
rect 357252 143724 396620 143780
rect 396676 143724 396686 143780
rect 449362 143724 449372 143780
rect 449428 143724 535164 143780
rect 535220 143724 535230 143780
rect 102498 143612 102508 143668
rect 102564 143612 264684 143668
rect 264740 143612 264750 143668
rect 350354 143612 350364 143668
rect 350420 143612 472892 143668
rect 472948 143612 472958 143668
rect 199154 143500 199164 143556
rect 199220 143500 268072 143556
rect 331912 143500 340396 143556
rect 340452 143500 340462 143556
rect 350578 143164 350588 143220
rect 350644 143164 369516 143220
rect 369572 143164 369582 143220
rect 102834 143052 102844 143108
rect 102900 143052 256172 143108
rect 256228 143052 256238 143108
rect 351922 143052 351932 143108
rect 351988 143052 373548 143108
rect 373604 143052 373614 143108
rect 435026 143052 435036 143108
rect 435092 143052 500892 143108
rect 500948 143052 500958 143108
rect 206658 142940 206668 142996
rect 206724 142940 268072 142996
rect 331912 142940 334348 142996
rect 334404 142940 334414 142996
rect 352146 142940 352156 142996
rect 352212 142940 438172 142996
rect 438228 142940 438238 142996
rect 40898 142828 40908 142884
rect 40964 142828 247996 142884
rect 248052 142828 248062 142884
rect 342066 142828 342076 142884
rect 342132 142828 372204 142884
rect 372260 142828 372270 142884
rect 393138 142828 393148 142884
rect 393204 142828 498204 142884
rect 498260 142828 498270 142884
rect 392242 142716 392252 142772
rect 392308 142716 396956 142772
rect 397012 142716 397022 142772
rect 390562 142604 390572 142660
rect 390628 142604 396732 142660
rect 396788 142604 396798 142660
rect 334450 142492 334460 142548
rect 334516 142492 517692 142548
rect 517748 142492 517758 142548
rect 192322 142380 192332 142436
rect 192388 142380 268072 142436
rect 331912 142380 435036 142436
rect 435092 142380 435102 142436
rect 352034 142268 352044 142324
rect 352100 142268 368172 142324
rect 368228 142268 368238 142324
rect 197474 142156 197484 142212
rect 197540 142156 265412 142212
rect 345202 142156 345212 142212
rect 345268 142156 375564 142212
rect 375620 142156 375630 142212
rect 99474 142044 99484 142100
rect 99540 142044 256172 142100
rect 256228 142044 256238 142100
rect 262052 142044 265188 142100
rect 262052 141988 262108 142044
rect 265132 141988 265188 142044
rect 265356 141988 265412 142156
rect 336802 142044 336812 142100
rect 336868 142044 376236 142100
rect 376292 142044 376302 142100
rect 452722 142044 452732 142100
rect 452788 142044 458892 142100
rect 458948 142044 458958 142100
rect 98578 141932 98588 141988
rect 98644 141932 262108 141988
rect 265122 141932 265132 141988
rect 265188 141932 265198 141988
rect 265346 141932 265356 141988
rect 265412 141932 265422 141988
rect 350242 141932 350252 141988
rect 350308 141932 583436 141988
rect 583492 141932 583502 141988
rect 187394 141820 187404 141876
rect 187460 141820 268072 141876
rect 331912 141820 517580 141876
rect 517636 141820 517646 141876
rect 256162 141708 256172 141764
rect 256228 141708 264908 141764
rect 264964 141708 264974 141764
rect 334450 141708 334460 141764
rect 334516 141708 334526 141764
rect 351026 141708 351036 141764
rect 351092 141708 492828 141764
rect 492884 141708 492894 141764
rect 334460 141652 334516 141708
rect 265346 141596 265356 141652
rect 265412 141596 268100 141652
rect 268044 141288 268100 141596
rect 331884 141596 334516 141652
rect 331884 141288 331940 141596
rect 352034 140812 352044 140868
rect 352100 140812 396844 140868
rect 396900 140812 396910 140868
rect 200834 140700 200844 140756
rect 200900 140700 268072 140756
rect 331912 140700 335132 140756
rect 335188 140700 335198 140756
rect 335794 140700 335804 140756
rect 335860 140700 413980 140756
rect 414036 140700 414046 140756
rect 334338 140588 334348 140644
rect 334404 140588 464492 140644
rect 464548 140588 464558 140644
rect 334450 140476 334460 140532
rect 334516 140476 475468 140532
rect 475524 140476 475534 140532
rect 345426 140364 345436 140420
rect 345492 140364 521052 140420
rect 521108 140364 521118 140420
rect 345202 140252 345212 140308
rect 345268 140252 583324 140308
rect 583380 140252 583390 140308
rect 205762 140140 205772 140196
rect 205828 140140 268072 140196
rect 331912 140140 519372 140196
rect 519428 140140 519438 140196
rect 143602 139804 143612 139860
rect 143668 139804 264012 139860
rect 264068 139804 264078 139860
rect 136882 139692 136892 139748
rect 136948 139692 263900 139748
rect 263956 139692 263966 139748
rect 142034 139580 142044 139636
rect 142100 139580 268072 139636
rect 331912 139580 393148 139636
rect 393204 139580 393214 139636
rect 80322 139468 80332 139524
rect 80388 139468 250236 139524
rect 250292 139468 250302 139524
rect 140914 139356 140924 139412
rect 140980 139356 142828 139412
rect 142884 139356 142894 139412
rect 595560 139272 597000 139496
rect 199266 139132 199276 139188
rect 199332 139132 252700 139188
rect 252756 139132 252766 139188
rect 252924 139132 258748 139188
rect 252924 139076 252980 139132
rect 195794 139020 195804 139076
rect 195860 139020 252980 139076
rect 258692 139076 258748 139132
rect 258692 139020 268072 139076
rect 331912 139020 334460 139076
rect 334516 139020 334526 139076
rect 252690 138908 252700 138964
rect 252756 138908 267148 138964
rect 267092 138852 267148 138908
rect 267092 138796 268100 138852
rect 189074 138572 189084 138628
rect 189140 138572 206668 138628
rect 206724 138572 206734 138628
rect 268044 138488 268100 138796
rect 331912 138460 351036 138516
rect 351092 138460 351102 138516
rect 263778 137900 263788 137956
rect 263844 137900 268072 137956
rect 331912 137900 350364 137956
rect 350420 137900 350430 137956
rect 248098 137340 248108 137396
rect 248164 137340 268072 137396
rect 331912 137340 335244 137396
rect 335300 137340 335310 137396
rect 263890 136780 263900 136836
rect 263956 136780 268072 136836
rect 331912 136780 338604 136836
rect 338660 136780 338670 136836
rect 123928 136668 127484 136724
rect 127540 136668 127550 136724
rect 264002 136220 264012 136276
rect 264068 136220 268072 136276
rect 331912 136220 348684 136276
rect 348740 136220 348750 136276
rect 392 135800 4508 135828
rect -960 135772 4508 135800
rect 4564 135772 4574 135828
rect -960 135576 480 135772
rect 256162 135660 256172 135716
rect 256228 135660 268072 135716
rect 331912 135660 352156 135716
rect 352212 135660 352222 135716
rect 393932 135324 396508 135380
rect 396564 135324 396574 135380
rect 265122 135100 265132 135156
rect 265188 135100 268072 135156
rect 331912 135100 335804 135156
rect 335860 135100 335870 135156
rect 393932 134680 393988 135324
rect 250226 134540 250236 134596
rect 250292 134540 268072 134596
rect 331912 134540 334460 134596
rect 334516 134540 334526 134596
rect 263890 133980 263900 134036
rect 263956 133980 268072 134036
rect 331912 133980 335356 134036
rect 335412 133980 335422 134036
rect 263778 133420 263788 133476
rect 263844 133420 268072 133476
rect 331912 133420 345212 133476
rect 345268 133420 345278 133476
rect 254482 132860 254492 132916
rect 254548 132860 268072 132916
rect 331912 132860 351932 132916
rect 351988 132860 351998 132916
rect 395826 132636 395836 132692
rect 395892 132636 397068 132692
rect 397124 132636 397134 132692
rect 264898 132300 264908 132356
rect 264964 132300 268072 132356
rect 331912 132300 334460 132356
rect 334516 132300 334526 132356
rect 263778 131740 263788 131796
rect 263844 131740 268072 131796
rect 331912 131740 334348 131796
rect 334404 131740 334414 131796
rect 264674 131180 264684 131236
rect 264740 131180 268072 131236
rect 331912 131180 338492 131236
rect 338548 131180 338558 131236
rect 264674 130620 264684 130676
rect 264740 130620 268072 130676
rect 331912 130620 341964 130676
rect 342020 130620 342030 130676
rect 263778 130060 263788 130116
rect 263844 130060 268072 130116
rect 331912 130060 342188 130116
rect 342244 130060 342254 130116
rect 263890 129500 263900 129556
rect 263956 129500 268072 129556
rect 331912 129500 336812 129556
rect 336868 129500 336878 129556
rect 341842 129276 341852 129332
rect 341908 129276 347788 129332
rect 347844 129276 347854 129332
rect 263890 128940 263900 128996
rect 263956 128940 268072 128996
rect 331912 128940 342076 128996
rect 342132 128940 342142 128996
rect 337652 128604 352044 128660
rect 352100 128604 352110 128660
rect 252914 128492 252924 128548
rect 252980 128492 264572 128548
rect 264628 128492 264638 128548
rect 337652 128436 337708 128604
rect 263778 128380 263788 128436
rect 263844 128380 268072 128436
rect 331912 128380 337708 128436
rect 352594 128380 352604 128436
rect 352660 128380 352670 128436
rect 352604 127988 352660 128380
rect 18386 127932 18396 127988
rect 18452 127932 20076 127988
rect 20132 127932 20142 127988
rect 141026 127932 141036 127988
rect 141092 127932 144060 127988
rect 144116 127932 144126 127988
rect 201618 127932 201628 127988
rect 201684 127932 206136 127988
rect 349346 127932 349356 127988
rect 349412 127960 352660 127988
rect 349412 127932 352632 127960
rect 473666 127932 473676 127988
rect 473732 127932 476028 127988
rect 476084 127932 476094 127988
rect 264002 127820 264012 127876
rect 264068 127820 268072 127876
rect 331912 127820 342636 127876
rect 342692 127820 342702 127876
rect 258066 127596 258076 127652
rect 258132 127596 263788 127652
rect 263844 127596 263854 127652
rect 18386 127260 18396 127316
rect 18452 127260 20104 127316
rect 82674 127260 82684 127316
rect 82740 127260 82750 127316
rect 263890 127260 263900 127316
rect 263956 127260 268072 127316
rect 331912 127260 341964 127316
rect 342020 127260 342030 127316
rect 530786 127260 530796 127316
rect 530852 127260 538104 127316
rect 579880 127260 582988 127316
rect 583044 127260 583054 127316
rect 20626 127148 20636 127204
rect 20692 127148 20702 127204
rect 20636 126616 20692 127148
rect 248098 126812 248108 126868
rect 248164 126812 263788 126868
rect 263844 126812 263854 126868
rect 263778 126700 263788 126756
rect 263844 126700 268072 126756
rect 331912 126700 334460 126756
rect 334516 126700 334526 126756
rect 61880 126588 64876 126644
rect 64932 126588 64942 126644
rect 123928 126588 127260 126644
rect 127316 126588 127326 126644
rect 185864 126588 199052 126644
rect 199108 126588 199118 126644
rect 247912 126588 257852 126644
rect 257908 126588 257918 126644
rect 393250 126588 393260 126644
rect 393316 126588 393326 126644
rect 472994 126588 473004 126644
rect 473060 126588 476056 126644
rect 517458 126588 517468 126644
rect 517524 126588 517534 126644
rect 579880 126588 581644 126644
rect 581700 126588 581710 126644
rect 248322 126140 248332 126196
rect 248388 126140 268072 126196
rect 331912 126140 350588 126196
rect 350644 126140 350654 126196
rect 595560 126056 597000 126280
rect 123928 125916 127372 125972
rect 127428 125916 127438 125972
rect 185864 125916 195692 125972
rect 195748 125916 195758 125972
rect 204866 125916 204876 125972
rect 204932 125916 206136 125972
rect 247912 125916 261324 125972
rect 261380 125916 261390 125972
rect 249442 125580 249452 125636
rect 249508 125580 268072 125636
rect 331912 125580 334460 125636
rect 334516 125580 334526 125636
rect 393372 125524 393428 125944
rect 411618 125916 411628 125972
rect 411684 125916 414120 125972
rect 517944 125916 519372 125972
rect 519428 125916 519438 125972
rect 579880 125916 583436 125972
rect 583492 125916 583502 125972
rect 82450 125468 82460 125524
rect 82516 125468 82526 125524
rect 393362 125468 393372 125524
rect 393428 125468 393438 125524
rect 61880 124572 69692 124628
rect 69748 124572 69758 124628
rect 82460 124600 82516 125468
rect 185864 125244 192332 125300
rect 192388 125244 192398 125300
rect 206098 125244 206108 125300
rect 206164 125244 206174 125300
rect 247912 125244 252812 125300
rect 252868 125244 252878 125300
rect 524962 125244 524972 125300
rect 525028 125244 538104 125300
rect 579880 125244 581532 125300
rect 581588 125244 581598 125300
rect 455410 125132 455420 125188
rect 455476 125132 455486 125188
rect 263778 125020 263788 125076
rect 263844 125020 268072 125076
rect 331912 125020 345212 125076
rect 345268 125020 345278 125076
rect 140802 124572 140812 124628
rect 140868 124572 144088 124628
rect 185864 124572 188972 124628
rect 189028 124572 189038 124628
rect 455420 124600 455476 125132
rect 523282 124572 523292 124628
rect 523348 124572 538104 124628
rect 579880 124572 583212 124628
rect 583268 124572 583278 124628
rect 264786 124460 264796 124516
rect 264852 124460 268072 124516
rect 331912 124460 351932 124516
rect 351988 124460 351998 124516
rect 61852 124012 81452 124068
rect 81508 124012 81518 124068
rect 393932 124012 396732 124068
rect 396788 124012 396798 124068
rect 61852 123928 61908 124012
rect 80322 123900 80332 123956
rect 80388 123900 82068 123956
rect 140914 123900 140924 123956
rect 140980 123900 144088 123956
rect 203074 123900 203084 123956
rect 203140 123900 206136 123956
rect 264674 123900 264684 123956
rect 264740 123900 268072 123956
rect 331912 123900 345324 123956
rect 345380 123900 345390 123956
rect 61880 123228 64204 123284
rect 64260 123228 64270 123284
rect 82012 123256 82068 123900
rect 247986 123452 247996 123508
rect 248052 123452 263900 123508
rect 263956 123452 263966 123508
rect 261426 123340 261436 123396
rect 261492 123340 268072 123396
rect 331912 123340 336812 123396
rect 336868 123340 336878 123396
rect 185864 123228 205772 123284
rect 205828 123228 205838 123284
rect 393932 123256 393988 124012
rect 455298 123900 455308 123956
rect 455364 123900 455374 123956
rect 464482 123900 464492 123956
rect 464548 123900 476056 123956
rect 579880 123900 581308 123956
rect 581364 123900 581374 123956
rect 526642 123228 526652 123284
rect 526708 123228 538104 123284
rect 579618 123228 579628 123284
rect 579684 123228 579694 123284
rect 251906 122780 251916 122836
rect 251972 122780 268072 122836
rect 331912 122780 352268 122836
rect 352324 122780 352334 122836
rect 141026 122668 141036 122724
rect 141092 122668 142044 122724
rect 142100 122668 142110 122724
rect 189756 122668 199164 122724
rect 199220 122668 199230 122724
rect 189756 122612 189812 122668
rect 82012 122500 82068 122584
rect 123928 122556 126924 122612
rect 126980 122556 126990 122612
rect 185864 122556 189812 122612
rect 247912 122556 259980 122612
rect 260036 122556 260046 122612
rect 80434 122444 80444 122500
rect 80500 122444 82068 122500
rect 393932 122500 393988 122584
rect 517944 122556 519260 122612
rect 519316 122556 519326 122612
rect 579880 122556 583324 122612
rect 583380 122556 583390 122612
rect 393932 122444 396844 122500
rect 396900 122444 396910 122500
rect 249442 122220 249452 122276
rect 249508 122220 268072 122276
rect 331912 122220 337036 122276
rect 337092 122220 337102 122276
rect 61880 121884 64764 121940
rect 64820 121884 64830 121940
rect 123928 121884 127148 121940
rect 127204 121884 127214 121940
rect 247912 121884 256396 121940
rect 256452 121884 256462 121940
rect 579880 121884 581420 121940
rect 581476 121884 581486 121940
rect -960 121464 480 121688
rect 259522 121660 259532 121716
rect 259588 121660 268072 121716
rect 331912 121660 351820 121716
rect 351876 121660 351886 121716
rect 18162 121212 18172 121268
rect 18228 121212 20104 121268
rect 61880 121212 64988 121268
rect 65044 121212 65054 121268
rect 185864 121212 189084 121268
rect 189140 121212 189150 121268
rect 189522 121212 189532 121268
rect 189588 121212 197484 121268
rect 197540 121212 197550 121268
rect 247912 121212 259756 121268
rect 259812 121212 259822 121268
rect 411170 121212 411180 121268
rect 411236 121212 414120 121268
rect 455896 121212 458780 121268
rect 458836 121212 458846 121268
rect 579880 121212 583100 121268
rect 583156 121212 583166 121268
rect 256162 121100 256172 121156
rect 256228 121100 268072 121156
rect 331912 121100 350252 121156
rect 350308 121100 350318 121156
rect 457762 121100 457772 121156
rect 457828 121100 458668 121156
rect 458724 121100 458734 121156
rect 259970 120876 259980 120932
rect 260036 120876 264684 120932
rect 264740 120876 264750 120932
rect 61880 120540 73836 120596
rect 73892 120540 73902 120596
rect 185864 120540 199276 120596
rect 199332 120540 199342 120596
rect 252802 120540 252812 120596
rect 252868 120540 268072 120596
rect 331912 120540 341852 120596
rect 341908 120540 341918 120596
rect 347778 120540 347788 120596
rect 347844 120540 352072 120596
rect 393932 120540 396620 120596
rect 396676 120540 396686 120596
rect 455896 120540 456988 120596
rect 457044 120540 457054 120596
rect 517944 120540 520828 120596
rect 520884 120540 520894 120596
rect 254482 119980 254492 120036
rect 254548 119980 268072 120036
rect 331912 119980 336924 120036
rect 336980 119980 336990 120036
rect 61880 119868 64204 119924
rect 64260 119868 64270 119924
rect 123928 119868 127036 119924
rect 127092 119868 127102 119924
rect 203186 119868 203196 119924
rect 203252 119868 206136 119924
rect 247912 119868 261212 119924
rect 261268 119868 261278 119924
rect 342178 119868 342188 119924
rect 342244 119868 352072 119924
rect 393932 119896 393988 120540
rect 455298 120316 455308 120372
rect 455364 120316 455374 120372
rect 455308 119896 455364 120316
rect 462802 120092 462812 120148
rect 462868 120092 472108 120148
rect 472164 120092 472174 120148
rect 461346 119868 461356 119924
rect 461412 119868 476056 119924
rect 517944 119868 521052 119924
rect 521108 119868 521118 119924
rect 535154 119868 535164 119924
rect 535220 119868 538104 119924
rect 517682 119756 517692 119812
rect 517748 119756 517758 119812
rect 579730 119756 579740 119812
rect 579796 119756 579806 119812
rect 264898 119420 264908 119476
rect 264964 119420 268072 119476
rect 331912 119420 348684 119476
rect 348740 119420 348750 119476
rect 188188 119308 197372 119364
rect 197428 119308 197438 119364
rect 395714 119308 395724 119364
rect 395780 119308 395790 119364
rect 188188 119252 188244 119308
rect 395724 119252 395780 119308
rect 18386 119196 18396 119252
rect 18452 119196 20104 119252
rect 123928 119196 126812 119252
rect 126868 119196 126878 119252
rect 185836 119196 188244 119252
rect 204082 119196 204092 119252
rect 204148 119196 206164 119252
rect 20066 118524 20076 118580
rect 20132 118524 20142 118580
rect 123928 118524 136892 118580
rect 136948 118524 136958 118580
rect 185836 118552 185892 119196
rect 206108 118552 206164 119196
rect 393932 119196 395780 119252
rect 264786 118860 264796 118916
rect 264852 118860 268072 118916
rect 331912 118860 345324 118916
rect 345380 118860 345390 118916
rect 393932 118552 393988 119196
rect 396452 119140 396508 119252
rect 396564 119196 396574 119252
rect 404002 119196 404012 119252
rect 404068 119196 414120 119252
rect 455896 119196 456092 119252
rect 456148 119196 456158 119252
rect 517692 119224 517748 119756
rect 579740 119224 579796 119756
rect 395602 119084 395612 119140
rect 395668 119084 396508 119140
rect 580402 118860 580412 118916
rect 580468 118860 580478 118916
rect 580412 118580 580468 118860
rect 455896 118524 459004 118580
rect 459060 118524 459070 118580
rect 579852 118524 580468 118580
rect 141922 118412 141932 118468
rect 141988 118412 144116 118468
rect 61880 117852 64652 117908
rect 64708 117852 64718 117908
rect 144060 117880 144116 118412
rect 257842 118300 257852 118356
rect 257908 118300 268072 118356
rect 331912 118300 338716 118356
rect 338772 118300 338782 118356
rect 185864 117852 189532 117908
rect 189588 117852 189598 117908
rect 247912 117852 252924 117908
rect 252980 117852 252990 117908
rect 342626 117852 342636 117908
rect 342692 117852 352072 117908
rect 455896 117852 458892 117908
rect 458948 117852 458958 117908
rect 472098 117852 472108 117908
rect 472164 117852 476056 117908
rect 579852 117880 579908 118524
rect 263218 117740 263228 117796
rect 263284 117740 268072 117796
rect 331912 117740 342188 117796
rect 342244 117740 342254 117796
rect 393932 117404 396508 117460
rect 396564 117404 396574 117460
rect 247884 117292 261436 117348
rect 261492 117292 261502 117348
rect 123928 117180 143612 117236
rect 143668 117180 143678 117236
rect 185864 117180 195804 117236
rect 195860 117180 195870 117236
rect 247884 117208 247940 117292
rect 256274 117180 256284 117236
rect 256340 117180 268072 117236
rect 331912 117180 335244 117236
rect 335300 117180 335310 117236
rect 341954 117180 341964 117236
rect 342020 117180 352072 117236
rect 393932 117208 393988 117404
rect 455896 117180 458668 117236
rect 458724 117180 458734 117236
rect 472882 117180 472892 117236
rect 472948 117180 476056 117236
rect 517944 117180 520940 117236
rect 520996 117180 521006 117236
rect 535042 117180 535052 117236
rect 535108 117180 538104 117236
rect 393932 117068 397068 117124
rect 397124 117068 397134 117124
rect 261202 116620 261212 116676
rect 261268 116620 268072 116676
rect 331912 116620 338604 116676
rect 338660 116620 338670 116676
rect 61880 116508 64204 116564
rect 64260 116508 64270 116564
rect 141026 116508 141036 116564
rect 141092 116508 144088 116564
rect 393932 116536 393988 117068
rect 410834 116508 410844 116564
rect 410900 116508 414120 116564
rect 455634 116508 455644 116564
rect 455700 116508 455710 116564
rect 517570 116508 517580 116564
rect 517636 116508 517646 116564
rect 259634 116060 259644 116116
rect 259700 116060 268072 116116
rect 331912 116060 335692 116116
rect 335748 116060 335758 116116
rect 393932 115780 393988 115864
rect 517944 115836 519148 115892
rect 519204 115836 519214 115892
rect 393932 115724 396956 115780
rect 397012 115724 397022 115780
rect 249666 115500 249676 115556
rect 249732 115500 268072 115556
rect 331912 115500 345212 115556
rect 345268 115500 345278 115556
rect 252914 114940 252924 114996
rect 252980 114940 268072 114996
rect 331912 114940 342076 114996
rect 342132 114940 342142 114996
rect 247912 114492 262892 114548
rect 262948 114492 262958 114548
rect 261426 114380 261436 114436
rect 261492 114380 268072 114436
rect 331912 114380 352044 114436
rect 352100 114380 352110 114436
rect 262882 113820 262892 113876
rect 262948 113820 268072 113876
rect 331912 113820 334348 113876
rect 334404 113820 334414 113876
rect 247874 113372 247884 113428
rect 247940 113372 264908 113428
rect 264964 113372 264974 113428
rect 335346 113372 335356 113428
rect 335412 113372 346892 113428
rect 346948 113372 346958 113428
rect 258066 113260 258076 113316
rect 258132 113260 268072 113316
rect 331912 113260 348684 113316
rect 348740 113260 348750 113316
rect 587122 113036 587132 113092
rect 587188 113064 595672 113092
rect 587188 113036 597000 113064
rect 335682 112812 335692 112868
rect 335748 112812 340172 112868
rect 340228 112812 340238 112868
rect 595560 112840 597000 113036
rect 256162 112700 256172 112756
rect 256228 112700 268072 112756
rect 331912 112700 335132 112756
rect 335188 112700 335198 112756
rect 263778 112140 263788 112196
rect 263844 112140 268072 112196
rect 331912 112140 335468 112196
rect 335524 112140 335534 112196
rect 264674 111580 264684 111636
rect 264740 111580 268072 111636
rect 331912 111580 338492 111636
rect 338548 111580 338558 111636
rect 261314 111020 261324 111076
rect 261380 111020 268072 111076
rect 331912 111020 340508 111076
rect 340564 111020 340574 111076
rect 253026 110460 253036 110516
rect 253092 110460 268072 110516
rect 331912 110460 335356 110516
rect 335412 110460 335422 110516
rect 335122 110012 335132 110068
rect 335188 110012 343532 110068
rect 343588 110012 343598 110068
rect 249442 109900 249452 109956
rect 249508 109900 268072 109956
rect 331912 109900 350364 109956
rect 350420 109900 350430 109956
rect 264114 109340 264124 109396
rect 264180 109340 268072 109396
rect 331912 109340 338940 109396
rect 338996 109340 339006 109396
rect 259522 109228 259532 109284
rect 259588 109228 263788 109284
rect 263844 109228 263854 109284
rect 265122 108780 265132 108836
rect 265188 108780 268072 108836
rect 331912 108780 345436 108836
rect 345492 108780 345502 108836
rect 248098 108332 248108 108388
rect 248164 108332 264796 108388
rect 264852 108332 264862 108388
rect 265010 108220 265020 108276
rect 265076 108220 268072 108276
rect 331912 108220 341852 108276
rect 341908 108220 341918 108276
rect 257954 107660 257964 107716
rect 258020 107660 268072 107716
rect 331912 107660 350476 107716
rect 350532 107660 350542 107716
rect -960 107380 480 107576
rect 334338 107436 334348 107492
rect 334404 107436 336812 107492
rect 336868 107436 336878 107492
rect -960 107352 4284 107380
rect 392 107324 4284 107352
rect 4340 107324 4350 107380
rect 259746 107100 259756 107156
rect 259812 107100 268072 107156
rect 331912 107100 352492 107156
rect 352548 107100 352558 107156
rect 256386 106540 256396 106596
rect 256452 106540 268072 106596
rect 331912 106540 335916 106596
rect 335972 106540 335982 106596
rect 261314 105980 261324 106036
rect 261380 105980 268072 106036
rect 331912 105980 340396 106036
rect 340452 105980 340462 106036
rect 258178 105420 258188 105476
rect 258244 105420 268072 105476
rect 331912 105420 345548 105476
rect 345604 105420 345614 105476
rect 262882 105308 262892 105364
rect 262948 105308 265020 105364
rect 265076 105308 265086 105364
rect 247762 104972 247772 105028
rect 247828 104972 264684 105028
rect 264740 104972 264750 105028
rect 263778 104860 263788 104916
rect 263844 104860 268072 104916
rect 331912 104860 348572 104916
rect 348628 104860 348638 104916
rect 263890 104300 263900 104356
rect 263956 104300 268072 104356
rect 331912 104300 351148 104356
rect 351204 104300 351214 104356
rect 264002 103740 264012 103796
rect 264068 103740 268072 103796
rect 331912 103740 350476 103796
rect 350532 103740 350542 103796
rect 133522 103292 133532 103348
rect 133588 103292 263788 103348
rect 263844 103292 263854 103348
rect 335234 103292 335244 103348
rect 335300 103292 530012 103348
rect 530068 103292 530078 103348
rect 264562 103180 264572 103236
rect 264628 103180 268072 103236
rect 331912 103180 353612 103236
rect 353668 103180 353678 103236
rect 195682 103068 195692 103124
rect 195748 103068 264124 103124
rect 264180 103068 264190 103124
rect 263778 102620 263788 102676
rect 263844 102620 268072 102676
rect 331912 102620 351932 102676
rect 351988 102620 351998 102676
rect 160850 101724 160860 101780
rect 160916 101724 187404 101780
rect 187460 101724 187470 101780
rect 230178 101724 230188 101780
rect 230244 101724 257852 101780
rect 257908 101724 257918 101780
rect 268044 101668 268100 102088
rect 331912 102060 334460 102116
rect 334516 102060 334526 102116
rect 410834 101948 410844 102004
rect 410900 101948 422044 102004
rect 422100 101948 422110 102004
rect 340274 101836 340284 101892
rect 340340 101836 368172 101892
rect 368228 101836 368238 101892
rect 412402 101836 412412 101892
rect 412468 101836 429436 101892
rect 429492 101836 429502 101892
rect 338482 101724 338492 101780
rect 338548 101724 368844 101780
rect 368900 101724 368910 101780
rect 398962 101724 398972 101780
rect 399028 101724 434140 101780
rect 434196 101724 434206 101780
rect 43652 101612 74732 101668
rect 74788 101612 74798 101668
rect 102834 101612 102844 101668
rect 102900 101612 125132 101668
rect 125188 101612 125198 101668
rect 136882 101612 136892 101668
rect 136948 101612 263900 101668
rect 263956 101612 263966 101668
rect 267698 101612 267708 101668
rect 267764 101612 268100 101668
rect 351138 101612 351148 101668
rect 351204 101612 411068 101668
rect 411124 101612 411134 101668
rect 414082 101612 414092 101668
rect 414148 101612 438844 101668
rect 438900 101612 438910 101668
rect 43586 101052 43596 101108
rect 43652 101052 43708 101612
rect 143602 101500 143612 101556
rect 143668 101500 268072 101556
rect 331912 101500 334572 101556
rect 334628 101500 334638 101556
rect 267698 101164 267708 101220
rect 267764 101164 267774 101220
rect 267708 101108 267764 101164
rect 45602 101052 45612 101108
rect 45668 101052 81452 101108
rect 81508 101052 81518 101108
rect 82002 101052 82012 101108
rect 82068 101052 267764 101108
rect 335458 101052 335468 101108
rect 335524 101052 517468 101108
rect 517524 101052 517534 101108
rect 536722 101052 536732 101108
rect 536788 101052 556892 101108
rect 556948 101052 556958 101108
rect 44258 100940 44268 100996
rect 44324 100940 133532 100996
rect 133588 100940 133598 100996
rect 160822 100940 160860 100996
rect 160916 100940 160926 100996
rect 165554 100940 165564 100996
rect 165620 100940 200844 100996
rect 200900 100940 200910 100996
rect 204082 100940 204092 100996
rect 204148 100940 268072 100996
rect 331912 100940 335244 100996
rect 335300 100940 335310 100996
rect 336914 100940 336924 100996
rect 336980 100940 498876 100996
rect 498932 100940 498942 100996
rect 37538 100828 37548 100884
rect 37604 100828 69692 100884
rect 69748 100828 69758 100884
rect 99474 100828 99484 100884
rect 99540 100828 263004 100884
rect 263060 100828 263070 100884
rect 335906 100828 335916 100884
rect 335972 100828 399196 100884
rect 399252 100828 399262 100884
rect 407362 100828 407372 100884
rect 407428 100828 444220 100884
rect 444276 100828 444286 100884
rect 472882 100828 472892 100884
rect 472948 100828 499548 100884
rect 499604 100828 499614 100884
rect 102806 100716 102844 100772
rect 102900 100716 102910 100772
rect 169586 100716 169596 100772
rect 169652 100716 187292 100772
rect 187348 100716 187358 100772
rect 230150 100716 230188 100772
rect 230244 100716 230254 100772
rect 232866 100716 232876 100772
rect 232932 100716 249564 100772
rect 249620 100716 249630 100772
rect 368134 100716 368172 100772
rect 368228 100716 368238 100772
rect 368806 100716 368844 100772
rect 368900 100716 368910 100772
rect 422006 100716 422044 100772
rect 422100 100716 422110 100772
rect 429398 100716 429436 100772
rect 429492 100716 429502 100772
rect 434102 100716 434140 100772
rect 434196 100716 434206 100772
rect 438806 100716 438844 100772
rect 438900 100716 438910 100772
rect 106866 100604 106876 100660
rect 106932 100604 130172 100660
rect 130228 100604 130238 100660
rect 170258 100604 170268 100660
rect 170324 100604 192332 100660
rect 192388 100604 192398 100660
rect 231522 100604 231532 100660
rect 231588 100604 252812 100660
rect 252868 100604 252878 100660
rect 341954 100604 341964 100660
rect 342020 100604 376908 100660
rect 376964 100604 376974 100660
rect 410722 100604 410732 100660
rect 410788 100604 435484 100660
rect 435540 100604 435550 100660
rect 474562 100604 474572 100660
rect 474628 100604 495516 100660
rect 495572 100604 495582 100660
rect 101490 100492 101500 100548
rect 101556 100492 254492 100548
rect 254548 100492 254558 100548
rect 350354 100492 350364 100548
rect 350420 100492 420028 100548
rect 420084 100492 420094 100548
rect 420466 100492 420476 100548
rect 420532 100492 500892 100548
rect 500948 100492 500958 100548
rect 249778 100380 249788 100436
rect 249844 100380 268072 100436
rect 331912 100380 338604 100436
rect 338660 100380 338670 100436
rect 414194 100268 414204 100324
rect 414260 100268 428764 100324
rect 428820 100268 428830 100324
rect 138562 99932 138572 99988
rect 138628 99932 264012 99988
rect 264068 99932 264078 99988
rect 334450 99932 334460 99988
rect 334516 99932 456988 99988
rect 457044 99932 457054 99988
rect 265010 99820 265020 99876
rect 265076 99820 268072 99876
rect 331912 99820 334348 99876
rect 334404 99820 334414 99876
rect 595560 99624 597000 99848
rect 264786 99260 264796 99316
rect 264852 99260 268072 99316
rect 331912 99260 334684 99316
rect 334740 99260 334750 99316
rect 42242 99036 42252 99092
rect 42308 99036 247996 99092
rect 248052 99036 248062 99092
rect 350242 99036 350252 99092
rect 350308 99036 564284 99092
rect 564340 99036 564350 99092
rect 38210 98924 38220 98980
rect 38276 98924 73052 98980
rect 73108 98924 73118 98980
rect 105522 98924 105532 98980
rect 105588 98924 258076 98980
rect 258132 98924 258142 98980
rect 348562 98924 348572 98980
rect 348628 98924 558908 98980
rect 558964 98924 558974 98980
rect 38882 98812 38892 98868
rect 38948 98812 62972 98868
rect 63028 98812 63038 98868
rect 104178 98812 104188 98868
rect 104244 98812 135212 98868
rect 135268 98812 135278 98868
rect 168914 98812 168924 98868
rect 168980 98812 204204 98868
rect 204260 98812 204270 98868
rect 227490 98812 227500 98868
rect 227556 98812 259644 98868
rect 259700 98812 259710 98868
rect 340386 98812 340396 98868
rect 340452 98812 492828 98868
rect 492884 98812 492894 98868
rect 533362 98812 533372 98868
rect 533428 98812 556220 98868
rect 556276 98812 556286 98868
rect 104850 98700 104860 98756
rect 104916 98700 125244 98756
rect 125300 98700 125310 98756
rect 166226 98700 166236 98756
rect 166292 98700 200732 98756
rect 200788 98700 200798 98756
rect 232194 98700 232204 98756
rect 232260 98700 263116 98756
rect 263172 98700 263182 98756
rect 263778 98700 263788 98756
rect 263844 98700 268072 98756
rect 331912 98700 341964 98756
rect 342020 98700 342030 98756
rect 343522 98700 343532 98756
rect 343588 98700 494172 98756
rect 494228 98700 494238 98756
rect 346882 98588 346892 98644
rect 346948 98588 430108 98644
rect 430164 98588 430174 98644
rect 200946 98252 200956 98308
rect 201012 98252 265132 98308
rect 265188 98252 265198 98308
rect 334338 98252 334348 98308
rect 334404 98252 394828 98308
rect 394884 98252 394894 98308
rect 78082 98140 78092 98196
rect 78148 98140 268072 98196
rect 331912 98140 334460 98196
rect 334516 98140 334526 98196
rect 135426 97580 135436 97636
rect 135492 97580 268072 97636
rect 331912 97580 340172 97636
rect 340228 97580 340238 97636
rect 334450 97132 334460 97188
rect 334516 97132 394940 97188
rect 394996 97132 395006 97188
rect 73042 97020 73052 97076
rect 73108 97020 268072 97076
rect 331912 97020 345212 97076
rect 345268 97020 345278 97076
rect 350466 96908 350476 96964
rect 350532 96908 438172 96964
rect 438228 96908 438238 96964
rect 351922 96796 351932 96852
rect 351988 96796 535164 96852
rect 535220 96796 535230 96852
rect 142706 96684 142716 96740
rect 142772 96684 264684 96740
rect 264740 96684 264750 96740
rect 342178 96684 342188 96740
rect 342244 96684 556892 96740
rect 556948 96684 556958 96740
rect 110002 96572 110012 96628
rect 110068 96572 263788 96628
rect 263844 96572 263854 96628
rect 338706 96572 338716 96628
rect 338772 96572 583436 96628
rect 583492 96572 583502 96628
rect 69682 96460 69692 96516
rect 69748 96460 268072 96516
rect 331912 96460 350252 96516
rect 350308 96460 350318 96516
rect 74722 95900 74732 95956
rect 74788 95900 268072 95956
rect 331912 95900 340284 95956
rect 340340 95900 340350 95956
rect 167346 95340 167356 95396
rect 167412 95340 268072 95396
rect 331912 95340 392252 95396
rect 392308 95340 392318 95396
rect 229506 95004 229516 95060
rect 229572 95004 256284 95060
rect 256340 95004 256350 95060
rect 334562 95004 334572 95060
rect 334628 95004 455308 95060
rect 455364 95004 455374 95060
rect 228162 94892 228172 94948
rect 228228 94892 261436 94948
rect 261492 94892 261502 94948
rect 340498 94892 340508 94948
rect 340564 94892 504252 94948
rect 504308 94892 504318 94948
rect 62962 94780 62972 94836
rect 63028 94780 268072 94836
rect 331912 94780 355292 94836
rect 355348 94780 355358 94836
rect 263778 94220 263788 94276
rect 263844 94220 268072 94276
rect 331912 94220 338492 94276
rect 338548 94220 338558 94276
rect 226706 93660 226716 93716
rect 226772 93660 268072 93716
rect 331912 93660 395612 93716
rect 395668 93660 395678 93716
rect -960 93268 480 93464
rect 73042 93324 73052 93380
rect 73108 93324 263788 93380
rect 263844 93324 263854 93380
rect 338930 93324 338940 93380
rect 338996 93324 521276 93380
rect 521332 93324 521342 93380
rect -960 93240 266252 93268
rect 392 93212 266252 93240
rect 266308 93212 266318 93268
rect 345314 93212 345324 93268
rect 345380 93212 554204 93268
rect 554260 93212 554270 93268
rect 257058 93100 257068 93156
rect 257124 93100 268072 93156
rect 331912 93100 338716 93156
rect 338772 93100 338782 93156
rect 230178 92540 230188 92596
rect 230244 92540 268072 92596
rect 331912 92540 524972 92596
rect 525028 92540 525038 92596
rect 261202 91980 261212 92036
rect 261268 91980 268072 92036
rect 331912 91980 523292 92036
rect 523348 91980 523358 92036
rect 188962 91868 188972 91924
rect 189028 91868 261436 91924
rect 261492 91868 261502 91924
rect 106194 91756 106204 91812
rect 106260 91756 258188 91812
rect 258244 91756 258254 91812
rect 81442 91644 81452 91700
rect 81508 91644 263788 91700
rect 263844 91644 263854 91700
rect 334674 91644 334684 91700
rect 334740 91644 396956 91700
rect 397012 91644 397022 91700
rect 4386 91532 4396 91588
rect 4452 91532 263116 91588
rect 263172 91532 263182 91588
rect 335346 91532 335356 91588
rect 335412 91532 519148 91588
rect 519204 91532 519214 91588
rect 263778 91420 263788 91476
rect 263844 91420 268072 91476
rect 331912 91420 461916 91476
rect 461972 91420 461982 91476
rect 249554 90860 249564 90916
rect 249620 90860 268072 90916
rect 331912 90860 579628 90916
rect 579684 90860 579694 90916
rect 227602 90300 227612 90356
rect 227668 90300 268072 90356
rect 331912 90300 464492 90356
rect 464548 90300 464558 90356
rect 202850 90188 202860 90244
rect 202916 90188 230188 90244
rect 230244 90188 230254 90244
rect 165554 90076 165564 90132
rect 165620 90076 253036 90132
rect 253092 90076 253102 90132
rect 42242 89964 42252 90020
rect 42308 89964 226716 90020
rect 226772 89964 226782 90020
rect 338594 89964 338604 90020
rect 338660 89964 372204 90020
rect 372260 89964 372270 90020
rect 69794 89852 69804 89908
rect 69860 89852 265020 89908
rect 265076 89852 265086 89908
rect 345426 89852 345436 89908
rect 345492 89852 520940 89908
rect 520996 89852 521006 89908
rect 225474 89740 225484 89796
rect 225540 89740 268072 89796
rect 331912 89740 581308 89796
rect 581364 89740 581374 89796
rect 252802 89180 252812 89236
rect 252868 89180 268072 89236
rect 331912 89180 432572 89236
rect 432628 89180 432638 89236
rect 225922 88620 225932 88676
rect 225988 88620 268072 88676
rect 331912 88620 581420 88676
rect 581476 88620 581486 88676
rect 168242 88396 168252 88452
rect 168308 88396 252924 88452
rect 252980 88396 252990 88452
rect 141922 88284 141932 88340
rect 141988 88284 264572 88340
rect 264628 88284 264638 88340
rect 345538 88284 345548 88340
rect 345604 88284 458668 88340
rect 458724 88284 458734 88340
rect 50306 88172 50316 88228
rect 50372 88172 257068 88228
rect 257124 88172 257134 88228
rect 352034 88172 352044 88228
rect 352100 88172 494844 88228
rect 494900 88172 494910 88228
rect 204866 88060 204876 88116
rect 204932 88060 268072 88116
rect 331912 88060 580412 88116
rect 580468 88060 580478 88116
rect 264898 87500 264908 87556
rect 264964 87500 268072 87556
rect 331912 87500 403228 87556
rect 403284 87500 403294 87556
rect 264562 86940 264572 86996
rect 264628 86940 268072 86996
rect 331912 86940 581532 86996
rect 581588 86940 581598 86996
rect 160850 86716 160860 86772
rect 160916 86716 249676 86772
rect 249732 86716 249742 86772
rect 104178 86604 104188 86660
rect 104244 86604 256396 86660
rect 256452 86604 256462 86660
rect 340386 86604 340396 86660
rect 340452 86604 458780 86660
rect 458836 86604 458846 86660
rect 74722 86492 74732 86548
rect 74788 86492 264796 86548
rect 264852 86492 264862 86548
rect 342066 86492 342076 86548
rect 342132 86492 498204 86548
rect 498260 86492 498270 86548
rect 205762 86380 205772 86436
rect 205828 86380 268072 86436
rect 331912 86380 579740 86436
rect 579796 86380 579806 86436
rect 595560 86408 597000 86632
rect 197362 85820 197372 85876
rect 197428 85820 268072 85876
rect 331912 85820 393932 85876
rect 393988 85820 393998 85876
rect 257954 85708 257964 85764
rect 258020 85708 263788 85764
rect 263844 85708 263854 85764
rect 140578 85260 140588 85316
rect 140644 85260 268072 85316
rect 331912 85260 499772 85316
rect 499828 85260 499838 85316
rect 41570 84924 41580 84980
rect 41636 84924 167356 84980
rect 167412 84924 167422 84980
rect 232194 84924 232204 84980
rect 232260 84924 263228 84980
rect 263284 84924 263294 84980
rect 335234 84924 335244 84980
rect 335300 84924 457100 84980
rect 457156 84924 457166 84980
rect 461906 84924 461916 84980
rect 461972 84924 560252 84980
rect 560308 84924 560318 84980
rect 126802 84812 126812 84868
rect 126868 84812 259756 84868
rect 259812 84812 259822 84868
rect 348674 84812 348684 84868
rect 348740 84812 472892 84868
rect 472948 84812 472958 84868
rect 167122 84700 167132 84756
rect 167188 84700 268072 84756
rect 331912 84700 375452 84756
rect 375508 84700 375518 84756
rect 199042 84140 199052 84196
rect 199108 84140 268072 84196
rect 331912 84140 462812 84196
rect 462868 84140 462878 84196
rect 140914 83580 140924 83636
rect 140980 83580 268072 83636
rect 331912 83580 461132 83636
rect 461188 83580 461198 83636
rect 146962 83020 146972 83076
rect 147028 83020 268072 83076
rect 331912 83020 519260 83076
rect 519316 83020 519326 83076
rect 145282 82460 145292 82516
rect 145348 82460 268072 82516
rect 331912 82460 517580 82516
rect 517636 82460 517646 82516
rect 187282 81900 187292 81956
rect 187348 81900 268072 81956
rect 331912 81900 407372 81956
rect 407428 81900 407438 81956
rect 403218 81452 403228 81508
rect 403284 81452 560924 81508
rect 560980 81452 560990 81508
rect 142034 81340 142044 81396
rect 142100 81340 268072 81396
rect 331912 81340 492156 81396
rect 492212 81340 492222 81396
rect 263778 80780 263788 80836
rect 263844 80780 268072 80836
rect 331912 80780 404796 80836
rect 404852 80780 404862 80836
rect 142594 80220 142604 80276
rect 142660 80220 268072 80276
rect 331912 80220 519372 80276
rect 519428 80220 519438 80276
rect 355282 79996 355292 80052
rect 355348 79996 379596 80052
rect 379652 79996 379662 80052
rect 350466 79884 350476 79940
rect 350532 79884 458892 79940
rect 458948 79884 458958 79940
rect 38882 79772 38892 79828
rect 38948 79772 135436 79828
rect 135492 79772 135502 79828
rect 162866 79772 162876 79828
rect 162932 79772 261324 79828
rect 261380 79772 261390 79828
rect 338594 79772 338604 79828
rect 338660 79772 583100 79828
rect 583156 79772 583166 79828
rect 144050 79660 144060 79716
rect 144116 79660 268072 79716
rect 331912 79660 518252 79716
rect 518308 79660 518318 79716
rect -960 79128 480 79352
rect 125122 79100 125132 79156
rect 125188 79100 268072 79156
rect 331912 79100 335916 79156
rect 335972 79100 335982 79156
rect 264674 78540 264684 78596
rect 264740 78540 268072 78596
rect 331912 78540 352044 78596
rect 352100 78540 352110 78596
rect 352482 78428 352492 78484
rect 352548 78428 436156 78484
rect 436212 78428 436222 78484
rect 203074 78316 203084 78372
rect 203140 78316 254492 78372
rect 254548 78316 254558 78372
rect 335906 78316 335916 78372
rect 335972 78316 371308 78372
rect 371364 78316 371374 78372
rect 404786 78316 404796 78372
rect 404852 78316 494172 78372
rect 494228 78316 494238 78372
rect 144274 78204 144284 78260
rect 144340 78204 263788 78260
rect 263844 78204 263854 78260
rect 352258 78204 352268 78260
rect 352324 78204 535388 78260
rect 535444 78204 535454 78260
rect 98802 78092 98812 78148
rect 98868 78092 257964 78148
rect 258020 78092 258030 78148
rect 348674 78092 348684 78148
rect 348740 78092 557564 78148
rect 557620 78092 557630 78148
rect 130162 77980 130172 78036
rect 130228 77980 268072 78036
rect 331912 77980 404012 78036
rect 404068 77980 404078 78036
rect 80210 77420 80220 77476
rect 80276 77420 268072 77476
rect 331912 77420 335132 77476
rect 335188 77420 335198 77476
rect 258178 77308 258188 77364
rect 258244 77308 264908 77364
rect 264964 77308 264974 77364
rect 188066 76860 188076 76916
rect 188132 76860 268072 76916
rect 331912 76860 457772 76916
rect 457828 76860 457838 76916
rect 134418 76300 134428 76356
rect 134484 76300 268072 76356
rect 331912 76300 402332 76356
rect 402388 76300 402398 76356
rect 263778 75740 263788 75796
rect 263844 75740 268072 75796
rect 331912 75740 334460 75796
rect 334516 75740 334526 75796
rect 82338 75180 82348 75236
rect 82404 75180 268072 75236
rect 331912 75180 334348 75236
rect 334404 75180 334414 75236
rect 371298 75068 371308 75124
rect 371364 75068 433468 75124
rect 433524 75068 433534 75124
rect 224130 74956 224140 75012
rect 224196 74956 228116 75012
rect 393922 74956 393932 75012
rect 393988 74956 497532 75012
rect 497588 74956 497598 75012
rect 100818 74844 100828 74900
rect 100884 74844 110012 74900
rect 110068 74844 110078 74900
rect 223458 74844 223468 74900
rect 223524 74844 225932 74900
rect 225988 74844 225998 74900
rect 228060 74788 228116 74956
rect 228834 74844 228844 74900
rect 228900 74844 248108 74900
rect 248164 74844 248174 74900
rect 375442 74844 375452 74900
rect 375508 74844 501564 74900
rect 501620 74844 501630 74900
rect 100146 74732 100156 74788
rect 100212 74732 134428 74788
rect 134484 74732 134494 74788
rect 163538 74732 163548 74788
rect 163604 74732 167132 74788
rect 167188 74732 167198 74788
rect 224802 74732 224812 74788
rect 224868 74732 227612 74788
rect 227668 74732 227678 74788
rect 228060 74732 247884 74788
rect 247940 74732 247950 74788
rect 252914 74732 252924 74788
rect 252980 74732 264572 74788
rect 264628 74732 264638 74788
rect 334450 74732 334460 74788
rect 334516 74732 399476 74788
rect 402322 74732 402332 74788
rect 402388 74732 432124 74788
rect 432180 74732 432190 74788
rect 432562 74732 432572 74788
rect 432628 74732 562268 74788
rect 562324 74732 562334 74788
rect 399420 74676 399476 74732
rect 105522 74620 105532 74676
rect 105588 74620 268072 74676
rect 331912 74620 398076 74676
rect 398132 74620 398142 74676
rect 399420 74620 402332 74676
rect 402388 74620 402398 74676
rect 499762 74620 499772 74676
rect 499828 74620 500892 74676
rect 500948 74620 500958 74676
rect 35522 74172 35532 74228
rect 35588 74172 248332 74228
rect 248388 74172 248398 74228
rect 348562 74172 348572 74228
rect 348628 74172 376908 74228
rect 376964 74172 376974 74228
rect 45602 74060 45612 74116
rect 45668 74060 83916 74116
rect 83972 74060 83982 74116
rect 135202 74060 135212 74116
rect 135268 74060 268072 74116
rect 331912 74060 334572 74116
rect 334628 74060 334638 74116
rect 352706 74060 352716 74116
rect 352772 74060 372876 74116
rect 372932 74060 372942 74116
rect 359538 73948 359548 74004
rect 359604 73948 368844 74004
rect 368900 73948 368910 74004
rect 102834 73500 102844 73556
rect 102900 73500 268072 73556
rect 331912 73500 334460 73556
rect 334516 73500 334526 73556
rect 348562 73500 348572 73556
rect 348628 73500 410732 73556
rect 410788 73500 410798 73556
rect 334338 73388 334348 73444
rect 334404 73388 455420 73444
rect 455476 73388 455486 73444
rect 203186 73276 203196 73332
rect 203252 73276 257852 73332
rect 257908 73276 257918 73332
rect 335122 73276 335132 73332
rect 335188 73276 519484 73332
rect 519540 73276 519550 73332
rect 595560 73220 597000 73416
rect 189074 73164 189084 73220
rect 189140 73164 258076 73220
rect 258132 73164 258142 73220
rect 333442 73164 333452 73220
rect 333508 73192 597000 73220
rect 333508 73164 595672 73192
rect 138674 73052 138684 73108
rect 138740 73052 263788 73108
rect 263844 73052 263854 73108
rect 337026 73052 337036 73108
rect 337092 73052 535276 73108
rect 535332 73052 535342 73108
rect 81554 72940 81564 72996
rect 81620 72940 268072 72996
rect 331912 72940 456092 72996
rect 456148 72940 456158 72996
rect 45266 72380 45276 72436
rect 45332 72380 268072 72436
rect 331912 72380 335356 72436
rect 335412 72380 335422 72436
rect 392242 72156 392252 72212
rect 392308 72156 396620 72212
rect 396676 72156 396686 72212
rect 83906 71820 83916 71876
rect 83972 71820 268072 71876
rect 331912 71820 346892 71876
rect 346948 71820 346958 71876
rect 353602 71708 353612 71764
rect 353668 71708 459116 71764
rect 459172 71708 459182 71764
rect 334450 71596 334460 71652
rect 334516 71596 457212 71652
rect 457268 71596 457278 71652
rect 189410 71484 189420 71540
rect 189476 71484 249452 71540
rect 249508 71484 249518 71540
rect 350242 71484 350252 71540
rect 350308 71484 535500 71540
rect 535556 71484 535566 71540
rect 80322 71372 80332 71428
rect 80388 71372 188076 71428
rect 188132 71372 188142 71428
rect 189186 71372 189196 71428
rect 189252 71372 259644 71428
rect 259700 71372 259710 71428
rect 336914 71372 336924 71428
rect 336980 71372 583212 71428
rect 583268 71372 583278 71428
rect 63074 71260 63084 71316
rect 63140 71260 268072 71316
rect 331912 71260 393932 71316
rect 393988 71260 393998 71316
rect 64642 70700 64652 70756
rect 64708 70700 268072 70756
rect 331912 70700 359548 70756
rect 359604 70700 359614 70756
rect 371158 70700 371196 70756
rect 371252 70700 371262 70756
rect 352258 70588 352268 70644
rect 352324 70588 377580 70644
rect 377636 70588 377646 70644
rect 43810 70476 43820 70532
rect 43876 70476 252700 70532
rect 252756 70476 252766 70532
rect 341842 70476 341852 70532
rect 341908 70476 583324 70532
rect 583380 70476 583390 70532
rect 140802 70364 140812 70420
rect 140868 70364 146972 70420
rect 147028 70364 147038 70420
rect 246932 70252 258748 70308
rect 246932 70196 246988 70252
rect 20626 70140 20636 70196
rect 20692 70140 246988 70196
rect 258692 70196 258748 70252
rect 258692 70140 268072 70196
rect 331912 70140 393148 70196
rect 393204 70140 393214 70196
rect 252690 70028 252700 70084
rect 252756 70028 267148 70084
rect 267092 69972 267148 70028
rect 202962 69916 202972 69972
rect 203028 69916 252812 69972
rect 252868 69916 252878 69972
rect 267092 69916 268100 69972
rect 338482 69916 338492 69972
rect 338548 69916 521052 69972
rect 521108 69916 521118 69972
rect 189298 69804 189308 69860
rect 189364 69804 262892 69860
rect 262948 69804 262958 69860
rect 126914 69692 126924 69748
rect 126980 69692 261324 69748
rect 261380 69692 261390 69748
rect 268044 69608 268100 69916
rect 345314 69804 345324 69860
rect 345380 69804 535612 69860
rect 535668 69804 535678 69860
rect 336802 69692 336812 69748
rect 336868 69692 535836 69748
rect 535892 69692 535902 69748
rect 331912 69580 337036 69636
rect 337092 69580 337102 69636
rect 361172 69132 371196 69188
rect 371252 69132 371262 69188
rect 361172 69076 361228 69132
rect 76402 69020 76412 69076
rect 76468 69020 268072 69076
rect 331912 69020 361228 69076
rect 80434 68796 80444 68852
rect 80500 68796 82348 68852
rect 82404 68796 82414 68852
rect 140690 68796 140700 68852
rect 140756 68796 145292 68852
rect 145348 68796 145358 68852
rect 334450 68572 334460 68628
rect 334516 68572 395052 68628
rect 395108 68572 395118 68628
rect 19954 68460 19964 68516
rect 20020 68460 268072 68516
rect 331912 68460 352716 68516
rect 352772 68460 352782 68516
rect 398066 68236 398076 68292
rect 398132 68236 459004 68292
rect 459060 68236 459070 68292
rect 334562 68124 334572 68180
rect 334628 68124 400652 68180
rect 400708 68124 400718 68180
rect 76514 68012 76524 68068
rect 76580 68012 252812 68068
rect 252868 68012 252878 68068
rect 253036 68012 258748 68068
rect 350354 68012 350364 68068
rect 350420 68012 521164 68068
rect 521220 68012 521230 68068
rect 253036 67956 253092 68012
rect 20066 67900 20076 67956
rect 20132 67900 253092 67956
rect 258692 67956 258748 68012
rect 258692 67900 268072 67956
rect 331912 67900 346780 67956
rect 346836 67900 346846 67956
rect 393138 67900 393148 67956
rect 393204 67900 396732 67956
rect 396788 67900 396798 67956
rect 252802 67788 252812 67844
rect 252868 67788 267148 67844
rect 334450 67788 334460 67844
rect 334516 67788 334526 67844
rect 267092 67732 267148 67788
rect 334460 67732 334516 67788
rect 267092 67676 268100 67732
rect 268044 67368 268100 67676
rect 331884 67676 334516 67732
rect 331884 67368 331940 67676
rect 18274 67228 18284 67284
rect 18340 67228 20636 67284
rect 20692 67228 20702 67284
rect 349412 66892 352268 66948
rect 352324 66892 352334 66948
rect 248322 66780 248332 66836
rect 248388 66780 268072 66836
rect 331912 66780 348572 66836
rect 348628 66780 348638 66836
rect 349412 66388 349468 66892
rect 64754 66332 64764 66388
rect 64820 66332 76412 66388
rect 76468 66332 76478 66388
rect 331884 66332 349468 66388
rect 123928 66220 138572 66276
rect 138628 66220 138638 66276
rect 264898 66220 264908 66276
rect 264964 66220 268072 66276
rect 331884 66248 331940 66332
rect 340274 66220 340284 66276
rect 340340 66220 352072 66276
rect 142706 65548 142716 65604
rect 142772 65548 144088 65604
rect 185864 65548 189420 65604
rect 189476 65548 189486 65604
rect 203186 65548 203196 65604
rect 203252 65548 206136 65604
rect -960 65044 480 65240
rect -960 65016 4396 65044
rect 392 64988 4396 65016
rect 4452 64988 4462 65044
rect 395042 60396 395052 60452
rect 395108 60396 396844 60452
rect 396900 60396 396910 60452
rect 595560 59976 597000 60200
rect 335346 59612 335356 59668
rect 335412 59612 348572 59668
rect 348628 59612 348638 59668
rect 349318 57036 349356 57092
rect 349412 57036 349422 57092
rect 18358 56812 18396 56868
rect 18452 56812 20104 56868
rect 82572 56308 82628 56840
rect 203186 56812 203196 56868
rect 203252 56840 206136 56868
rect 203252 56812 206164 56840
rect 206108 56308 206164 56812
rect 352604 56308 352660 56840
rect 414652 56308 414708 56840
rect 82562 56252 82572 56308
rect 82628 56252 82638 56308
rect 123900 56252 143612 56308
rect 143668 56252 143678 56308
rect 206098 56252 206108 56308
rect 206164 56252 206174 56308
rect 352594 56252 352604 56308
rect 352660 56252 352670 56308
rect 414642 56252 414652 56308
rect 414708 56252 414718 56308
rect 123900 56168 123956 56252
rect 141026 56140 141036 56196
rect 141092 56140 144060 56196
rect 144116 56140 144126 56196
rect 204866 56140 204876 56196
rect 204932 56140 206136 56196
rect 473666 56140 473676 56196
rect 473732 56140 476056 56196
rect 534258 56140 534268 56196
rect 534324 56140 538104 56196
rect 20066 55468 20076 55524
rect 20132 55468 20142 55524
rect 123928 55468 138684 55524
rect 138740 55468 138750 55524
rect 185864 55468 195692 55524
rect 195748 55468 195758 55524
rect 411058 55468 411068 55524
rect 411124 55468 414120 55524
rect 455896 55468 457100 55524
rect 457156 55468 457166 55524
rect 579880 55468 581420 55524
rect 581476 55468 581486 55524
rect 123928 54796 141932 54852
rect 141988 54796 141998 54852
rect 185864 54796 189308 54852
rect 189364 54796 189374 54852
rect 400642 54796 400652 54852
rect 400708 54796 414120 54852
rect 455896 54796 458668 54852
rect 458724 54796 458734 54852
rect 535826 54796 535836 54852
rect 535892 54796 538104 54852
rect 579880 54796 581532 54852
rect 581588 54796 581598 54852
rect 80322 54124 80332 54180
rect 80388 54124 82040 54180
rect 123928 54124 126924 54180
rect 126980 54124 126990 54180
rect 140802 54124 140812 54180
rect 140868 54124 144088 54180
rect 185864 54124 188972 54180
rect 189028 54124 189038 54180
rect 202850 54124 202860 54180
rect 202916 54124 206136 54180
rect 346770 54124 346780 54180
rect 346836 54124 352072 54180
rect 393960 54124 396956 54180
rect 397012 54124 397022 54180
rect 455896 54124 458780 54180
rect 458836 54124 458846 54180
rect 61880 53452 76412 53508
rect 76468 53452 76478 53508
rect 140690 53452 140700 53508
rect 140756 53452 144088 53508
rect 203074 53452 203084 53508
rect 203140 53452 206136 53508
rect 247912 53452 256172 53508
rect 256228 53452 256238 53508
rect 393960 53452 396732 53508
rect 396788 53452 396798 53508
rect 455298 53452 455308 53508
rect 455364 53452 455374 53508
rect 517944 53452 521164 53508
rect 521220 53452 521230 53508
rect 393922 53228 393932 53284
rect 393988 53228 393998 53284
rect 455868 53228 459116 53284
rect 459172 53228 459182 53284
rect 4386 52892 4396 52948
rect 4452 52892 10892 52948
rect 10948 52892 10958 52948
rect 61880 52780 74732 52836
rect 74788 52780 74798 52836
rect 142594 52780 142604 52836
rect 142660 52780 144088 52836
rect 202962 52780 202972 52836
rect 203028 52780 206136 52836
rect 247912 52780 259532 52836
rect 259588 52780 259598 52836
rect 346882 52780 346892 52836
rect 346948 52780 352072 52836
rect 393932 52808 393988 53228
rect 402322 52780 402332 52836
rect 402388 52780 414120 52836
rect 455868 52808 455924 53228
rect 457762 52892 457772 52948
rect 457828 52892 457838 52948
rect 457772 52612 457828 52892
rect 462802 52780 462812 52836
rect 462868 52780 476056 52836
rect 517944 52780 521052 52836
rect 521108 52780 521118 52836
rect 523282 52780 523292 52836
rect 523348 52780 538104 52836
rect 579618 52780 579628 52836
rect 579684 52780 579694 52836
rect 455868 52556 457828 52612
rect 61880 52108 64764 52164
rect 64820 52108 64830 52164
rect 185864 52108 189196 52164
rect 189252 52108 189262 52164
rect 247912 52108 261212 52164
rect 261268 52108 261278 52164
rect 341954 52108 341964 52164
rect 342020 52108 352072 52164
rect 410722 52108 410732 52164
rect 410788 52108 414120 52164
rect 455868 52136 455924 52556
rect 517570 52108 517580 52164
rect 517636 52108 517646 52164
rect 535378 52108 535388 52164
rect 535444 52108 538104 52164
rect 579880 52108 583324 52164
rect 583380 52108 583390 52164
rect 395602 51996 395612 52052
rect 395668 51996 396508 52052
rect 396564 51996 396574 52052
rect 61880 51436 64652 51492
rect 64708 51436 64718 51492
rect 455896 51436 456988 51492
rect 457044 51436 457054 51492
rect 517944 51436 520940 51492
rect 520996 51436 521006 51492
rect 64306 51324 64316 51380
rect 64372 51324 73052 51380
rect 73108 51324 73118 51380
rect 64082 51212 64092 51268
rect 64148 51212 78092 51268
rect 78148 51212 78158 51268
rect 392 51128 4172 51156
rect -960 51100 4172 51128
rect 4228 51100 4238 51156
rect -960 50904 480 51100
rect 123928 50764 126812 50820
rect 126868 50764 126878 50820
rect 455896 50764 457212 50820
rect 457268 50764 457278 50820
rect 517944 50764 519148 50820
rect 519204 50764 519214 50820
rect 524962 50764 524972 50820
rect 525028 50764 538104 50820
rect 579730 50764 579740 50820
rect 579796 50764 579806 50820
rect 127586 50540 127596 50596
rect 127652 50540 130172 50596
rect 130228 50540 130238 50596
rect 61852 50204 81452 50260
rect 81508 50204 81518 50260
rect 61852 50120 61908 50204
rect 81554 50092 81564 50148
rect 81620 50092 82040 50148
rect 123928 50092 136892 50148
rect 136948 50092 136958 50148
rect 144274 50092 144284 50148
rect 144340 50092 144350 50148
rect 185864 50092 200956 50148
rect 201012 50092 201022 50148
rect 247912 50092 257964 50148
rect 258020 50092 258030 50148
rect 393960 50092 394940 50148
rect 394996 50092 395006 50148
rect 455896 50092 458892 50148
rect 458948 50092 458958 50148
rect 123928 49420 133532 49476
rect 133588 49420 133598 49476
rect 144050 49420 144060 49476
rect 144116 49420 144126 49476
rect 185864 49420 189084 49476
rect 189140 49420 189150 49476
rect 247912 49420 251916 49476
rect 251972 49420 251982 49476
rect 340162 49420 340172 49476
rect 340228 49420 352072 49476
rect 455896 49420 459004 49476
rect 459060 49420 459070 49476
rect 535602 49420 535612 49476
rect 535668 49420 538104 49476
rect 579880 49420 583212 49476
rect 583268 49420 583278 49476
rect 142034 49196 142044 49252
rect 142100 49196 144116 49252
rect 61880 48748 64316 48804
rect 64372 48748 64382 48804
rect 144060 48776 144116 49196
rect 517944 48748 519372 48804
rect 519428 48748 519438 48804
rect 530002 48748 530012 48804
rect 530068 48748 538104 48804
rect 64194 48636 64204 48692
rect 64260 48636 69692 48692
rect 69748 48636 69758 48692
rect 189522 48636 189532 48692
rect 189588 48636 199052 48692
rect 199108 48636 199118 48692
rect 19954 48188 19964 48244
rect 20020 48188 20132 48244
rect 20076 47432 20132 48188
rect 61880 48076 64092 48132
rect 64148 48076 64158 48132
rect 393960 48076 394828 48132
rect 394884 48076 394894 48132
rect 399186 48076 399196 48132
rect 399252 48076 414120 48132
rect 455410 48076 455420 48132
rect 455476 48076 455486 48132
rect 517944 48076 519260 48132
rect 519316 48076 519326 48132
rect 535154 48076 535164 48132
rect 535220 48076 538104 48132
rect 517916 47852 518252 47908
rect 518308 47852 518318 47908
rect 455868 47516 456092 47572
rect 456148 47516 456158 47572
rect 82002 47404 82012 47460
rect 82068 47404 82078 47460
rect 185864 47404 197372 47460
rect 197428 47404 197438 47460
rect 247912 47404 258188 47460
rect 258244 47404 258254 47460
rect 345202 47404 345212 47460
rect 345268 47404 352072 47460
rect 125972 47068 135212 47124
rect 135268 47068 135278 47124
rect 125972 46788 126028 47068
rect 80434 46732 80444 46788
rect 80500 46732 82040 46788
rect 123928 46732 126028 46788
rect 455868 46760 455924 47516
rect 517916 47432 517972 47852
rect 579880 47404 581308 47460
rect 581364 47404 581374 47460
rect 580402 47068 580412 47124
rect 580468 47068 580478 47124
rect 580412 46788 580468 47068
rect 579852 46732 580468 46788
rect 595560 46760 597000 46984
rect 80210 46060 80220 46116
rect 80276 46060 82040 46116
rect 123928 46060 127596 46116
rect 127652 46060 127662 46116
rect 140578 46060 140588 46116
rect 140644 46060 144088 46116
rect 185864 46060 189532 46116
rect 189588 46060 189598 46116
rect 393960 46060 396620 46116
rect 396676 46060 396686 46116
rect 535266 46060 535276 46116
rect 535332 46060 538104 46116
rect 579852 46088 579908 46732
rect 205762 45948 205772 46004
rect 205828 45948 206164 46004
rect 18274 45388 18284 45444
rect 18340 45388 20104 45444
rect 61880 45388 64204 45444
rect 64260 45388 64270 45444
rect 140914 45388 140924 45444
rect 140980 45388 144088 45444
rect 206108 45416 206164 45948
rect 247912 45388 252924 45444
rect 252980 45388 252990 45444
rect 393960 45388 396844 45444
rect 396900 45388 396910 45444
rect 535490 45388 535500 45444
rect 535556 45388 538104 45444
rect 579880 45388 583436 45444
rect 583492 45388 583502 45444
rect 61880 44716 69804 44772
rect 69860 44716 69870 44772
rect 393960 44716 396508 44772
rect 396564 44716 396574 44772
rect 472882 44716 472892 44772
rect 472948 44716 476056 44772
rect 517458 44716 517468 44772
rect 517524 44716 517534 44772
rect 579880 44716 583100 44772
rect 583156 44716 583166 44772
rect 517944 44044 519484 44100
rect 519540 44044 519550 44100
rect 517944 43372 521276 43428
rect 521332 43372 521342 43428
rect -960 36792 480 37016
rect 585442 33740 585452 33796
rect 585508 33768 595672 33796
rect 585508 33740 597000 33768
rect 595560 33544 597000 33740
rect 122658 31276 122668 31332
rect 122724 31276 264684 31332
rect 264740 31276 264750 31332
rect 61282 31164 61292 31220
rect 61348 31164 264908 31220
rect 264964 31164 264974 31220
rect 4274 31052 4284 31108
rect 4340 31052 265468 31108
rect 265524 31052 265534 31108
rect 335122 31052 335132 31108
rect 335188 31052 414092 31108
rect 414148 31052 414158 31108
rect 270022 29932 270060 29988
rect 270116 29932 270126 29988
rect 226818 29820 226828 29876
rect 226884 29820 249452 29876
rect 249508 29820 249518 29876
rect 76402 29708 76412 29764
rect 76468 29708 274316 29764
rect 274372 29708 274382 29764
rect 350242 29708 350252 29764
rect 350308 29708 372204 29764
rect 372260 29708 372270 29764
rect 12562 29596 12572 29652
rect 12628 29596 278572 29652
rect 278628 29596 278638 29652
rect 338706 29596 338716 29652
rect 338772 29596 370860 29652
rect 370916 29596 370926 29652
rect 404002 29596 404012 29652
rect 404068 29596 434812 29652
rect 434868 29596 434878 29652
rect 14242 29484 14252 29540
rect 14308 29484 282828 29540
rect 282884 29484 282894 29540
rect 351922 29484 351932 29540
rect 351988 29484 434140 29540
rect 434196 29484 434206 29540
rect 7522 29372 7532 29428
rect 7588 29372 291340 29428
rect 291396 29372 291406 29428
rect 338482 29372 338492 29428
rect 338548 29372 377580 29428
rect 377636 29372 377646 29428
rect 407362 29372 407372 29428
rect 407428 29372 498204 29428
rect 498260 29372 498270 29428
rect 230178 29260 230188 29316
rect 230244 29260 231868 29316
rect 231812 29204 231868 29260
rect 290612 29260 295596 29316
rect 295652 29260 295662 29316
rect 341842 29260 341852 29316
rect 341908 29260 436828 29316
rect 436884 29260 436894 29316
rect 461122 29260 461132 29316
rect 461188 29260 499548 29316
rect 499604 29260 499614 29316
rect 290612 29204 290668 29260
rect 231812 29148 252812 29204
rect 252868 29148 252878 29204
rect 266354 29148 266364 29204
rect 266420 29148 290668 29204
rect 19282 29036 19292 29092
rect 19348 29036 304108 29092
rect 304164 29036 304174 29092
rect 15922 28476 15932 28532
rect 15988 28476 299852 28532
rect 299908 28476 299918 28532
rect 345202 28476 345212 28532
rect 345268 28476 495516 28532
rect 495572 28476 495582 28532
rect 43586 28364 43596 28420
rect 43652 28364 63084 28420
rect 63140 28364 63150 28420
rect 78082 28364 78092 28420
rect 78148 28364 287084 28420
rect 287140 28364 287150 28420
rect 160850 28252 160860 28308
rect 160916 28252 187292 28308
rect 187348 28252 187358 28308
rect 222114 28252 222124 28308
rect 222180 28252 261212 28308
rect 261268 28252 261278 28308
rect 264562 28252 264572 28308
rect 264628 28252 308364 28308
rect 308420 28252 308430 28308
rect 231522 28140 231532 28196
rect 231588 28140 249564 28196
rect 249620 28140 249630 28196
rect 55682 26796 55692 26852
rect 55748 26796 74732 26852
rect 74788 26796 74798 26852
rect 107538 26796 107548 26852
rect 107604 26796 125132 26852
rect 125188 26796 125198 26852
rect 227490 26796 227500 26852
rect 227556 26796 247772 26852
rect 247828 26796 247838 26852
rect 336802 26796 336812 26852
rect 336868 26796 494172 26852
rect 494228 26796 494238 26852
rect 42914 26684 42924 26740
rect 42980 26684 249788 26740
rect 249844 26684 249854 26740
rect 265458 26684 265468 26740
rect 265524 26684 321132 26740
rect 321188 26684 321198 26740
rect 340162 26684 340172 26740
rect 340228 26684 492156 26740
rect 492212 26684 492222 26740
rect 39554 26572 39564 26628
rect 39620 26572 73052 26628
rect 73108 26572 73118 26628
rect 103506 26572 103516 26628
rect 103572 26572 262892 26628
rect 262948 26572 262958 26628
rect 263106 26572 263116 26628
rect 263172 26572 316876 26628
rect 316932 26572 316942 26628
rect 352034 26572 352044 26628
rect 352100 26572 432796 26628
rect 432852 26572 432862 26628
rect 464482 26572 464492 26628
rect 464548 26572 562268 26628
rect 562324 26572 562334 26628
rect 38882 26460 38892 26516
rect 38948 26460 62972 26516
rect 63028 26460 63038 26516
rect 89394 26460 89404 26516
rect 89460 26460 204092 26516
rect 204148 26460 204158 26516
rect 205762 26460 205772 26516
rect 205828 26460 312620 26516
rect 312676 26460 312686 26516
rect 337026 26460 337036 26516
rect 337092 26460 376908 26516
rect 376964 26460 376974 26516
rect 414082 26460 414092 26516
rect 414148 26460 438844 26516
rect 438900 26460 438910 26516
rect 40226 26348 40236 26404
rect 40292 26348 61292 26404
rect 61348 26348 61358 26404
rect 104178 26348 104188 26404
rect 104244 26348 122668 26404
rect 122724 26348 122734 26404
rect 169586 26348 169596 26404
rect 169652 26348 259532 26404
rect 259588 26348 259598 26404
rect 348562 26348 348572 26404
rect 348628 26348 374892 26404
rect 374948 26348 374958 26404
rect 167570 26236 167580 26292
rect 167636 26236 256172 26292
rect 256228 26236 256238 26292
rect 10882 26124 10892 26180
rect 10948 26124 325388 26180
rect 325444 26124 325454 26180
rect 4162 24332 4172 24388
rect 4228 24332 329644 24388
rect 329700 24332 329710 24388
rect 392 22904 4172 22932
rect -960 22876 4172 22904
rect 4228 22876 4238 22932
rect -960 22680 480 22876
rect 595560 20328 597000 20552
rect -960 8596 480 8792
rect -960 8568 200844 8596
rect 392 8540 200844 8568
rect 200900 8540 200910 8596
rect 595560 7112 597000 7336
rect 11554 5068 11564 5124
rect 11620 5068 18396 5124
rect 18452 5068 18462 5124
<< via3 >>
rect 319116 571228 319172 571284
rect 330764 571228 330820 571284
rect 317996 569996 318052 570052
rect 290444 569772 290500 569828
rect 303660 569548 303716 569604
rect 315756 569548 315812 569604
rect 317996 569324 318052 569380
rect 270284 568876 270340 568932
rect 271404 568876 271460 568932
rect 272524 568876 272580 568932
rect 289324 568876 289380 568932
rect 300524 568876 300580 568932
rect 301644 568876 301700 568932
rect 302764 568876 302820 568932
rect 302764 568652 302820 568708
rect 270284 567756 270340 567812
rect 300524 567644 300580 567700
rect 272524 567532 272580 567588
rect 303660 567420 303716 567476
rect 301644 567308 301700 567364
rect 315756 567196 315812 567252
rect 319116 567084 319172 567140
rect 271404 566972 271460 567028
rect 141036 563948 141092 564004
rect 583212 563948 583268 564004
rect 141036 556108 141092 556164
rect 141932 556108 141988 556164
rect 18396 555884 18452 555940
rect 141036 555884 141092 555940
rect 80108 555212 80164 555268
rect 144060 555212 144116 555268
rect 352716 555212 352772 555268
rect 473676 555212 473732 555268
rect 414652 555100 414708 555156
rect 80444 554540 80500 554596
rect 126924 554540 126980 554596
rect 201628 554540 201684 554596
rect 476028 554764 476084 554820
rect 18396 554428 18452 554484
rect 82684 553868 82740 553924
rect 252812 553868 252868 553924
rect 347788 553868 347844 553924
rect 410956 553868 411012 553924
rect 473452 553868 473508 553924
rect 519036 553868 519092 553924
rect 18284 553196 18340 553252
rect 340284 553196 340340 553252
rect 410732 553196 410788 553252
rect 458780 553196 458836 553252
rect 472892 553196 472948 553252
rect 583436 553196 583492 553252
rect 65100 552524 65156 552580
rect 127260 552524 127316 552580
rect 204876 552524 204932 552580
rect 261324 552524 261380 552580
rect 473228 552524 473284 552580
rect 535500 552524 535556 552580
rect 583324 552524 583380 552580
rect 18396 551852 18452 551908
rect 141036 551852 141092 551908
rect 203196 551852 203252 551908
rect 396844 551852 396900 551908
rect 458668 551852 458724 551908
rect 521276 551852 521332 551908
rect 341964 551628 342020 551684
rect 347788 551628 347844 551684
rect 80332 551180 80388 551236
rect 140924 551180 140980 551236
rect 189084 551180 189140 551236
rect 262892 551180 262948 551236
rect 348572 551180 348628 551236
rect 394828 551180 394884 551236
rect 459004 551180 459060 551236
rect 535276 551180 535332 551236
rect 579628 551180 579684 551236
rect 518252 551068 518308 551124
rect 582428 551068 582484 551124
rect 345212 550508 345268 550564
rect 473116 550508 473172 550564
rect 205772 549948 205828 550004
rect 74732 549836 74788 549892
rect 188972 549836 189028 549892
rect 348684 549836 348740 549892
rect 410844 549836 410900 549892
rect 520940 549836 520996 549892
rect 534268 549836 534324 549892
rect 74844 549164 74900 549220
rect 82012 549164 82068 549220
rect 338492 549164 338548 549220
rect 458892 549164 458948 549220
rect 64652 548492 64708 548548
rect 143612 548492 143668 548548
rect 189196 548492 189252 548548
rect 257852 548492 257908 548548
rect 402332 548492 402388 548548
rect 456988 548492 457044 548548
rect 461132 548492 461188 548548
rect 473228 548492 473284 548548
rect 523292 548492 523348 548548
rect 534268 548492 534324 548548
rect 583100 548492 583156 548548
rect 126812 547820 126868 547876
rect 264572 547820 264628 547876
rect 473228 547820 473284 547876
rect 535164 547820 535220 547876
rect 456092 547708 456148 547764
rect 458668 547708 458724 547764
rect 82236 547148 82292 547204
rect 127036 547148 127092 547204
rect 251916 547148 251972 547204
rect 393372 547148 393428 547204
rect 521052 547148 521108 547204
rect 535052 547148 535108 547204
rect 82124 546476 82180 546532
rect 142044 546476 142100 546532
rect 411068 546476 411124 546532
rect 458668 546476 458724 546532
rect 473004 546476 473060 546532
rect 519260 546476 519316 546532
rect 581308 546476 581364 546532
rect 141036 546028 141092 546084
rect 143724 546028 143780 546084
rect 457772 546028 457828 546084
rect 458780 546028 458836 546084
rect 20076 545804 20132 545860
rect 64764 545804 64820 545860
rect 127148 545804 127204 545860
rect 197372 545804 197428 545860
rect 254492 545804 254548 545860
rect 473340 545804 473396 545860
rect 18172 545132 18228 545188
rect 138572 545132 138628 545188
rect 140812 545132 140868 545188
rect 189420 545132 189476 545188
rect 259980 545132 260036 545188
rect 341852 545132 341908 545188
rect 458780 545132 458836 545188
rect 581420 545804 581476 545860
rect 519932 544796 519988 544852
rect 64988 544460 65044 544516
rect 80220 544460 80276 544516
rect 141036 544460 141092 544516
rect 203084 544460 203140 544516
rect 256284 544460 256340 544516
rect 394940 544460 394996 544516
rect 519148 544460 519204 544516
rect 203196 544348 203252 544404
rect 204092 544348 204148 544404
rect 18060 543788 18116 543844
rect 203084 543788 203140 543844
rect 261212 543788 261268 543844
rect 340172 543788 340228 543844
rect 398972 543788 399028 543844
rect 535388 543788 535444 543844
rect 395612 543228 395668 543284
rect 142716 543116 142772 543172
rect 520828 543116 520884 543172
rect 396732 542668 396788 542724
rect 396620 542444 396676 542500
rect 455308 542444 455364 542500
rect 521164 541772 521220 541828
rect 64876 538412 64932 538468
rect 464492 536732 464548 536788
rect 473452 536732 473508 536788
rect 252812 533372 252868 533428
rect 263900 533372 263956 533428
rect 519036 533372 519092 533428
rect 535388 533372 535444 533428
rect 254492 531580 254548 531636
rect 263788 531020 263844 531076
rect 523292 530460 523348 530516
rect 140812 530236 140868 530292
rect 205996 530236 206052 530292
rect 65100 530124 65156 530180
rect 259532 530124 259588 530180
rect 456876 530124 456932 530180
rect 583212 530124 583268 530180
rect 18172 530012 18228 530068
rect 256172 530012 256228 530068
rect 205772 529900 205828 529956
rect 582428 529900 582484 529956
rect 263900 529340 263956 529396
rect 140924 529116 140980 529172
rect 146076 529116 146132 529172
rect 261324 528780 261380 528836
rect 332668 528332 332724 528388
rect 18060 528220 18116 528276
rect 261548 528220 261604 528276
rect 80220 527996 80276 528052
rect 252812 527996 252868 528052
rect 519036 528220 519092 528276
rect 354396 527996 354452 528052
rect 535500 527996 535556 528052
rect 357756 527884 357812 527940
rect 520828 527884 520884 527940
rect 332668 527772 332724 527828
rect 127260 526652 127316 526708
rect 249452 526652 249508 526708
rect 259980 526540 260036 526596
rect 456876 526540 456932 526596
rect 354396 525980 354452 526036
rect 256284 524860 256340 524916
rect 251916 524300 251972 524356
rect 521164 523740 521220 523796
rect 203084 523516 203140 523572
rect 246092 523516 246148 523572
rect 348796 523292 348852 523348
rect 473340 523292 473396 523348
rect 146076 523180 146132 523236
rect 197372 522620 197428 522676
rect 518252 522620 518308 522676
rect 189196 522060 189252 522116
rect 357756 522060 357812 522116
rect 351932 521948 351988 522004
rect 396732 521948 396788 522004
rect 126924 521724 126980 521780
rect 256508 521724 256564 521780
rect 18284 521612 18340 521668
rect 256284 521612 256340 521668
rect 189420 521500 189476 521556
rect 205996 520940 206052 520996
rect 142716 520380 142772 520436
rect 355292 520156 355348 520212
rect 411068 520156 411124 520212
rect 80444 520044 80500 520100
rect 247772 520044 247828 520100
rect 380492 520044 380548 520100
rect 459004 520044 459060 520100
rect 82236 519932 82292 519988
rect 263788 519932 263844 519988
rect 336812 519932 336868 519988
rect 521052 519932 521108 519988
rect 143724 519820 143780 519876
rect 519260 519260 519316 519316
rect 461132 518700 461188 518756
rect 82124 518364 82180 518420
rect 264908 518364 264964 518420
rect 80332 518252 80388 518308
rect 263116 518252 263172 518308
rect 353612 518252 353668 518308
rect 583324 518252 583380 518308
rect 519932 518140 519988 518196
rect 464492 517020 464548 517076
rect 353724 516684 353780 516740
rect 535276 516684 535332 516740
rect 335244 516572 335300 516628
rect 519148 516572 519204 516628
rect 141932 516460 141988 516516
rect 82012 515900 82068 515956
rect 398972 515900 399028 515956
rect 80108 514892 80164 514948
rect 257964 514892 258020 514948
rect 142044 514780 142100 514836
rect 456988 514780 457044 514836
rect 263788 514220 263844 514276
rect 127036 513660 127092 513716
rect 380492 513660 380548 513716
rect 342076 513324 342132 513380
rect 473228 513324 473284 513380
rect 345548 513212 345604 513268
rect 583100 513212 583156 513268
rect 126812 513100 126868 513156
rect 456092 513100 456148 513156
rect 264908 512540 264964 512596
rect 457772 512540 457828 512596
rect 355292 511980 355348 512036
rect 334460 511868 334516 511924
rect 402332 511868 402388 511924
rect 141036 511644 141092 511700
rect 247884 511644 247940 511700
rect 354396 511644 354452 511700
rect 458892 511644 458948 511700
rect 340396 511532 340452 511588
rect 520940 511532 520996 511588
rect 127148 510860 127204 510916
rect 354396 510300 354452 510356
rect 334348 510188 334404 510244
rect 394828 510188 394884 510244
rect 335468 510076 335524 510132
rect 455308 510076 455364 510132
rect 345324 509964 345380 510020
rect 473116 509964 473172 510020
rect 74844 509852 74900 509908
rect 263788 509852 263844 509908
rect 353836 509852 353892 509908
rect 535164 509852 535220 509908
rect 334460 509740 334516 509796
rect 138572 509180 138628 509236
rect 143612 508620 143668 508676
rect 342188 508284 342244 508340
rect 410844 508284 410900 508340
rect 263788 508060 263844 508116
rect 341964 508060 342020 508116
rect 261548 507500 261604 507556
rect 334348 507500 334404 507556
rect 350588 506828 350644 506884
rect 410956 506828 411012 506884
rect 189084 506716 189140 506772
rect 247996 506716 248052 506772
rect 352156 506716 352212 506772
rect 458668 506716 458724 506772
rect 335132 506604 335188 506660
rect 393372 506604 393428 506660
rect 402332 506604 402388 506660
rect 535052 506604 535108 506660
rect 338716 506492 338772 506548
rect 521276 506492 521332 506548
rect 64652 506380 64708 506436
rect 337708 505372 337764 505428
rect 396620 505372 396676 505428
rect 64764 505260 64820 505316
rect 348908 505148 348964 505204
rect 410732 505148 410788 505204
rect 338604 505036 338660 505092
rect 458780 505036 458836 505092
rect 352268 504924 352324 504980
rect 473004 504924 473060 504980
rect 74732 504812 74788 504868
rect 264684 504812 264740 504868
rect 335356 504812 335412 504868
rect 394940 504812 394996 504868
rect 64988 504700 65044 504756
rect 340284 504700 340340 504756
rect 18396 504140 18452 504196
rect 338492 503580 338548 503636
rect 335916 503468 335972 503524
rect 348684 503468 348740 503524
rect 349020 503468 349076 503524
rect 396844 503468 396900 503524
rect 188972 503244 189028 503300
rect 251916 503244 251972 503300
rect 393932 503132 393988 503188
rect 583436 503132 583492 503188
rect 395612 503020 395668 503076
rect 64876 502460 64932 502516
rect 20076 501900 20132 501956
rect 335916 501900 335972 501956
rect 203196 501452 203252 501508
rect 246876 501452 246932 501508
rect 344092 501452 344148 501508
rect 472892 501452 472948 501508
rect 337708 501340 337764 501396
rect 257852 500220 257908 500276
rect 581420 500220 581476 500276
rect 262892 500108 262948 500164
rect 263900 500108 263956 500164
rect 264572 499660 264628 499716
rect 353836 499660 353892 499716
rect 261212 499100 261268 499156
rect 345548 499100 345604 499156
rect 581308 498540 581364 498596
rect 263900 497980 263956 498036
rect 579628 497980 579684 498036
rect 246876 497532 246932 497588
rect 353724 497420 353780 497476
rect 204092 496860 204148 496916
rect 402332 496860 402388 496916
rect 393932 495740 393988 495796
rect 246092 495180 246148 495236
rect 353612 494956 353668 495012
rect 348796 493500 348852 493556
rect 143612 493388 143668 493444
rect 459228 493388 459284 493444
rect 247884 492940 247940 492996
rect 336812 492940 336868 492996
rect 69692 492716 69748 492772
rect 140924 492716 140980 492772
rect 345324 491820 345380 491876
rect 352268 491260 352324 491316
rect 247996 490700 248052 490756
rect 342076 490140 342132 490196
rect 344092 489580 344148 489636
rect 335244 488460 335300 488516
rect 335580 488012 335636 488068
rect 345212 488012 345268 488068
rect 340396 487900 340452 487956
rect 251916 487340 251972 487396
rect 338716 487340 338772 487396
rect 247772 486780 247828 486836
rect 257964 486220 258020 486276
rect 348908 485660 348964 485716
rect 256508 485100 256564 485156
rect 534268 484652 534324 484708
rect 249452 484540 249508 484596
rect 350588 484540 350644 484596
rect 476028 484316 476084 484372
rect 18396 483980 18452 484036
rect 20076 483980 20132 484036
rect 342188 483980 342244 484036
rect 473676 483980 473732 484036
rect 141036 483756 141092 483812
rect 335804 483756 335860 483812
rect 340172 483756 340228 483812
rect 252812 483420 252868 483476
rect 335468 483420 335524 483476
rect 64764 483308 64820 483364
rect 82684 483308 82740 483364
rect 201628 483308 201684 483364
rect 352716 483308 352772 483364
rect 396844 483308 396900 483364
rect 458668 483308 458724 483364
rect 519148 483308 519204 483364
rect 189084 482636 189140 482692
rect 259644 482636 259700 482692
rect 396732 482636 396788 482692
rect 410844 482636 410900 482692
rect 458780 482636 458836 482692
rect 472108 482636 472164 482692
rect 206668 482300 206724 482356
rect 136892 482076 136948 482132
rect 82236 481964 82292 482020
rect 127596 481964 127652 482020
rect 262892 481964 262948 482020
rect 411180 481964 411236 482020
rect 456988 481964 457044 482020
rect 472220 481964 472276 482020
rect 581308 482636 581364 482692
rect 534268 481964 534324 482020
rect 518252 481852 518308 481908
rect 263116 481740 263172 481796
rect 352156 481740 352212 481796
rect 461132 481404 461188 481460
rect 472108 481404 472164 481460
rect 64876 481292 64932 481348
rect 142044 481292 142100 481348
rect 203196 481292 203252 481348
rect 410956 481292 411012 481348
rect 459004 481292 459060 481348
rect 462812 481292 462868 481348
rect 535052 481292 535108 481348
rect 338604 481180 338660 481236
rect 414652 481068 414708 481124
rect 18172 480620 18228 480676
rect 141036 480620 141092 480676
rect 261324 480620 261380 480676
rect 458892 480620 458948 480676
rect 583324 480620 583380 480676
rect 127596 480396 127652 480452
rect 130172 480396 130228 480452
rect 140924 480396 140980 480452
rect 143724 480396 143780 480452
rect 349020 480060 349076 480116
rect 18284 479948 18340 480004
rect 133532 479948 133588 480004
rect 197372 479948 197428 480004
rect 348796 479948 348852 480004
rect 394828 479948 394884 480004
rect 455308 479948 455364 480004
rect 472892 479948 472948 480004
rect 517468 479948 517524 480004
rect 523292 479612 523348 479668
rect 534268 479612 534324 479668
rect 259532 479500 259588 479556
rect 348572 479500 348628 479556
rect 65100 479276 65156 479332
rect 80556 479276 80612 479332
rect 204204 479276 204260 479332
rect 348684 479276 348740 479332
rect 394940 479276 394996 479332
rect 455420 479276 455476 479332
rect 473116 479276 473172 479332
rect 521164 479276 521220 479332
rect 581420 479276 581476 479332
rect 264684 478940 264740 478996
rect 73164 478604 73220 478660
rect 80332 478604 80388 478660
rect 127596 478604 127652 478660
rect 188972 478604 189028 478660
rect 206556 478604 206612 478660
rect 251020 478604 251076 478660
rect 342076 478604 342132 478660
rect 396508 478604 396564 478660
rect 459116 478604 459172 478660
rect 582988 478604 583044 478660
rect 341852 478380 341908 478436
rect 579628 478380 579684 478436
rect 194908 477932 194964 477988
rect 250908 477932 250964 477988
rect 404012 477932 404068 477988
rect 457324 477932 457380 477988
rect 467852 477932 467908 477988
rect 256172 477820 256228 477876
rect 17948 477260 18004 477316
rect 140924 477260 140980 477316
rect 252812 477260 252868 477316
rect 335356 477260 335412 477316
rect 518476 477148 518532 477204
rect 78316 476588 78372 476644
rect 80444 476588 80500 476644
rect 135212 476588 135268 476644
rect 140812 476588 140868 476644
rect 259532 476588 259588 476644
rect 340172 476588 340228 476644
rect 396620 476588 396676 476644
rect 519260 476588 519316 476644
rect 127596 476252 127652 476308
rect 138572 476252 138628 476308
rect 251020 476252 251076 476308
rect 264572 476252 264628 476308
rect 335132 476140 335188 476196
rect 18060 475916 18116 475972
rect 64652 475916 64708 475972
rect 189532 475916 189588 475972
rect 261212 475916 261268 475972
rect 393372 475916 393428 475972
rect 400652 475916 400708 475972
rect 455532 475916 455588 475972
rect 520940 475916 520996 475972
rect 579404 475916 579460 475972
rect 141036 475468 141092 475524
rect 141932 475468 141988 475524
rect 335356 475468 335412 475524
rect 339388 475468 339444 475524
rect 457772 475468 457828 475524
rect 458668 475468 458724 475524
rect 395612 475356 395668 475412
rect 396844 475356 396900 475412
rect 20076 475244 20132 475300
rect 256284 475020 256340 475076
rect 351932 475020 351988 475076
rect 250908 474796 250964 474852
rect 256508 474796 256564 474852
rect 126812 474572 126868 474628
rect 335580 474460 335636 474516
rect 535164 474572 535220 474628
rect 579628 474572 579684 474628
rect 456092 474460 456148 474516
rect 457212 474012 457268 474068
rect 82124 473900 82180 473956
rect 127036 473900 127092 473956
rect 189532 473900 189588 473956
rect 262108 473900 262164 473956
rect 335804 473900 335860 473956
rect 348572 473900 348628 473956
rect 402332 473900 402388 473956
rect 457100 473900 457156 473956
rect 521052 473900 521108 473956
rect 345212 473788 345268 473844
rect 348684 473788 348740 473844
rect 263788 473340 263844 473396
rect 334460 473340 334516 473396
rect 69804 473228 69860 473284
rect 199052 473228 199108 473284
rect 257852 473228 257908 473284
rect 396844 473228 396900 473284
rect 410732 473228 410788 473284
rect 73052 472556 73108 472612
rect 395052 471884 395108 471940
rect 247996 471660 248052 471716
rect 351036 471660 351092 471716
rect 64988 471212 65044 471268
rect 144396 471212 144452 471268
rect 334348 471100 334404 471156
rect 334460 470540 334516 470596
rect 262108 469980 262164 470036
rect 579292 469868 579348 469924
rect 334460 468860 334516 468916
rect 189084 467852 189140 467908
rect 204092 467852 204148 467908
rect 261324 467740 261380 467796
rect 249452 466172 249508 466228
rect 263900 466172 263956 466228
rect 259532 466060 259588 466116
rect 81452 465164 81508 465220
rect 263788 464940 263844 464996
rect 334460 464380 334516 464436
rect 264684 463820 264740 463876
rect 263900 463260 263956 463316
rect 398972 462812 399028 462868
rect 410844 462812 410900 462868
rect 263788 462700 263844 462756
rect 249564 462140 249620 462196
rect 264012 461580 264068 461636
rect 82012 461132 82068 461188
rect 142156 461132 142212 461188
rect 188972 461132 189028 461188
rect 205772 461132 205828 461188
rect 334460 461020 334516 461076
rect 264124 460460 264180 460516
rect 334348 460460 334404 460516
rect 335356 459900 335412 459956
rect 518252 459340 518308 459396
rect 143724 459116 143780 459172
rect 204204 458780 204260 458836
rect 518476 458780 518532 458836
rect 230860 458108 230916 458164
rect 354396 458108 354452 458164
rect 459116 458108 459172 458164
rect 160860 457996 160916 458052
rect 336028 457996 336084 458052
rect 459004 457996 459060 458052
rect 142044 457884 142100 457940
rect 263900 457884 263956 457940
rect 493724 457884 493780 457940
rect 69692 457772 69748 457828
rect 264684 457772 264740 457828
rect 130172 457660 130228 457716
rect 133532 456988 133588 457044
rect 392476 457100 392532 457156
rect 396732 457100 396788 457156
rect 493724 457100 493780 457156
rect 457324 456988 457380 457044
rect 160860 456876 160916 456932
rect 230860 456876 230916 456932
rect 354396 456652 354452 456708
rect 336140 456316 336196 456372
rect 411180 456316 411236 456372
rect 354396 456204 354452 456260
rect 459228 456204 459284 456260
rect 82012 456092 82068 456148
rect 263788 456092 263844 456148
rect 337708 456092 337764 456148
rect 458892 456092 458948 456148
rect 135212 455980 135268 456036
rect 136892 455420 136948 455476
rect 455532 455420 455588 455476
rect 457212 454860 457268 454916
rect 138572 454300 138628 454356
rect 456092 454300 456148 454356
rect 263900 453740 263956 453796
rect 337708 453740 337764 453796
rect 80332 452844 80388 452900
rect 258188 452844 258244 452900
rect 263788 452620 263844 452676
rect 336140 452620 336196 452676
rect 336028 452060 336084 452116
rect 82124 451500 82180 451556
rect 457772 451500 457828 451556
rect 335132 451164 335188 451220
rect 393372 451164 393428 451220
rect 20076 451052 20132 451108
rect 264908 451052 264964 451108
rect 142156 450940 142212 450996
rect 398972 450940 399028 450996
rect 143612 450380 143668 450436
rect 354396 450380 354452 450436
rect 345212 449820 345268 449876
rect 351932 449708 351988 449764
rect 396620 449708 396676 449764
rect 342188 449596 342244 449652
rect 396844 449596 396900 449652
rect 392364 449484 392420 449540
rect 535052 449484 535108 449540
rect 17948 449372 18004 449428
rect 247772 449372 247828 449428
rect 352156 449372 352212 449428
rect 520940 449372 520996 449428
rect 64764 449260 64820 449316
rect 395052 449260 395108 449316
rect 65100 448700 65156 448756
rect 18172 448140 18228 448196
rect 336812 447804 336868 447860
rect 458780 447804 458836 447860
rect 355292 447692 355348 447748
rect 535164 447692 535220 447748
rect 64876 447580 64932 447636
rect 392476 447580 392532 447636
rect 395612 447020 395668 447076
rect 344428 446572 344484 446628
rect 396508 446572 396564 446628
rect 73164 446460 73220 446516
rect 353612 446348 353668 446404
rect 410732 446348 410788 446404
rect 342300 446236 342356 446292
rect 410956 446236 411012 446292
rect 370412 446124 370468 446180
rect 521164 446124 521220 446180
rect 127036 446012 127092 446068
rect 261324 446012 261380 446068
rect 335804 446012 335860 446068
rect 348796 446012 348852 446068
rect 391356 446012 391412 446068
rect 583324 446012 583380 446068
rect 78316 445900 78372 445956
rect 18060 444780 18116 444836
rect 344428 444780 344484 444836
rect 335916 444668 335972 444724
rect 394940 444668 394996 444724
rect 338492 444556 338548 444612
rect 472892 444556 472948 444612
rect 140812 444444 140868 444500
rect 253148 444444 253204 444500
rect 81452 444220 81508 444276
rect 342076 444220 342132 444276
rect 264908 443100 264964 443156
rect 335916 443100 335972 443156
rect 264684 442540 264740 442596
rect 335804 442540 335860 442596
rect 203196 441980 203252 442036
rect 261212 441868 261268 441924
rect 581308 441420 581364 441476
rect 64988 441084 65044 441140
rect 256172 441084 256228 441140
rect 64652 440972 64708 441028
rect 259532 440972 259588 441028
rect 256508 440860 256564 440916
rect 391356 440300 391412 440356
rect 252812 439740 252868 439796
rect 392364 439740 392420 439796
rect 69804 439516 69860 439572
rect 264684 439516 264740 439572
rect 257852 439180 257908 439236
rect 581420 439180 581476 439236
rect 259644 438060 259700 438116
rect 523292 438060 523348 438116
rect 126812 437948 126868 438004
rect 247884 437948 247940 438004
rect 18284 437612 18340 437668
rect 261212 437612 261268 437668
rect 335356 437612 335412 437668
rect 394828 437612 394884 437668
rect 262892 437500 262948 437556
rect 264572 436380 264628 436436
rect 355292 435820 355348 435876
rect 205772 434700 205828 434756
rect 80556 434364 80612 434420
rect 263340 434364 263396 434420
rect 73052 434252 73108 434308
rect 264572 434252 264628 434308
rect 204092 433580 204148 433636
rect 519260 433580 519316 433636
rect 141932 433020 141988 433076
rect 519148 433020 519204 433076
rect 80444 432572 80500 432628
rect 255612 432572 255668 432628
rect 335804 432572 335860 432628
rect 455420 432572 455476 432628
rect 517468 432460 517524 432516
rect 467852 431900 467908 431956
rect 461132 430780 461188 430836
rect 352156 430556 352212 430612
rect 370412 429660 370468 429716
rect 253148 429100 253204 429156
rect 338492 429100 338548 429156
rect 255612 428540 255668 428596
rect 404012 428540 404068 428596
rect 402332 427980 402388 428036
rect 334460 427532 334516 427588
rect 455308 427532 455364 427588
rect 457100 427420 457156 427476
rect 436828 426972 436884 427028
rect 438172 426972 438228 427028
rect 335804 426860 335860 426916
rect 173852 426636 173908 426692
rect 400652 426636 400708 426692
rect 82236 426524 82292 426580
rect 170268 426412 170324 426468
rect 222796 426412 222852 426468
rect 232204 426412 232260 426468
rect 173740 426300 173796 426356
rect 436828 426188 436884 426244
rect 438172 426188 438228 426244
rect 170268 426076 170324 426132
rect 173852 426076 173908 426132
rect 222796 426076 222852 426132
rect 232204 425964 232260 426020
rect 173740 425852 173796 425908
rect 263340 425740 263396 425796
rect 353612 425740 353668 425796
rect 258188 425180 258244 425236
rect 342300 425180 342356 425236
rect 456988 424620 457044 424676
rect 247884 424060 247940 424116
rect 336812 424060 336868 424116
rect 261324 423500 261380 423556
rect 334460 423500 334516 423556
rect 348796 421484 348852 421540
rect 396620 421484 396676 421540
rect 410732 421484 410788 421540
rect 472108 421484 472164 421540
rect 348572 421260 348628 421316
rect 259532 420700 259588 420756
rect 335132 420700 335188 420756
rect 261212 420140 261268 420196
rect 340172 420140 340228 420196
rect 395612 419916 395668 419972
rect 247772 419580 247828 419636
rect 342188 419580 342244 419636
rect 256172 419020 256228 419076
rect 335356 419020 335412 419076
rect 264572 418460 264628 418516
rect 264684 416220 264740 416276
rect 351932 416220 351988 416276
rect 263900 415100 263956 415156
rect 334460 415100 334516 415156
rect 206668 414988 206724 415044
rect 334460 414540 334516 414596
rect 262892 413980 262948 414036
rect 263340 413420 263396 413476
rect 334460 413420 334516 413476
rect 472108 413420 472164 413476
rect 263788 412860 263844 412916
rect 351036 412860 351092 412916
rect 82684 412748 82740 412804
rect 141036 412748 141092 412804
rect 144060 412748 144116 412804
rect 334348 412300 334404 412356
rect 18396 411740 18452 411796
rect 201628 412076 201684 412132
rect 262108 412076 262164 412132
rect 472108 412076 472164 412132
rect 334460 411740 334516 411796
rect 19964 411628 20020 411684
rect 18060 411404 18116 411460
rect 135212 411404 135268 411460
rect 352716 411404 352772 411460
rect 411516 411404 411572 411460
rect 414652 411404 414708 411460
rect 464492 411404 464548 411460
rect 534380 411404 534436 411460
rect 334460 411180 334516 411236
rect 19852 410732 19908 410788
rect 69692 410732 69748 410788
rect 127036 410732 127092 410788
rect 457324 410732 457380 410788
rect 473116 410732 473172 410788
rect 530012 410732 530068 410788
rect 579292 410732 579348 410788
rect 262108 410620 262164 410676
rect 579628 410620 579684 410676
rect 263900 410172 263956 410228
rect 19740 410060 19796 410116
rect 74732 410060 74788 410116
rect 82684 410060 82740 410116
rect 126812 410060 126868 410116
rect 142716 410060 142772 410116
rect 334348 410060 334404 410116
rect 338604 410060 338660 410116
rect 394828 410060 394884 410116
rect 402332 410060 402388 410116
rect 144284 409836 144340 409892
rect 79772 409388 79828 409444
rect 126252 409388 126308 409444
rect 334460 409500 334516 409556
rect 521052 410060 521108 410116
rect 534268 410060 534324 410116
rect 203196 409388 203252 409444
rect 347788 409388 347844 409444
rect 456092 409388 456148 409444
rect 533372 409388 533428 409444
rect 579292 409388 579348 409444
rect 334348 409052 334404 409108
rect 350364 409052 350420 409108
rect 260316 408940 260372 408996
rect 127260 408716 127316 408772
rect 206108 408716 206164 408772
rect 458892 408716 458948 408772
rect 467852 408716 467908 408772
rect 144284 408380 144340 408436
rect 18284 408044 18340 408100
rect 76412 407372 76468 407428
rect 188972 408044 189028 408100
rect 204876 408044 204932 408100
rect 263340 408044 263396 408100
rect 338492 408044 338548 408100
rect 394940 408044 394996 408100
rect 458780 408044 458836 408100
rect 519148 408044 519204 408100
rect 535052 408044 535108 408100
rect 334460 407820 334516 407876
rect 199836 407372 199892 407428
rect 256172 407372 256228 407428
rect 411180 407372 411236 407428
rect 455532 407372 455588 407428
rect 581308 407372 581364 407428
rect 82348 407260 82404 407316
rect 144396 407260 144452 407316
rect 263788 407260 263844 407316
rect 20636 406700 20692 406756
rect 81452 406700 81508 406756
rect 136108 406700 136164 406756
rect 259532 406700 259588 406756
rect 260316 406700 260372 406756
rect 411068 406700 411124 406756
rect 457100 406700 457156 406756
rect 579628 406700 579684 406756
rect 144284 406588 144340 406644
rect 579852 406476 579908 406532
rect 262108 406140 262164 406196
rect 64652 406028 64708 406084
rect 127148 406028 127204 406084
rect 191548 406028 191604 406084
rect 253148 406028 253204 406084
rect 341852 406028 341908 406084
rect 395052 406028 395108 406084
rect 406588 406028 406644 406084
rect 458668 406028 458724 406084
rect 472892 406028 472948 406084
rect 336028 405580 336084 405636
rect 73052 405356 73108 405412
rect 204988 405356 205044 405412
rect 456988 405356 457044 405412
rect 583100 405356 583156 405412
rect 519932 405244 519988 405300
rect 263900 405020 263956 405076
rect 81564 404684 81620 404740
rect 189420 404684 189476 404740
rect 396508 404684 396564 404740
rect 411180 404684 411236 404740
rect 459004 404684 459060 404740
rect 263788 404460 263844 404516
rect 126924 404012 126980 404068
rect 189532 404012 189588 404068
rect 457212 404012 457268 404068
rect 461132 404012 461188 404068
rect 473116 404012 473172 404068
rect 263452 403900 263508 403956
rect 334460 403900 334516 403956
rect 252812 403452 252868 403508
rect 141036 403340 141092 403396
rect 189308 403340 189364 403396
rect 262892 403340 262948 403396
rect 396732 403340 396788 403396
rect 455308 403340 455364 403396
rect 472108 403340 472164 403396
rect 340508 403228 340564 403284
rect 347788 403228 347844 403284
rect 579740 403116 579796 403172
rect 263788 402780 263844 402836
rect 334460 402780 334516 402836
rect 20076 402668 20132 402724
rect 143612 402668 143668 402724
rect 259644 402668 259700 402724
rect 345212 402668 345268 402724
rect 401212 402668 401268 402724
rect 455420 402668 455476 402724
rect 520940 402668 520996 402724
rect 579628 402556 579684 402612
rect 398972 402332 399028 402388
rect 411180 402332 411236 402388
rect 189532 401996 189588 402052
rect 204764 401996 204820 402052
rect 411180 401996 411236 402052
rect 461132 401996 461188 402052
rect 517468 401996 517524 402052
rect 534268 401996 534324 402052
rect 263900 401660 263956 401716
rect 350252 401660 350308 401716
rect 18172 401324 18228 401380
rect 64876 401324 64932 401380
rect 133532 401324 133588 401380
rect 192332 401324 192388 401380
rect 517244 401324 517300 401380
rect 334348 401100 334404 401156
rect 82348 400652 82404 400708
rect 535612 400652 535668 400708
rect 262108 400540 262164 400596
rect 262220 399980 262276 400036
rect 336252 399420 336308 399476
rect 336812 398972 336868 399028
rect 348796 398972 348852 399028
rect 334460 398860 334516 398916
rect 533484 398524 533540 398580
rect 535612 398524 535668 398580
rect 263788 398300 263844 398356
rect 351036 398300 351092 398356
rect 263788 397740 263844 397796
rect 334460 397180 334516 397236
rect 249452 396620 249508 396676
rect 334348 396620 334404 396676
rect 334460 396060 334516 396116
rect 188972 395612 189028 395668
rect 205772 395612 205828 395668
rect 263788 395500 263844 395556
rect 334348 395500 334404 395556
rect 74844 395276 74900 395332
rect 263900 394940 263956 394996
rect 334460 394380 334516 394436
rect 334348 393820 334404 393876
rect 263788 392700 263844 392756
rect 334348 392700 334404 392756
rect 334460 392140 334516 392196
rect 263788 391020 263844 391076
rect 579628 391020 579684 391076
rect 263900 390460 263956 390516
rect 455532 390460 455588 390516
rect 263788 389900 263844 389956
rect 253148 388892 253204 388948
rect 265020 388892 265076 388948
rect 340508 388220 340564 388276
rect 20076 387996 20132 388052
rect 263900 387996 263956 388052
rect 81564 387884 81620 387940
rect 263788 387884 263844 387940
rect 74732 387660 74788 387716
rect 338604 387660 338660 387716
rect 349468 387660 349524 387716
rect 396620 387660 396676 387716
rect 347788 387212 347844 387268
rect 583100 387212 583156 387268
rect 73052 387100 73108 387156
rect 19852 386540 19908 386596
rect 336812 386540 336868 386596
rect 259532 386316 259588 386372
rect 263788 386316 263844 386372
rect 503132 385756 503188 385812
rect 520940 385756 520996 385812
rect 371308 385644 371364 385700
rect 535052 385644 535108 385700
rect 395612 385532 395668 385588
rect 400652 385532 400708 385588
rect 472892 385532 472948 385588
rect 476252 385532 476308 385588
rect 521052 385532 521108 385588
rect 81452 385420 81508 385476
rect 367052 385308 367108 385364
rect 367052 384972 367108 385028
rect 19964 384860 20020 384916
rect 349468 384524 349524 384580
rect 74844 384300 74900 384356
rect 203196 383740 203252 383796
rect 581308 383740 581364 383796
rect 259644 383180 259700 383236
rect 347788 383180 347844 383236
rect 263788 382620 263844 382676
rect 265020 382060 265076 382116
rect 206108 381500 206164 381556
rect 371308 381500 371364 381556
rect 392252 381276 392308 381332
rect 396732 381276 396788 381332
rect 579628 380940 579684 380996
rect 133532 380716 133588 380772
rect 264908 380716 264964 380772
rect 335244 380492 335300 380548
rect 455420 380492 455476 380548
rect 204876 380380 204932 380436
rect 533372 379820 533428 379876
rect 530012 379260 530068 379316
rect 79772 379036 79828 379092
rect 264796 379036 264852 379092
rect 18172 378924 18228 378980
rect 257852 378924 257908 378980
rect 19740 378812 19796 378868
rect 264572 378812 264628 378868
rect 335132 378812 335188 378868
rect 395052 378812 395108 378868
rect 256172 378700 256228 378756
rect 533484 377580 533540 377636
rect 69692 377132 69748 377188
rect 264684 377132 264740 377188
rect 141036 377020 141092 377076
rect 476252 377020 476308 377076
rect 519148 376460 519204 376516
rect 519932 375900 519988 375956
rect 336140 375452 336196 375508
rect 458780 375452 458836 375508
rect 461132 375340 461188 375396
rect 400652 374780 400708 374836
rect 142716 374220 142772 374276
rect 517468 373660 517524 373716
rect 467852 372540 467908 372596
rect 76412 372092 76468 372148
rect 263788 372092 263844 372148
rect 192332 371980 192388 372036
rect 464492 371980 464548 372036
rect 205772 371420 205828 371476
rect 503132 371420 503188 371476
rect 264908 370300 264964 370356
rect 336140 370300 336196 370356
rect 335244 369740 335300 369796
rect 127036 369180 127092 369236
rect 457212 369180 457268 369236
rect 334572 368732 334628 368788
rect 394940 368732 394996 368788
rect 455308 368620 455364 368676
rect 127260 368060 127316 368116
rect 457324 367500 457380 367556
rect 334348 367052 334404 367108
rect 402332 367052 402388 367108
rect 398972 366940 399028 366996
rect 126924 366380 126980 366436
rect 457100 366380 457156 366436
rect 334460 365484 334516 365540
rect 396508 365484 396564 365540
rect 393148 365372 393204 365428
rect 459004 365372 459060 365428
rect 126812 365260 126868 365316
rect 456092 365260 456148 365316
rect 127148 364700 127204 364756
rect 334348 364700 334404 364756
rect 143612 364140 143668 364196
rect 393148 364140 393204 364196
rect 257852 363580 257908 363636
rect 335132 363580 335188 363636
rect 263788 363020 263844 363076
rect 334460 363020 334516 363076
rect 18284 362460 18340 362516
rect 334572 362460 334628 362516
rect 335916 362012 335972 362068
rect 394828 362012 394884 362068
rect 18060 361900 18116 361956
rect 392252 361900 392308 361956
rect 264684 361340 264740 361396
rect 345212 360780 345268 360836
rect 64876 360220 64932 360276
rect 341852 360220 341908 360276
rect 64652 359660 64708 359716
rect 264796 358540 264852 358596
rect 338492 357980 338548 358036
rect 264572 357420 264628 357476
rect 335916 357420 335972 357476
rect 205660 356860 205716 356916
rect 581308 356300 581364 356356
rect 581420 355852 581476 355908
rect 206668 355740 206724 355796
rect 583100 355740 583156 355796
rect 518252 355404 518308 355460
rect 264796 355180 264852 355236
rect 206220 354172 206276 354228
rect 204764 354060 204820 354116
rect 580412 354060 580468 354116
rect 351036 353052 351092 353108
rect 535164 353052 535220 353108
rect 265132 352940 265188 352996
rect 579628 352940 579684 352996
rect 352604 352828 352660 352884
rect 583212 352828 583268 352884
rect 202972 352604 203028 352660
rect 206668 352604 206724 352660
rect 264572 352380 264628 352436
rect 351036 352380 351092 352436
rect 263340 351820 263396 351876
rect 352604 351260 352660 351316
rect 202860 351036 202916 351092
rect 205660 351036 205716 351092
rect 334460 350700 334516 350756
rect 263788 350140 263844 350196
rect 393372 349916 393428 349972
rect 473228 349692 473284 349748
rect 263788 347900 263844 347956
rect 260092 347340 260148 347396
rect 262108 346220 262164 346276
rect 263788 345660 263844 345716
rect 334460 345660 334516 345716
rect 263900 345100 263956 345156
rect 334348 345100 334404 345156
rect 263788 343980 263844 344036
rect 334460 343420 334516 343476
rect 263788 342300 263844 342356
rect 334348 342300 334404 342356
rect 580412 341740 580468 341796
rect 20076 341628 20132 341684
rect 82684 341628 82740 341684
rect 141036 341628 141092 341684
rect 144060 341628 144116 341684
rect 473676 341628 473732 341684
rect 476028 341628 476084 341684
rect 534268 341628 534324 341684
rect 263788 341180 263844 341236
rect 334460 341180 334516 341236
rect 352604 341180 352660 341236
rect 201292 340956 201348 341012
rect 263900 340620 263956 340676
rect 334348 340620 334404 340676
rect 414652 340956 414708 341012
rect 394044 340396 394100 340452
rect 455420 340396 455476 340452
rect 82460 340284 82516 340340
rect 127484 340284 127540 340340
rect 141036 340284 141092 340340
rect 189532 340284 189588 340340
rect 264572 340284 264628 340340
rect 65212 339612 65268 339668
rect 334460 340060 334516 340116
rect 518252 340284 518308 340340
rect 581420 340284 581476 340340
rect 393372 339724 393428 339780
rect 200956 339612 201012 339668
rect 345212 339612 345268 339668
rect 455532 339612 455588 339668
rect 473228 339612 473284 339668
rect 263788 339500 263844 339556
rect 457772 339500 457828 339556
rect 126140 339276 126196 339332
rect 130060 339276 130116 339332
rect 18060 338940 18116 338996
rect 334348 338940 334404 338996
rect 341852 338940 341908 338996
rect 472892 338940 472948 338996
rect 517468 338716 517524 338772
rect 127484 338492 127540 338548
rect 143612 338492 143668 338548
rect 189532 338492 189588 338548
rect 204092 338492 204148 338548
rect 337708 338380 337764 338436
rect 127596 338268 127652 338324
rect 206108 338268 206164 338324
rect 334460 337820 334516 337876
rect 455308 337820 455364 337876
rect 82236 337596 82292 337652
rect 140924 337596 140980 337652
rect 192444 337596 192500 337652
rect 261212 337596 261268 337652
rect 141932 337372 141988 337428
rect 334348 337260 334404 337316
rect 517468 337596 517524 337652
rect 583100 337596 583156 337652
rect 393484 337036 393540 337092
rect 64092 336924 64148 336980
rect 127596 336924 127652 336980
rect 188972 336924 189028 336980
rect 265132 336924 265188 336980
rect 264572 336700 264628 336756
rect 334460 336700 334516 336756
rect 520828 336924 520884 336980
rect 581308 336924 581364 336980
rect 455308 336812 455364 336868
rect 20636 336364 20692 336420
rect 80556 336364 80612 336420
rect 396508 336364 396564 336420
rect 18284 336252 18340 336308
rect 64204 336252 64260 336308
rect 195804 336252 195860 336308
rect 204876 336252 204932 336308
rect 264796 336252 264852 336308
rect 334460 336140 334516 336196
rect 394828 336028 394884 336084
rect 64764 335580 64820 335636
rect 195692 335580 195748 335636
rect 264012 335580 264068 335636
rect 351148 335580 351204 335636
rect 455532 335580 455588 335636
rect 519148 335580 519204 335636
rect 260316 335020 260372 335076
rect 334460 335020 334516 335076
rect 18396 334908 18452 334964
rect 334460 334460 334516 334516
rect 461132 334908 461188 334964
rect 582988 334908 583044 334964
rect 206220 334236 206276 334292
rect 251020 334236 251076 334292
rect 264908 333900 264964 333956
rect 394940 334236 394996 334292
rect 399756 334236 399812 334292
rect 535164 334236 535220 334292
rect 393372 333676 393428 333732
rect 126140 333564 126196 333620
rect 189084 333564 189140 333620
rect 202972 333564 203028 333620
rect 455644 333564 455700 333620
rect 473116 333564 473172 333620
rect 534268 333564 534324 333620
rect 579628 333564 579684 333620
rect 264684 333340 264740 333396
rect 334460 333340 334516 333396
rect 20076 332892 20132 332948
rect 64652 332892 64708 332948
rect 127596 332892 127652 332948
rect 192332 332892 192388 332948
rect 204764 332892 204820 332948
rect 456092 333452 456148 333508
rect 473228 333452 473284 333508
rect 263788 332780 263844 332836
rect 521052 332892 521108 332948
rect 523292 332892 523348 332948
rect 396844 332668 396900 332724
rect 18172 332220 18228 332276
rect 69692 332220 69748 332276
rect 205772 332220 205828 332276
rect 261324 332220 261380 332276
rect 393932 332220 393988 332276
rect 455308 332220 455364 332276
rect 520940 332220 520996 332276
rect 523292 332220 523348 332276
rect 263900 331660 263956 331716
rect 334460 331660 334516 331716
rect 579628 331660 579684 331716
rect 64204 331548 64260 331604
rect 189420 331548 189476 331604
rect 80556 331436 80612 331492
rect 81452 331436 81508 331492
rect 455308 331212 455364 331268
rect 263788 331100 263844 331156
rect 203084 330876 203140 330932
rect 395612 330876 395668 330932
rect 396508 330876 396564 330932
rect 535052 330876 535108 330932
rect 205996 330652 206052 330708
rect 126812 330204 126868 330260
rect 263788 330540 263844 330596
rect 251916 330204 251972 330260
rect 338492 330204 338548 330260
rect 334460 329980 334516 330036
rect 80444 329644 80500 329700
rect 407372 330204 407428 330260
rect 394828 329644 394884 329700
rect 127596 329532 127652 329588
rect 202860 329532 202916 329588
rect 259532 329532 259588 329588
rect 393260 329532 393316 329588
rect 344428 329420 344484 329476
rect 80556 329308 80612 329364
rect 197372 328860 197428 328916
rect 263900 328860 263956 328916
rect 338604 328860 338660 328916
rect 455532 328860 455588 328916
rect 455420 328636 455476 328692
rect 263788 327740 263844 327796
rect 334460 327740 334516 327796
rect 334460 327180 334516 327236
rect 350252 326620 350308 326676
rect 334348 326060 334404 326116
rect 263788 325500 263844 325556
rect 583212 325500 583268 325556
rect 251020 324940 251076 324996
rect 334460 324380 334516 324436
rect 263788 323820 263844 323876
rect 334460 323820 334516 323876
rect 259532 322700 259588 322756
rect 334348 322700 334404 322756
rect 261212 322140 261268 322196
rect 251916 321580 251972 321636
rect 334460 321580 334516 321636
rect 261324 320460 261380 320516
rect 351932 320460 351988 320516
rect 334460 319900 334516 319956
rect 140924 319116 140980 319172
rect 142828 319116 142884 319172
rect 334460 318780 334516 318836
rect 456876 318444 456932 318500
rect 473116 318444 473172 318500
rect 188972 318332 189028 318388
rect 204988 318332 205044 318388
rect 456204 318332 456260 318388
rect 472892 318332 472948 318388
rect 520828 317548 520884 317604
rect 204988 316988 205044 317044
rect 142828 316540 142884 316596
rect 519148 316540 519204 316596
rect 204092 315980 204148 316036
rect 456876 315420 456932 315476
rect 80444 314636 80500 314692
rect 161308 314636 161364 314692
rect 261436 314524 261492 314580
rect 456092 314860 456148 314916
rect 141036 314300 141092 314356
rect 261436 314300 261492 314356
rect 517468 314300 517524 314356
rect 562940 314076 562996 314132
rect 205772 313628 205828 313684
rect 126812 313292 126868 313348
rect 198156 313292 198212 313348
rect 456204 313180 456260 313236
rect 200956 312620 201012 312676
rect 80556 312060 80612 312116
rect 161308 311500 161364 311556
rect 143612 310380 143668 310436
rect 198156 309260 198212 309316
rect 69692 308252 69748 308308
rect 263788 308252 263844 308308
rect 81452 308140 81508 308196
rect 141932 307580 141988 307636
rect 393932 307580 393988 307636
rect 457772 305900 457828 305956
rect 345212 305340 345268 305396
rect 64764 304780 64820 304836
rect 263788 304220 263844 304276
rect 64652 303660 64708 303716
rect 396844 302540 396900 302596
rect 18284 301980 18340 302036
rect 341852 300860 341908 300916
rect 18172 299740 18228 299796
rect 338492 299740 338548 299796
rect 18396 299180 18452 299236
rect 395612 299180 395668 299236
rect 264572 298620 264628 298676
rect 202972 295820 203028 295876
rect 583548 295260 583604 295316
rect 203084 294700 203140 294756
rect 582092 294700 582148 294756
rect 580412 294140 580468 294196
rect 204764 293580 204820 293636
rect 581308 293580 581364 293636
rect 206108 293020 206164 293076
rect 523292 293020 523348 293076
rect 252812 292460 252868 292516
rect 580524 292460 580580 292516
rect 430108 291900 430164 291956
rect 204876 291340 204932 291396
rect 502348 291340 502404 291396
rect 263788 290780 263844 290836
rect 335916 290780 335972 290836
rect 189196 290220 189252 290276
rect 449372 290220 449428 290276
rect 140924 289772 140980 289828
rect 263788 289772 263844 289828
rect 335916 289772 335972 289828
rect 517468 289772 517524 289828
rect 517580 289660 517636 289716
rect 188972 289100 189028 289156
rect 519148 289100 519204 289156
rect 334460 288092 334516 288148
rect 200732 287980 200788 288036
rect 334460 287868 334516 287924
rect 352716 286860 352772 286916
rect 502348 286412 502404 286468
rect 583100 286412 583156 286468
rect 263788 285740 263844 285796
rect 464492 285740 464548 285796
rect 259532 285628 259588 285684
rect 264572 285628 264628 285684
rect 144060 284844 144116 284900
rect 261212 284844 261268 284900
rect 449372 284844 449428 284900
rect 521052 284844 521108 284900
rect 430108 284732 430164 284788
rect 535164 284732 535220 284788
rect 205772 284620 205828 284676
rect 473116 284508 473172 284564
rect 261212 284396 261268 284452
rect 342636 284060 342692 284116
rect 204092 283500 204148 283556
rect 142716 283164 142772 283220
rect 263788 283164 263844 283220
rect 342636 283164 342692 283220
rect 472892 283164 472948 283220
rect 473116 283164 473172 283220
rect 520828 283164 520884 283220
rect 352716 283052 352772 283108
rect 520940 283052 520996 283108
rect 523292 283052 523348 283108
rect 583212 283052 583268 283108
rect 138572 282940 138628 282996
rect 456988 282940 457044 282996
rect 80332 282380 80388 282436
rect 455308 282380 455364 282436
rect 136892 281820 136948 281876
rect 456092 281820 456148 281876
rect 130284 281596 130340 281652
rect 334460 281596 334516 281652
rect 458780 281596 458836 281652
rect 82012 281484 82068 281540
rect 457772 281484 457828 281540
rect 263788 279580 263844 279636
rect 334460 279580 334516 279636
rect 455420 279356 455476 279412
rect 204764 279132 204820 279188
rect 263340 279020 263396 279076
rect 334460 278460 334516 278516
rect 520828 278460 520884 278516
rect 262108 277340 262164 277396
rect 64204 277116 64260 277172
rect 455308 277116 455364 277172
rect 263788 276780 263844 276836
rect 334460 276780 334516 276836
rect 262220 275660 262276 275716
rect 334348 275660 334404 275716
rect 249452 275100 249508 275156
rect 336924 275100 336980 275156
rect 334572 274540 334628 274596
rect 334460 273980 334516 274036
rect 334348 273420 334404 273476
rect 262108 272860 262164 272916
rect 351036 272860 351092 272916
rect 263788 272300 263844 272356
rect 334460 272300 334516 272356
rect 263900 271740 263956 271796
rect 464492 271292 464548 271348
rect 473004 271292 473060 271348
rect 141036 271068 141092 271124
rect 144060 271068 144116 271124
rect 201628 271068 201684 271124
rect 20076 270396 20132 270452
rect 82460 270396 82516 270452
rect 127596 270396 127652 270452
rect 534268 270396 534324 270452
rect 64204 269724 64260 269780
rect 334460 270060 334516 270116
rect 130172 269724 130228 269780
rect 457212 269724 457268 269780
rect 473676 269724 473732 269780
rect 263788 269500 263844 269556
rect 414652 269500 414708 269556
rect 64092 269052 64148 269108
rect 127484 269052 127540 269108
rect 404012 269052 404068 269108
rect 458892 269052 458948 269108
rect 472108 269052 472164 269108
rect 583212 269052 583268 269108
rect 335692 268940 335748 268996
rect 457772 268716 457828 268772
rect 458668 268716 458724 268772
rect 18396 268380 18452 268436
rect 141036 268380 141092 268436
rect 189532 268380 189588 268436
rect 20076 267708 20132 267764
rect 64204 267708 64260 267764
rect 205772 267708 205828 267764
rect 334348 268380 334404 268436
rect 352716 268380 352772 268436
rect 410732 268380 410788 268436
rect 455532 268380 455588 268436
rect 472108 268380 472164 268436
rect 534268 268380 534324 268436
rect 263788 267820 263844 267876
rect 338492 267708 338548 267764
rect 206444 267596 206500 267652
rect 583100 267708 583156 267764
rect 334460 267260 334516 267316
rect 517468 267260 517524 267316
rect 203084 267036 203140 267092
rect 262444 267036 262500 267092
rect 345212 267036 345268 267092
rect 395052 267036 395108 267092
rect 579292 267036 579348 267092
rect 82460 266924 82516 266980
rect 263788 266700 263844 266756
rect 189532 266588 189588 266644
rect 199836 266588 199892 266644
rect 130284 266364 130340 266420
rect 142604 266364 142660 266420
rect 189532 266364 189588 266420
rect 204876 266364 204932 266420
rect 259532 266364 259588 266420
rect 407372 266364 407428 266420
rect 472108 266364 472164 266420
rect 583548 266364 583604 266420
rect 335692 266252 335748 266308
rect 347788 266252 347844 266308
rect 393372 266252 393428 266308
rect 206332 266140 206388 266196
rect 263788 266140 263844 266196
rect 334460 266140 334516 266196
rect 64652 265692 64708 265748
rect 80444 265692 80500 265748
rect 126812 265692 126868 265748
rect 262220 265692 262276 265748
rect 336812 265692 336868 265748
rect 582092 266140 582148 266196
rect 456988 265692 457044 265748
rect 461132 265692 461188 265748
rect 517804 265692 517860 265748
rect 260316 265580 260372 265636
rect 69692 265020 69748 265076
rect 127596 265020 127652 265076
rect 133532 265020 133588 265076
rect 140924 265020 140980 265076
rect 206108 265020 206164 265076
rect 394940 265020 394996 265076
rect 402332 265020 402388 265076
rect 458668 265020 458724 265076
rect 393372 264796 393428 264852
rect 264012 264460 264068 264516
rect 334460 264460 334516 264516
rect 136892 264348 136948 264404
rect 202972 264348 203028 264404
rect 348572 264348 348628 264404
rect 464492 264572 464548 264628
rect 472108 264572 472164 264628
rect 473004 264348 473060 264404
rect 520940 264348 520996 264404
rect 579292 264348 579348 264404
rect 334460 263900 334516 263956
rect 580412 263788 580468 263844
rect 64204 263676 64260 263732
rect 126812 263676 126868 263732
rect 64204 263004 64260 263060
rect 80332 263004 80388 263060
rect 127596 263004 127652 263060
rect 189196 263676 189252 263732
rect 396620 263676 396676 263732
rect 472892 263676 472948 263732
rect 262332 263340 262388 263396
rect 579628 263228 579684 263284
rect 204092 263004 204148 263060
rect 144284 262780 144340 262836
rect 394828 263004 394884 263060
rect 534268 263004 534324 263060
rect 262108 262780 262164 262836
rect 334460 262780 334516 262836
rect 82684 262332 82740 262388
rect 396956 262332 397012 262388
rect 521052 262332 521108 262388
rect 582988 262332 583044 262388
rect 194908 261996 194964 262052
rect 468636 261996 468692 262052
rect 580524 261996 580580 262052
rect 64764 261660 64820 261716
rect 262220 261660 262276 261716
rect 334460 261660 334516 261716
rect 396844 261660 396900 261716
rect 398972 261660 399028 261716
rect 457100 261660 457156 261716
rect 206444 261548 206500 261604
rect 64204 261212 64260 261268
rect 81452 261212 81508 261268
rect 135212 260988 135268 261044
rect 142716 260988 142772 261044
rect 393484 261436 393540 261492
rect 262444 261100 262500 261156
rect 262108 260988 262164 261044
rect 348796 260988 348852 261044
rect 458780 260988 458836 261044
rect 472220 260988 472276 261044
rect 579292 260988 579348 261044
rect 334460 260540 334516 260596
rect 64652 260316 64708 260372
rect 82012 260316 82068 260372
rect 138572 260316 138628 260372
rect 144060 260316 144116 260372
rect 200732 260316 200788 260372
rect 393260 260316 393316 260372
rect 472108 260316 472164 260372
rect 519148 260316 519204 260372
rect 263788 259980 263844 260036
rect 334460 259980 334516 260036
rect 133532 259644 133588 259700
rect 346892 259644 346948 259700
rect 396620 259644 396676 259700
rect 581308 259644 581364 259700
rect 395612 259532 395668 259588
rect 456876 259532 456932 259588
rect 472220 259532 472276 259588
rect 263900 259420 263956 259476
rect 188972 258972 189028 259028
rect 262332 258972 262388 259028
rect 334460 258860 334516 258916
rect 456092 258636 456148 258692
rect 81564 258300 81620 258356
rect 252812 258300 252868 258356
rect 263788 258300 263844 258356
rect 334460 258300 334516 258356
rect 517692 258300 517748 258356
rect 535164 258300 535220 258356
rect 517468 258076 517524 258132
rect 263900 257740 263956 257796
rect 334348 257740 334404 257796
rect 264012 257628 264068 257684
rect 455308 257628 455364 257684
rect 259980 257180 260036 257236
rect 262556 256620 262612 256676
rect 351932 256620 351988 256676
rect 351036 256060 351092 256116
rect 334572 255500 334628 255556
rect 334460 254940 334516 254996
rect 334684 254380 334740 254436
rect 263788 253820 263844 253876
rect 334348 253820 334404 253876
rect 263788 253260 263844 253316
rect 64764 252812 64820 252868
rect 80556 252812 80612 252868
rect 263900 252700 263956 252756
rect 334460 252700 334516 252756
rect 334460 251580 334516 251636
rect 263788 251020 263844 251076
rect 351036 251020 351092 251076
rect 263788 250460 263844 250516
rect 334348 250460 334404 250516
rect 260316 248780 260372 248836
rect 334460 248780 334516 248836
rect 334460 248220 334516 248276
rect 351036 247660 351092 247716
rect 338492 247100 338548 247156
rect 346892 246540 346948 246596
rect 336028 246204 336084 246260
rect 348572 246204 348628 246260
rect 348796 245980 348852 246036
rect 351036 245756 351092 245812
rect 410732 245756 410788 245812
rect 18396 245308 18452 245364
rect 20972 245308 21028 245364
rect 64652 245196 64708 245252
rect 80556 244860 80612 244916
rect 345212 244860 345268 244916
rect 345996 244412 346052 244468
rect 396620 244412 396676 244468
rect 81564 244300 81620 244356
rect 336812 244300 336868 244356
rect 336028 243740 336084 243796
rect 69692 243180 69748 243236
rect 81452 242620 81508 242676
rect 395052 242620 395108 242676
rect 20972 242060 21028 242116
rect 394940 241500 394996 241556
rect 20076 240940 20132 240996
rect 345996 240940 346052 240996
rect 248556 239820 248612 239876
rect 335916 239820 335972 239876
rect 263788 239260 263844 239316
rect 263900 238700 263956 238756
rect 335692 238700 335748 238756
rect 335132 237020 335188 237076
rect 203196 236460 203252 236516
rect 400652 236460 400708 236516
rect 204876 236012 204932 236068
rect 263788 236012 263844 236068
rect 264908 235900 264964 235956
rect 257852 235340 257908 235396
rect 263900 235340 263956 235396
rect 581308 235340 581364 235396
rect 262892 235116 262948 235172
rect 261212 234780 261268 234836
rect 203084 234556 203140 234612
rect 248556 234556 248612 234612
rect 256172 234220 256228 234276
rect 459452 234220 459508 234276
rect 583436 233660 583492 233716
rect 257964 233436 258020 233492
rect 140588 232540 140644 232596
rect 462812 231980 462868 232036
rect 140700 231420 140756 231476
rect 518364 231420 518420 231476
rect 335916 230972 335972 231028
rect 583100 230972 583156 231028
rect 140812 230300 140868 230356
rect 140924 229740 140980 229796
rect 519932 229740 519988 229796
rect 418348 229180 418404 229236
rect 520156 228620 520212 228676
rect 189196 228060 189252 228116
rect 396172 228060 396228 228116
rect 188972 227500 189028 227556
rect 518252 226940 518308 226996
rect 197372 226380 197428 226436
rect 263900 225820 263956 225876
rect 263788 225260 263844 225316
rect 338492 225260 338548 225316
rect 80332 224700 80388 224756
rect 418348 224364 418404 224420
rect 520940 224364 520996 224420
rect 144060 224252 144116 224308
rect 263788 224252 263844 224308
rect 335132 224252 335188 224308
rect 581420 224252 581476 224308
rect 126812 223580 126868 223636
rect 419132 223580 419188 223636
rect 80108 223020 80164 223076
rect 192332 222572 192388 222628
rect 263900 222572 263956 222628
rect 80444 222460 80500 222516
rect 455308 222460 455364 222516
rect 126924 221900 126980 221956
rect 83132 221340 83188 221396
rect 351932 221340 351988 221396
rect 130172 220780 130228 220836
rect 335916 220780 335972 220836
rect 263788 220220 263844 220276
rect 407372 219660 407428 219716
rect 82012 219212 82068 219268
rect 263788 219212 263844 219268
rect 335692 219212 335748 219268
rect 579628 219212 579684 219268
rect 339276 219100 339332 219156
rect 263788 218540 263844 218596
rect 356188 217980 356244 218036
rect 82236 217532 82292 217588
rect 263788 217532 263844 217588
rect 335916 217532 335972 217588
rect 456988 217532 457044 217588
rect 263788 216300 263844 216356
rect 336028 216300 336084 216356
rect 252812 215852 252868 215908
rect 264908 215852 264964 215908
rect 263900 215740 263956 215796
rect 337036 215180 337092 215236
rect 74732 214620 74788 214676
rect 340396 214620 340452 214676
rect 356188 214396 356244 214452
rect 410732 214396 410788 214452
rect 336028 214284 336084 214340
rect 396732 214284 396788 214340
rect 419132 214284 419188 214340
rect 458892 214284 458948 214340
rect 459452 214284 459508 214340
rect 535276 214284 535332 214340
rect 81452 214172 81508 214228
rect 263788 214172 263844 214228
rect 338492 214172 338548 214228
rect 472108 214172 472164 214228
rect 206668 214060 206724 214116
rect 340620 214060 340676 214116
rect 263788 213500 263844 213556
rect 340172 213500 340228 213556
rect 73052 213276 73108 213332
rect 263900 213276 263956 213332
rect 261100 213164 261156 213220
rect 339276 213164 339332 213220
rect 458780 213164 458836 213220
rect 395836 213052 395892 213108
rect 396172 213052 396228 213108
rect 521164 213052 521220 213108
rect 160188 212828 160244 212884
rect 231532 212828 231588 212884
rect 334460 212828 334516 212884
rect 370860 212828 370916 212884
rect 375788 212828 375844 212884
rect 231756 212716 231812 212772
rect 160188 212604 160244 212660
rect 334460 212604 334516 212660
rect 375788 212604 375844 212660
rect 396620 212604 396676 212660
rect 231532 212380 231588 212436
rect 231756 212380 231812 212436
rect 370860 212380 370916 212436
rect 261100 212156 261156 212212
rect 74844 212044 74900 212100
rect 263788 212044 263844 212100
rect 338492 211820 338548 211876
rect 79996 211596 80052 211652
rect 83132 211596 83188 211652
rect 396396 211260 396452 211316
rect 80220 211148 80276 211204
rect 130172 211148 130228 211204
rect 351932 211148 351988 211204
rect 410844 211148 410900 211204
rect 462812 211148 462868 211204
rect 521052 211148 521108 211204
rect 64652 211036 64708 211092
rect 206668 211036 206724 211092
rect 400652 210924 400708 210980
rect 583324 210924 583380 210980
rect 81676 210700 81732 210756
rect 396844 210700 396900 210756
rect 351148 210588 351204 210644
rect 535164 210588 535220 210644
rect 345996 210476 346052 210532
rect 535500 210476 535556 210532
rect 20076 210364 20132 210420
rect 263788 210364 263844 210420
rect 351036 210364 351092 210420
rect 583212 210364 583268 210420
rect 340284 210140 340340 210196
rect 263788 209580 263844 209636
rect 251916 209020 251972 209076
rect 351036 209020 351092 209076
rect 144060 208572 144116 208628
rect 472108 208572 472164 208628
rect 351148 207900 351204 207956
rect 262108 206780 262164 206836
rect 258076 206220 258132 206276
rect 334460 206220 334516 206276
rect 261212 205884 261268 205940
rect 264796 205660 264852 205716
rect 264572 205100 264628 205156
rect 334460 204540 334516 204596
rect 345996 203420 346052 203476
rect 334460 202300 334516 202356
rect 341852 201740 341908 201796
rect 334460 200620 334516 200676
rect 141036 199836 141092 199892
rect 201628 199836 201684 199892
rect 396508 199164 396564 199220
rect 534268 199164 534324 199220
rect 414652 199052 414708 199108
rect 18396 198940 18452 198996
rect 263788 198940 263844 198996
rect 334460 198940 334516 198996
rect 82684 198492 82740 198548
rect 140700 198492 140756 198548
rect 352716 198492 352772 198548
rect 455308 198492 455364 198548
rect 80332 197820 80388 197876
rect 263900 197820 263956 197876
rect 334348 197820 334404 197876
rect 473676 197820 473732 197876
rect 263788 197260 263844 197316
rect 334460 197260 334516 197316
rect 64204 197148 64260 197204
rect 197372 197148 197428 197204
rect 579628 197148 579684 197204
rect 248556 196700 248612 196756
rect 455420 196700 455476 196756
rect 395836 196588 395892 196644
rect 396508 196588 396564 196644
rect 196588 196476 196644 196532
rect 337036 196476 337092 196532
rect 394828 196476 394884 196532
rect 410844 196476 410900 196532
rect 467852 196476 467908 196532
rect 520940 196476 520996 196532
rect 524972 196476 525028 196532
rect 583324 196476 583380 196532
rect 520156 196364 520212 196420
rect 263788 196140 263844 196196
rect 334460 196140 334516 196196
rect 20636 196028 20692 196084
rect 189532 195804 189588 195860
rect 340620 195804 340676 195860
rect 535500 195804 535556 195860
rect 581420 195804 581476 195860
rect 64204 195132 64260 195188
rect 80444 195132 80500 195188
rect 127484 195132 127540 195188
rect 189196 195132 189252 195188
rect 202972 195132 203028 195188
rect 262892 195132 262948 195188
rect 340396 195132 340452 195188
rect 396732 195132 396788 195188
rect 411180 195132 411236 195188
rect 535276 195132 535332 195188
rect 20300 194908 20356 194964
rect 20076 194460 20132 194516
rect 81676 194572 81732 194628
rect 79996 194460 80052 194516
rect 127596 194460 127652 194516
rect 257964 194460 258020 194516
rect 334460 194460 334516 194516
rect 340172 194460 340228 194516
rect 411292 194460 411348 194516
rect 455308 194012 455364 194068
rect 81452 193900 81508 193956
rect 334348 193900 334404 193956
rect 80220 193788 80276 193844
rect 192332 193788 192388 193844
rect 264796 193788 264852 193844
rect 456988 193788 457044 193844
rect 472108 193788 472164 193844
rect 264012 193340 264068 193396
rect 334460 193340 334516 193396
rect 519932 193228 519988 193284
rect 188972 193116 189028 193172
rect 396508 193116 396564 193172
rect 535164 193116 535220 193172
rect 583100 193116 583156 193172
rect 334348 192668 334404 192724
rect 351820 192668 351876 192724
rect 74844 192444 74900 192500
rect 126924 192444 126980 192500
rect 140812 192444 140868 192500
rect 340284 192444 340340 192500
rect 411180 192444 411236 192500
rect 521052 192444 521108 192500
rect 189532 192332 189588 192388
rect 204988 192332 205044 192388
rect 463596 192332 463652 192388
rect 472108 192332 472164 192388
rect 334460 192220 334516 192276
rect 205660 191772 205716 191828
rect 256172 191772 256228 191828
rect 396732 191772 396788 191828
rect 410732 191772 410788 191828
rect 458892 191772 458948 191828
rect 263788 191660 263844 191716
rect 518364 191436 518420 191492
rect 127596 191100 127652 191156
rect 264572 191212 264628 191268
rect 258412 191100 258468 191156
rect 338492 191100 338548 191156
rect 407372 191100 407428 191156
rect 458780 191100 458836 191156
rect 472108 191100 472164 191156
rect 334348 190540 334404 190596
rect 80108 190428 80164 190484
rect 252812 190428 252868 190484
rect 579740 190988 579796 191044
rect 262108 189980 262164 190036
rect 336028 189980 336084 190036
rect 73052 189756 73108 189812
rect 189532 189756 189588 189812
rect 257852 189756 257908 189812
rect 472108 189756 472164 189812
rect 519148 189756 519204 189812
rect 583436 189756 583492 189812
rect 263788 189420 263844 189476
rect 347788 189420 347844 189476
rect 126812 189084 126868 189140
rect 204876 189084 204932 189140
rect 258076 189084 258132 189140
rect 396620 189084 396676 189140
rect 581308 189084 581364 189140
rect 455420 188972 455476 189028
rect 74732 188412 74788 188468
rect 134428 188412 134484 188468
rect 140924 188412 140980 188468
rect 346108 188412 346164 188468
rect 396844 188412 396900 188468
rect 263900 188300 263956 188356
rect 20076 188188 20132 188244
rect 82124 187740 82180 187796
rect 140588 187740 140644 187796
rect 197484 187740 197540 187796
rect 203084 187740 203140 187796
rect 64652 187068 64708 187124
rect 82236 187068 82292 187124
rect 203196 187068 203252 187124
rect 251916 187068 251972 187124
rect 472108 187068 472164 187124
rect 583212 187068 583268 187124
rect 258636 186620 258692 186676
rect 342636 186620 342692 186676
rect 82684 186396 82740 186452
rect 393260 186396 393316 186452
rect 455308 186396 455364 186452
rect 456092 186284 456148 186340
rect 263788 185500 263844 185556
rect 346108 185500 346164 185556
rect 248556 184940 248612 184996
rect 336140 184380 336196 184436
rect 263900 183820 263956 183876
rect 335132 183260 335188 183316
rect 261436 182140 261492 182196
rect 521164 181692 521220 181748
rect 264572 181580 264628 181636
rect 338492 181020 338548 181076
rect 252812 179900 252868 179956
rect 345212 179900 345268 179956
rect 262892 179340 262948 179396
rect 257852 178780 257908 178836
rect 256396 178220 256452 178276
rect 264684 177660 264740 177716
rect 335356 177660 335412 177716
rect 350252 177100 350308 177156
rect 334460 176540 334516 176596
rect 518252 176316 518308 176372
rect 263788 175980 263844 176036
rect 348572 175980 348628 176036
rect 341852 175420 341908 175476
rect 351932 174860 351988 174916
rect 206108 173964 206164 174020
rect 263788 173964 263844 174020
rect 334460 173852 334516 173908
rect 579628 173852 579684 173908
rect 140812 173740 140868 173796
rect 462812 173740 462868 173796
rect 517468 173180 517524 173236
rect 350364 172620 350420 172676
rect 204876 172172 204932 172228
rect 264684 172172 264740 172228
rect 345436 172060 345492 172116
rect 336028 171500 336084 171556
rect 380492 170940 380548 170996
rect 336028 170492 336084 170548
rect 520828 170492 520884 170548
rect 461356 170380 461412 170436
rect 188972 169820 189028 169876
rect 338940 169260 338996 169316
rect 263900 168700 263956 168756
rect 263788 168140 263844 168196
rect 197372 167580 197428 167636
rect 519148 167580 519204 167636
rect 199052 167020 199108 167076
rect 356972 166460 357028 166516
rect 455308 165340 455364 165396
rect 338604 164780 338660 164836
rect 127148 164220 127204 164276
rect 195692 163772 195748 163828
rect 263788 163772 263844 163828
rect 341852 163772 341908 163828
rect 582988 163772 583044 163828
rect 126924 163660 126980 163716
rect 127372 163100 127428 163156
rect 452732 163100 452788 163156
rect 127260 162540 127316 162596
rect 457772 162540 457828 162596
rect 192332 162092 192388 162148
rect 263900 162092 263956 162148
rect 456092 161980 456148 162036
rect 126812 161420 126868 161476
rect 127484 160860 127540 160916
rect 338940 160524 338996 160580
rect 520940 160524 520996 160580
rect 390572 160300 390628 160356
rect 127036 159740 127092 159796
rect 335356 158732 335412 158788
rect 581308 158732 581364 158788
rect 64876 158620 64932 158676
rect 352044 158620 352100 158676
rect 395612 158060 395668 158116
rect 64988 157500 65044 157556
rect 390460 157500 390516 157556
rect 390572 157276 390628 157332
rect 459004 157276 459060 157332
rect 338604 157164 338660 157220
rect 410844 157164 410900 157220
rect 348572 157052 348628 157108
rect 583212 157052 583268 157108
rect 64764 156940 64820 156996
rect 395724 156940 395780 156996
rect 18172 156380 18228 156436
rect 341852 156380 341908 156436
rect 357196 155820 357252 155876
rect 356972 155596 357028 155652
rect 458780 155596 458836 155652
rect 338492 155484 338548 155540
rect 535052 155484 535108 155540
rect 351932 155372 351988 155428
rect 583100 155372 583156 155428
rect 395836 155260 395892 155316
rect 64652 154700 64708 154756
rect 392252 154700 392308 154756
rect 264684 153020 264740 153076
rect 380492 152124 380548 152180
rect 473004 152124 473060 152180
rect 263788 151340 263844 151396
rect 396508 151340 396564 151396
rect 261324 150780 261380 150836
rect 81452 150444 81508 150500
rect 263788 150444 263844 150500
rect 259980 150220 260036 150276
rect 526652 150220 526708 150276
rect 259756 149660 259812 149716
rect 524972 149660 525028 149716
rect 523292 149100 523348 149156
rect 449372 148540 449428 148596
rect 203084 147420 203140 147476
rect 581532 147420 581588 147476
rect 69692 146972 69748 147028
rect 264684 146972 264740 147028
rect 261212 146860 261268 146916
rect 579740 146860 579796 146916
rect 581420 146300 581476 146356
rect 203196 145180 203252 145236
rect 581644 145180 581700 145236
rect 204092 144732 204148 144788
rect 580412 144620 580468 144676
rect 142828 144060 142884 144116
rect 519260 144060 519316 144116
rect 357196 143724 357252 143780
rect 396620 143724 396676 143780
rect 449372 143724 449428 143780
rect 535164 143724 535220 143780
rect 350364 143612 350420 143668
rect 472892 143612 472948 143668
rect 199164 143500 199220 143556
rect 206668 142940 206724 142996
rect 334348 142940 334404 142996
rect 392252 142716 392308 142772
rect 396956 142716 397012 142772
rect 390572 142604 390628 142660
rect 396732 142604 396788 142660
rect 334460 142492 334516 142548
rect 517692 142492 517748 142548
rect 197484 142156 197540 142212
rect 256172 142044 256228 142100
rect 452732 142044 452788 142100
rect 458892 142044 458948 142100
rect 350252 141932 350308 141988
rect 583436 141932 583492 141988
rect 517580 141820 517636 141876
rect 256172 141708 256228 141764
rect 334460 141708 334516 141764
rect 352044 140812 352100 140868
rect 396844 140812 396900 140868
rect 334348 140588 334404 140644
rect 464492 140588 464548 140644
rect 345436 140364 345492 140420
rect 521052 140364 521108 140420
rect 345212 140252 345268 140308
rect 583324 140252 583380 140308
rect 205772 140140 205828 140196
rect 519372 140140 519428 140196
rect 143612 139804 143668 139860
rect 264012 139804 264068 139860
rect 136892 139692 136948 139748
rect 263900 139692 263956 139748
rect 142044 139580 142100 139636
rect 80332 139468 80388 139524
rect 250236 139468 250292 139524
rect 140924 139356 140980 139412
rect 142828 139356 142884 139412
rect 199276 139132 199332 139188
rect 195804 139020 195860 139076
rect 189084 138572 189140 138628
rect 206668 138572 206724 138628
rect 263788 137900 263844 137956
rect 263900 136780 263956 136836
rect 127484 136668 127540 136724
rect 264012 136220 264068 136276
rect 396508 135324 396564 135380
rect 250236 134540 250292 134596
rect 334460 134540 334516 134596
rect 263900 133980 263956 134036
rect 263788 133420 263844 133476
rect 345212 133420 345268 133476
rect 351932 132860 351988 132916
rect 395836 132636 395892 132692
rect 397068 132636 397124 132692
rect 334460 132300 334516 132356
rect 334348 131740 334404 131796
rect 338492 131180 338548 131236
rect 264684 130620 264740 130676
rect 263788 130060 263844 130116
rect 342188 130060 342244 130116
rect 263900 129500 263956 129556
rect 341852 129276 341908 129332
rect 347788 129276 347844 129332
rect 263900 128940 263956 128996
rect 252924 128492 252980 128548
rect 264572 128492 264628 128548
rect 263788 128380 263844 128436
rect 352604 128380 352660 128436
rect 20076 127932 20132 127988
rect 141036 127932 141092 127988
rect 144060 127932 144116 127988
rect 201628 127932 201684 127988
rect 473676 127932 473732 127988
rect 476028 127932 476084 127988
rect 264012 127820 264068 127876
rect 342636 127820 342692 127876
rect 18396 127260 18452 127316
rect 82684 127260 82740 127316
rect 341964 127260 342020 127316
rect 530796 127260 530852 127316
rect 582988 127260 583044 127316
rect 20636 127148 20692 127204
rect 263788 126700 263844 126756
rect 334460 126700 334516 126756
rect 64876 126588 64932 126644
rect 127260 126588 127316 126644
rect 199052 126588 199108 126644
rect 257852 126588 257908 126644
rect 393260 126588 393316 126644
rect 473004 126588 473060 126644
rect 517468 126588 517524 126644
rect 581644 126588 581700 126644
rect 127372 125916 127428 125972
rect 195692 125916 195748 125972
rect 204876 125916 204932 125972
rect 261324 125916 261380 125972
rect 334460 125580 334516 125636
rect 411628 125916 411684 125972
rect 519372 125916 519428 125972
rect 583436 125916 583492 125972
rect 82460 125468 82516 125524
rect 393372 125468 393428 125524
rect 69692 124572 69748 124628
rect 192332 125244 192388 125300
rect 206108 125244 206164 125300
rect 252812 125244 252868 125300
rect 524972 125244 525028 125300
rect 581532 125244 581588 125300
rect 455420 125132 455476 125188
rect 140812 124572 140868 124628
rect 188972 124572 189028 124628
rect 523292 124572 523348 124628
rect 583212 124572 583268 124628
rect 264796 124460 264852 124516
rect 81452 124012 81508 124068
rect 396732 124012 396788 124068
rect 80332 123900 80388 123956
rect 140924 123900 140980 123956
rect 203084 123900 203140 123956
rect 64204 123228 64260 123284
rect 336812 123340 336868 123396
rect 205772 123228 205828 123284
rect 455308 123900 455364 123956
rect 464492 123900 464548 123956
rect 581308 123900 581364 123956
rect 526652 123228 526708 123284
rect 579628 123228 579684 123284
rect 251916 122780 251972 122836
rect 352268 122780 352324 122836
rect 141036 122668 141092 122724
rect 142044 122668 142100 122724
rect 199164 122668 199220 122724
rect 126924 122556 126980 122612
rect 259980 122556 260036 122612
rect 80444 122444 80500 122500
rect 519260 122556 519316 122612
rect 583324 122556 583380 122612
rect 396844 122444 396900 122500
rect 337036 122220 337092 122276
rect 64764 121884 64820 121940
rect 127148 121884 127204 121940
rect 256396 121884 256452 121940
rect 581420 121884 581476 121940
rect 259532 121660 259588 121716
rect 351820 121660 351876 121716
rect 18172 121212 18228 121268
rect 64988 121212 65044 121268
rect 189084 121212 189140 121268
rect 189532 121212 189588 121268
rect 197484 121212 197540 121268
rect 259756 121212 259812 121268
rect 411180 121212 411236 121268
rect 458780 121212 458836 121268
rect 583100 121212 583156 121268
rect 256172 121100 256228 121156
rect 350252 121100 350308 121156
rect 457772 121100 457828 121156
rect 458668 121100 458724 121156
rect 259980 120876 260036 120932
rect 264684 120876 264740 120932
rect 73836 120540 73892 120596
rect 199276 120540 199332 120596
rect 252812 120540 252868 120596
rect 341852 120540 341908 120596
rect 347788 120540 347844 120596
rect 396620 120540 396676 120596
rect 456988 120540 457044 120596
rect 520828 120540 520884 120596
rect 254492 119980 254548 120036
rect 336924 119980 336980 120036
rect 64204 119868 64260 119924
rect 127036 119868 127092 119924
rect 203196 119868 203252 119924
rect 261212 119868 261268 119924
rect 342188 119868 342244 119924
rect 455308 120316 455364 120372
rect 462812 120092 462868 120148
rect 472108 120092 472164 120148
rect 461356 119868 461412 119924
rect 521052 119868 521108 119924
rect 535164 119868 535220 119924
rect 517692 119756 517748 119812
rect 579740 119756 579796 119812
rect 197372 119308 197428 119364
rect 395724 119308 395780 119364
rect 18396 119196 18452 119252
rect 126812 119196 126868 119252
rect 204092 119196 204148 119252
rect 20076 118524 20132 118580
rect 136892 118524 136948 118580
rect 345324 118860 345380 118916
rect 396508 119196 396564 119252
rect 404012 119196 404068 119252
rect 456092 119196 456148 119252
rect 395612 119084 395668 119140
rect 580412 118860 580468 118916
rect 459004 118524 459060 118580
rect 141932 118412 141988 118468
rect 64652 117852 64708 117908
rect 257852 118300 257908 118356
rect 338716 118300 338772 118356
rect 189532 117852 189588 117908
rect 252924 117852 252980 117908
rect 342636 117852 342692 117908
rect 458892 117852 458948 117908
rect 472108 117852 472164 117908
rect 396508 117404 396564 117460
rect 261436 117292 261492 117348
rect 143612 117180 143668 117236
rect 195804 117180 195860 117236
rect 335244 117180 335300 117236
rect 341964 117180 342020 117236
rect 458668 117180 458724 117236
rect 472892 117180 472948 117236
rect 520940 117180 520996 117236
rect 535052 117180 535108 117236
rect 397068 117068 397124 117124
rect 338604 116620 338660 116676
rect 64204 116508 64260 116564
rect 141036 116508 141092 116564
rect 410844 116508 410900 116564
rect 455644 116508 455700 116564
rect 517580 116508 517636 116564
rect 259644 116060 259700 116116
rect 519148 115836 519204 115892
rect 396956 115724 397012 115780
rect 262892 114492 262948 114548
rect 261436 114380 261492 114436
rect 262892 113820 262948 113876
rect 258076 113260 258132 113316
rect 348684 113260 348740 113316
rect 335132 112700 335188 112756
rect 335468 112140 335524 112196
rect 264684 111580 264740 111636
rect 338492 111580 338548 111636
rect 335356 110460 335412 110516
rect 249452 109900 249508 109956
rect 350364 109900 350420 109956
rect 264124 109340 264180 109396
rect 338940 109340 338996 109396
rect 265132 108780 265188 108836
rect 345436 108780 345492 108836
rect 259756 107100 259812 107156
rect 335916 106540 335972 106596
rect 261324 105980 261380 106036
rect 340396 105980 340452 106036
rect 345548 105420 345604 105476
rect 263788 104860 263844 104916
rect 348572 104860 348628 104916
rect 263900 104300 263956 104356
rect 351148 104300 351204 104356
rect 264012 103740 264068 103796
rect 350476 103740 350532 103796
rect 133532 103292 133588 103348
rect 263788 103292 263844 103348
rect 335244 103292 335300 103348
rect 530012 103292 530068 103348
rect 264572 103180 264628 103236
rect 353612 103180 353668 103236
rect 195692 103068 195748 103124
rect 264124 103068 264180 103124
rect 160860 101724 160916 101780
rect 230188 101724 230244 101780
rect 334460 102060 334516 102116
rect 422044 101948 422100 102004
rect 368172 101836 368228 101892
rect 429436 101836 429492 101892
rect 368844 101724 368900 101780
rect 434140 101724 434196 101780
rect 102844 101612 102900 101668
rect 136892 101612 136948 101668
rect 263900 101612 263956 101668
rect 351148 101612 351204 101668
rect 411068 101612 411124 101668
rect 438844 101612 438900 101668
rect 143612 101500 143668 101556
rect 334572 101500 334628 101556
rect 82012 101052 82068 101108
rect 335468 101052 335524 101108
rect 517468 101052 517524 101108
rect 160860 100940 160916 100996
rect 335244 100940 335300 100996
rect 335916 100828 335972 100884
rect 399196 100828 399252 100884
rect 102844 100716 102900 100772
rect 230188 100716 230244 100772
rect 368172 100716 368228 100772
rect 368844 100716 368900 100772
rect 422044 100716 422100 100772
rect 429436 100716 429492 100772
rect 434140 100716 434196 100772
rect 438844 100716 438900 100772
rect 138572 99932 138628 99988
rect 264012 99932 264068 99988
rect 334460 99932 334516 99988
rect 456988 99932 457044 99988
rect 265020 99820 265076 99876
rect 334348 99820 334404 99876
rect 264796 99260 264852 99316
rect 334684 99260 334740 99316
rect 263788 98700 263844 98756
rect 341964 98700 342020 98756
rect 200956 98252 201012 98308
rect 265132 98252 265188 98308
rect 334348 98252 334404 98308
rect 394828 98252 394884 98308
rect 78092 98140 78148 98196
rect 334460 98140 334516 98196
rect 340172 97580 340228 97636
rect 334460 97132 334516 97188
rect 394940 97132 394996 97188
rect 73052 97020 73108 97076
rect 345212 97020 345268 97076
rect 351932 96796 351988 96852
rect 535164 96796 535220 96852
rect 142716 96684 142772 96740
rect 264684 96684 264740 96740
rect 338716 96572 338772 96628
rect 583436 96572 583492 96628
rect 69692 96460 69748 96516
rect 340284 95900 340340 95956
rect 392252 95340 392308 95396
rect 334572 95004 334628 95060
rect 455308 95004 455364 95060
rect 395612 93660 395668 93716
rect 338940 93324 338996 93380
rect 521276 93324 521332 93380
rect 230188 92540 230244 92596
rect 524972 92540 525028 92596
rect 261212 91980 261268 92036
rect 523292 91980 523348 92036
rect 188972 91868 189028 91924
rect 261436 91868 261492 91924
rect 81452 91644 81508 91700
rect 263788 91644 263844 91700
rect 334684 91644 334740 91700
rect 396956 91644 397012 91700
rect 335356 91532 335412 91588
rect 519148 91532 519204 91588
rect 263788 91420 263844 91476
rect 579628 90860 579684 90916
rect 202860 90188 202916 90244
rect 230188 90188 230244 90244
rect 69804 89852 69860 89908
rect 265020 89852 265076 89908
rect 345436 89852 345492 89908
rect 520940 89852 520996 89908
rect 581308 89740 581364 89796
rect 581420 88620 581476 88676
rect 141932 88284 141988 88340
rect 264572 88284 264628 88340
rect 345548 88284 345604 88340
rect 458668 88284 458724 88340
rect 204876 88060 204932 88116
rect 580412 88060 580468 88116
rect 264908 87500 264964 87556
rect 264572 86940 264628 86996
rect 581532 86940 581588 86996
rect 340396 86604 340452 86660
rect 458780 86604 458836 86660
rect 74732 86492 74788 86548
rect 264796 86492 264852 86548
rect 205772 86380 205828 86436
rect 579740 86380 579796 86436
rect 197372 85820 197428 85876
rect 257964 85708 258020 85764
rect 263788 85708 263844 85764
rect 140588 85260 140644 85316
rect 335244 84924 335300 84980
rect 457100 84924 457156 84980
rect 126812 84812 126868 84868
rect 259756 84812 259812 84868
rect 348684 84812 348740 84868
rect 472892 84812 472948 84868
rect 199052 84140 199108 84196
rect 462812 84140 462868 84196
rect 140924 83580 140980 83636
rect 146972 83020 147028 83076
rect 519260 83020 519316 83076
rect 145292 82460 145348 82516
rect 517580 82460 517636 82516
rect 142044 81340 142100 81396
rect 263788 80780 263844 80836
rect 142604 80220 142660 80276
rect 519372 80220 519428 80276
rect 350476 79884 350532 79940
rect 458892 79884 458948 79940
rect 338604 79772 338660 79828
rect 583100 79772 583156 79828
rect 144060 79660 144116 79716
rect 518252 79660 518308 79716
rect 203084 78316 203140 78372
rect 254492 78316 254548 78372
rect 144284 78204 144340 78260
rect 263788 78204 263844 78260
rect 352268 78204 352324 78260
rect 535388 78204 535444 78260
rect 130172 77980 130228 78036
rect 80220 77420 80276 77476
rect 258188 77308 258244 77364
rect 264908 77308 264964 77364
rect 188076 76860 188132 76916
rect 457772 76860 457828 76916
rect 263788 75740 263844 75796
rect 334460 75740 334516 75796
rect 82348 75180 82404 75236
rect 334348 75180 334404 75236
rect 252924 74732 252980 74788
rect 264572 74732 264628 74788
rect 334460 74732 334516 74788
rect 398076 74620 398132 74676
rect 402332 74620 402388 74676
rect 135212 74060 135268 74116
rect 334572 74060 334628 74116
rect 334460 73500 334516 73556
rect 348572 73500 348628 73556
rect 410732 73500 410788 73556
rect 334348 73388 334404 73444
rect 455420 73388 455476 73444
rect 203196 73276 203252 73332
rect 257852 73276 257908 73332
rect 335132 73276 335188 73332
rect 519484 73276 519540 73332
rect 189084 73164 189140 73220
rect 258076 73164 258132 73220
rect 333452 73164 333508 73220
rect 138684 73052 138740 73108
rect 263788 73052 263844 73108
rect 337036 73052 337092 73108
rect 535276 73052 535332 73108
rect 81564 72940 81620 72996
rect 456092 72940 456148 72996
rect 392252 72156 392308 72212
rect 396620 72156 396676 72212
rect 346892 71820 346948 71876
rect 353612 71708 353668 71764
rect 459116 71708 459172 71764
rect 334460 71596 334516 71652
rect 457212 71596 457268 71652
rect 189420 71484 189476 71540
rect 249452 71484 249508 71540
rect 350252 71484 350308 71540
rect 535500 71484 535556 71540
rect 80332 71372 80388 71428
rect 188076 71372 188132 71428
rect 189196 71372 189252 71428
rect 259644 71372 259700 71428
rect 336924 71372 336980 71428
rect 583212 71372 583268 71428
rect 393932 71260 393988 71316
rect 64652 70700 64708 70756
rect 371196 70700 371252 70756
rect 341852 70476 341908 70532
rect 583324 70476 583380 70532
rect 140812 70364 140868 70420
rect 146972 70364 147028 70420
rect 20636 70140 20692 70196
rect 393148 70140 393204 70196
rect 202972 69916 203028 69972
rect 252812 69916 252868 69972
rect 338492 69916 338548 69972
rect 521052 69916 521108 69972
rect 189308 69804 189364 69860
rect 262892 69804 262948 69860
rect 126924 69692 126980 69748
rect 261324 69692 261380 69748
rect 345324 69804 345380 69860
rect 535612 69804 535668 69860
rect 336812 69692 336868 69748
rect 535836 69692 535892 69748
rect 371196 69132 371252 69188
rect 76412 69020 76468 69076
rect 80444 68796 80500 68852
rect 82348 68796 82404 68852
rect 140700 68796 140756 68852
rect 145292 68796 145348 68852
rect 395052 68572 395108 68628
rect 19964 68460 20020 68516
rect 398076 68236 398132 68292
rect 459004 68236 459060 68292
rect 334572 68124 334628 68180
rect 400652 68124 400708 68180
rect 76524 68012 76580 68068
rect 252812 68012 252868 68068
rect 350364 68012 350420 68068
rect 521164 68012 521220 68068
rect 20076 67900 20132 67956
rect 346780 67900 346836 67956
rect 393148 67900 393204 67956
rect 396732 67900 396788 67956
rect 252812 67788 252868 67844
rect 18284 67228 18340 67284
rect 20636 67228 20692 67284
rect 64764 66332 64820 66388
rect 76412 66332 76468 66388
rect 138572 66220 138628 66276
rect 340284 66220 340340 66276
rect 142716 65548 142772 65604
rect 189420 65548 189476 65604
rect 203196 65548 203252 65604
rect 395052 60396 395108 60452
rect 396844 60396 396900 60452
rect 349356 57036 349412 57092
rect 18396 56812 18452 56868
rect 203196 56812 203252 56868
rect 82572 56252 82628 56308
rect 143612 56252 143668 56308
rect 206108 56252 206164 56308
rect 352604 56252 352660 56308
rect 414652 56252 414708 56308
rect 141036 56140 141092 56196
rect 144060 56140 144116 56196
rect 204876 56140 204932 56196
rect 473676 56140 473732 56196
rect 534268 56140 534324 56196
rect 20076 55468 20132 55524
rect 138684 55468 138740 55524
rect 195692 55468 195748 55524
rect 411068 55468 411124 55524
rect 457100 55468 457156 55524
rect 581420 55468 581476 55524
rect 141932 54796 141988 54852
rect 189308 54796 189364 54852
rect 400652 54796 400708 54852
rect 458668 54796 458724 54852
rect 535836 54796 535892 54852
rect 581532 54796 581588 54852
rect 80332 54124 80388 54180
rect 126924 54124 126980 54180
rect 140812 54124 140868 54180
rect 188972 54124 189028 54180
rect 202860 54124 202916 54180
rect 346780 54124 346836 54180
rect 396956 54124 397012 54180
rect 458780 54124 458836 54180
rect 76412 53452 76468 53508
rect 140700 53452 140756 53508
rect 203084 53452 203140 53508
rect 256172 53452 256228 53508
rect 396732 53452 396788 53508
rect 455308 53452 455364 53508
rect 521164 53452 521220 53508
rect 393932 53228 393988 53284
rect 459116 53228 459172 53284
rect 74732 52780 74788 52836
rect 142604 52780 142660 52836
rect 202972 52780 203028 52836
rect 259532 52780 259588 52836
rect 346892 52780 346948 52836
rect 402332 52780 402388 52836
rect 457772 52892 457828 52948
rect 462812 52780 462868 52836
rect 521052 52780 521108 52836
rect 523292 52780 523348 52836
rect 579628 52780 579684 52836
rect 64764 52108 64820 52164
rect 189196 52108 189252 52164
rect 261212 52108 261268 52164
rect 341964 52108 342020 52164
rect 410732 52108 410788 52164
rect 517580 52108 517636 52164
rect 535388 52108 535444 52164
rect 583324 52108 583380 52164
rect 395612 51996 395668 52052
rect 396508 51996 396564 52052
rect 64652 51436 64708 51492
rect 456988 51436 457044 51492
rect 520940 51436 520996 51492
rect 64316 51324 64372 51380
rect 73052 51324 73108 51380
rect 64092 51212 64148 51268
rect 78092 51212 78148 51268
rect 126812 50764 126868 50820
rect 457212 50764 457268 50820
rect 519148 50764 519204 50820
rect 524972 50764 525028 50820
rect 579740 50764 579796 50820
rect 127596 50540 127652 50596
rect 130172 50540 130228 50596
rect 81452 50204 81508 50260
rect 81564 50092 81620 50148
rect 136892 50092 136948 50148
rect 144284 50092 144340 50148
rect 200956 50092 201012 50148
rect 257964 50092 258020 50148
rect 394940 50092 394996 50148
rect 458892 50092 458948 50148
rect 133532 49420 133588 49476
rect 144060 49420 144116 49476
rect 189084 49420 189140 49476
rect 251916 49420 251972 49476
rect 340172 49420 340228 49476
rect 459004 49420 459060 49476
rect 535612 49420 535668 49476
rect 583212 49420 583268 49476
rect 142044 49196 142100 49252
rect 64316 48748 64372 48804
rect 519372 48748 519428 48804
rect 530012 48748 530068 48804
rect 64204 48636 64260 48692
rect 69692 48636 69748 48692
rect 189532 48636 189588 48692
rect 199052 48636 199108 48692
rect 19964 48188 20020 48244
rect 64092 48076 64148 48132
rect 394828 48076 394884 48132
rect 399196 48076 399252 48132
rect 455420 48076 455476 48132
rect 519260 48076 519316 48132
rect 535164 48076 535220 48132
rect 518252 47852 518308 47908
rect 456092 47516 456148 47572
rect 82012 47404 82068 47460
rect 197372 47404 197428 47460
rect 258188 47404 258244 47460
rect 345212 47404 345268 47460
rect 135212 47068 135268 47124
rect 80444 46732 80500 46788
rect 581308 47404 581364 47460
rect 580412 47068 580468 47124
rect 80220 46060 80276 46116
rect 127596 46060 127652 46116
rect 140588 46060 140644 46116
rect 189532 46060 189588 46116
rect 396620 46060 396676 46116
rect 535276 46060 535332 46116
rect 205772 45948 205828 46004
rect 18284 45388 18340 45444
rect 64204 45388 64260 45444
rect 140924 45388 140980 45444
rect 252924 45388 252980 45444
rect 396844 45388 396900 45444
rect 535500 45388 535556 45444
rect 583436 45388 583492 45444
rect 69804 44716 69860 44772
rect 396508 44716 396564 44772
rect 472892 44716 472948 44772
rect 517468 44716 517524 44772
rect 583100 44716 583156 44772
rect 519484 44044 519540 44100
rect 521276 43372 521332 43428
rect 585452 33740 585508 33796
rect 270060 29932 270116 29988
rect 200844 8540 200900 8596
rect 18396 5068 18452 5124
<< metal4 >>
rect -1916 598172 -1296 598268
rect -1916 598116 -1820 598172
rect -1764 598116 -1696 598172
rect -1640 598116 -1572 598172
rect -1516 598116 -1448 598172
rect -1392 598116 -1296 598172
rect -1916 598048 -1296 598116
rect -1916 597992 -1820 598048
rect -1764 597992 -1696 598048
rect -1640 597992 -1572 598048
rect -1516 597992 -1448 598048
rect -1392 597992 -1296 598048
rect -1916 597924 -1296 597992
rect -1916 597868 -1820 597924
rect -1764 597868 -1696 597924
rect -1640 597868 -1572 597924
rect -1516 597868 -1448 597924
rect -1392 597868 -1296 597924
rect -1916 597800 -1296 597868
rect -1916 597744 -1820 597800
rect -1764 597744 -1696 597800
rect -1640 597744 -1572 597800
rect -1516 597744 -1448 597800
rect -1392 597744 -1296 597800
rect -1916 586350 -1296 597744
rect -1916 586294 -1820 586350
rect -1764 586294 -1696 586350
rect -1640 586294 -1572 586350
rect -1516 586294 -1448 586350
rect -1392 586294 -1296 586350
rect -1916 586226 -1296 586294
rect -1916 586170 -1820 586226
rect -1764 586170 -1696 586226
rect -1640 586170 -1572 586226
rect -1516 586170 -1448 586226
rect -1392 586170 -1296 586226
rect -1916 586102 -1296 586170
rect -1916 586046 -1820 586102
rect -1764 586046 -1696 586102
rect -1640 586046 -1572 586102
rect -1516 586046 -1448 586102
rect -1392 586046 -1296 586102
rect -1916 585978 -1296 586046
rect -1916 585922 -1820 585978
rect -1764 585922 -1696 585978
rect -1640 585922 -1572 585978
rect -1516 585922 -1448 585978
rect -1392 585922 -1296 585978
rect -1916 568350 -1296 585922
rect -1916 568294 -1820 568350
rect -1764 568294 -1696 568350
rect -1640 568294 -1572 568350
rect -1516 568294 -1448 568350
rect -1392 568294 -1296 568350
rect -1916 568226 -1296 568294
rect -1916 568170 -1820 568226
rect -1764 568170 -1696 568226
rect -1640 568170 -1572 568226
rect -1516 568170 -1448 568226
rect -1392 568170 -1296 568226
rect -1916 568102 -1296 568170
rect -1916 568046 -1820 568102
rect -1764 568046 -1696 568102
rect -1640 568046 -1572 568102
rect -1516 568046 -1448 568102
rect -1392 568046 -1296 568102
rect -1916 567978 -1296 568046
rect -1916 567922 -1820 567978
rect -1764 567922 -1696 567978
rect -1640 567922 -1572 567978
rect -1516 567922 -1448 567978
rect -1392 567922 -1296 567978
rect -1916 550350 -1296 567922
rect -1916 550294 -1820 550350
rect -1764 550294 -1696 550350
rect -1640 550294 -1572 550350
rect -1516 550294 -1448 550350
rect -1392 550294 -1296 550350
rect -1916 550226 -1296 550294
rect -1916 550170 -1820 550226
rect -1764 550170 -1696 550226
rect -1640 550170 -1572 550226
rect -1516 550170 -1448 550226
rect -1392 550170 -1296 550226
rect -1916 550102 -1296 550170
rect -1916 550046 -1820 550102
rect -1764 550046 -1696 550102
rect -1640 550046 -1572 550102
rect -1516 550046 -1448 550102
rect -1392 550046 -1296 550102
rect -1916 549978 -1296 550046
rect -1916 549922 -1820 549978
rect -1764 549922 -1696 549978
rect -1640 549922 -1572 549978
rect -1516 549922 -1448 549978
rect -1392 549922 -1296 549978
rect -1916 532350 -1296 549922
rect -1916 532294 -1820 532350
rect -1764 532294 -1696 532350
rect -1640 532294 -1572 532350
rect -1516 532294 -1448 532350
rect -1392 532294 -1296 532350
rect -1916 532226 -1296 532294
rect -1916 532170 -1820 532226
rect -1764 532170 -1696 532226
rect -1640 532170 -1572 532226
rect -1516 532170 -1448 532226
rect -1392 532170 -1296 532226
rect -1916 532102 -1296 532170
rect -1916 532046 -1820 532102
rect -1764 532046 -1696 532102
rect -1640 532046 -1572 532102
rect -1516 532046 -1448 532102
rect -1392 532046 -1296 532102
rect -1916 531978 -1296 532046
rect -1916 531922 -1820 531978
rect -1764 531922 -1696 531978
rect -1640 531922 -1572 531978
rect -1516 531922 -1448 531978
rect -1392 531922 -1296 531978
rect -1916 514350 -1296 531922
rect -1916 514294 -1820 514350
rect -1764 514294 -1696 514350
rect -1640 514294 -1572 514350
rect -1516 514294 -1448 514350
rect -1392 514294 -1296 514350
rect -1916 514226 -1296 514294
rect -1916 514170 -1820 514226
rect -1764 514170 -1696 514226
rect -1640 514170 -1572 514226
rect -1516 514170 -1448 514226
rect -1392 514170 -1296 514226
rect -1916 514102 -1296 514170
rect -1916 514046 -1820 514102
rect -1764 514046 -1696 514102
rect -1640 514046 -1572 514102
rect -1516 514046 -1448 514102
rect -1392 514046 -1296 514102
rect -1916 513978 -1296 514046
rect -1916 513922 -1820 513978
rect -1764 513922 -1696 513978
rect -1640 513922 -1572 513978
rect -1516 513922 -1448 513978
rect -1392 513922 -1296 513978
rect -1916 496350 -1296 513922
rect -1916 496294 -1820 496350
rect -1764 496294 -1696 496350
rect -1640 496294 -1572 496350
rect -1516 496294 -1448 496350
rect -1392 496294 -1296 496350
rect -1916 496226 -1296 496294
rect -1916 496170 -1820 496226
rect -1764 496170 -1696 496226
rect -1640 496170 -1572 496226
rect -1516 496170 -1448 496226
rect -1392 496170 -1296 496226
rect -1916 496102 -1296 496170
rect -1916 496046 -1820 496102
rect -1764 496046 -1696 496102
rect -1640 496046 -1572 496102
rect -1516 496046 -1448 496102
rect -1392 496046 -1296 496102
rect -1916 495978 -1296 496046
rect -1916 495922 -1820 495978
rect -1764 495922 -1696 495978
rect -1640 495922 -1572 495978
rect -1516 495922 -1448 495978
rect -1392 495922 -1296 495978
rect -1916 478350 -1296 495922
rect -1916 478294 -1820 478350
rect -1764 478294 -1696 478350
rect -1640 478294 -1572 478350
rect -1516 478294 -1448 478350
rect -1392 478294 -1296 478350
rect -1916 478226 -1296 478294
rect -1916 478170 -1820 478226
rect -1764 478170 -1696 478226
rect -1640 478170 -1572 478226
rect -1516 478170 -1448 478226
rect -1392 478170 -1296 478226
rect -1916 478102 -1296 478170
rect -1916 478046 -1820 478102
rect -1764 478046 -1696 478102
rect -1640 478046 -1572 478102
rect -1516 478046 -1448 478102
rect -1392 478046 -1296 478102
rect -1916 477978 -1296 478046
rect -1916 477922 -1820 477978
rect -1764 477922 -1696 477978
rect -1640 477922 -1572 477978
rect -1516 477922 -1448 477978
rect -1392 477922 -1296 477978
rect -1916 460350 -1296 477922
rect -1916 460294 -1820 460350
rect -1764 460294 -1696 460350
rect -1640 460294 -1572 460350
rect -1516 460294 -1448 460350
rect -1392 460294 -1296 460350
rect -1916 460226 -1296 460294
rect -1916 460170 -1820 460226
rect -1764 460170 -1696 460226
rect -1640 460170 -1572 460226
rect -1516 460170 -1448 460226
rect -1392 460170 -1296 460226
rect -1916 460102 -1296 460170
rect -1916 460046 -1820 460102
rect -1764 460046 -1696 460102
rect -1640 460046 -1572 460102
rect -1516 460046 -1448 460102
rect -1392 460046 -1296 460102
rect -1916 459978 -1296 460046
rect -1916 459922 -1820 459978
rect -1764 459922 -1696 459978
rect -1640 459922 -1572 459978
rect -1516 459922 -1448 459978
rect -1392 459922 -1296 459978
rect -1916 442350 -1296 459922
rect -1916 442294 -1820 442350
rect -1764 442294 -1696 442350
rect -1640 442294 -1572 442350
rect -1516 442294 -1448 442350
rect -1392 442294 -1296 442350
rect -1916 442226 -1296 442294
rect -1916 442170 -1820 442226
rect -1764 442170 -1696 442226
rect -1640 442170 -1572 442226
rect -1516 442170 -1448 442226
rect -1392 442170 -1296 442226
rect -1916 442102 -1296 442170
rect -1916 442046 -1820 442102
rect -1764 442046 -1696 442102
rect -1640 442046 -1572 442102
rect -1516 442046 -1448 442102
rect -1392 442046 -1296 442102
rect -1916 441978 -1296 442046
rect -1916 441922 -1820 441978
rect -1764 441922 -1696 441978
rect -1640 441922 -1572 441978
rect -1516 441922 -1448 441978
rect -1392 441922 -1296 441978
rect -1916 424350 -1296 441922
rect -1916 424294 -1820 424350
rect -1764 424294 -1696 424350
rect -1640 424294 -1572 424350
rect -1516 424294 -1448 424350
rect -1392 424294 -1296 424350
rect -1916 424226 -1296 424294
rect -1916 424170 -1820 424226
rect -1764 424170 -1696 424226
rect -1640 424170 -1572 424226
rect -1516 424170 -1448 424226
rect -1392 424170 -1296 424226
rect -1916 424102 -1296 424170
rect -1916 424046 -1820 424102
rect -1764 424046 -1696 424102
rect -1640 424046 -1572 424102
rect -1516 424046 -1448 424102
rect -1392 424046 -1296 424102
rect -1916 423978 -1296 424046
rect -1916 423922 -1820 423978
rect -1764 423922 -1696 423978
rect -1640 423922 -1572 423978
rect -1516 423922 -1448 423978
rect -1392 423922 -1296 423978
rect -1916 406350 -1296 423922
rect -1916 406294 -1820 406350
rect -1764 406294 -1696 406350
rect -1640 406294 -1572 406350
rect -1516 406294 -1448 406350
rect -1392 406294 -1296 406350
rect -1916 406226 -1296 406294
rect -1916 406170 -1820 406226
rect -1764 406170 -1696 406226
rect -1640 406170 -1572 406226
rect -1516 406170 -1448 406226
rect -1392 406170 -1296 406226
rect -1916 406102 -1296 406170
rect -1916 406046 -1820 406102
rect -1764 406046 -1696 406102
rect -1640 406046 -1572 406102
rect -1516 406046 -1448 406102
rect -1392 406046 -1296 406102
rect -1916 405978 -1296 406046
rect -1916 405922 -1820 405978
rect -1764 405922 -1696 405978
rect -1640 405922 -1572 405978
rect -1516 405922 -1448 405978
rect -1392 405922 -1296 405978
rect -1916 388350 -1296 405922
rect -1916 388294 -1820 388350
rect -1764 388294 -1696 388350
rect -1640 388294 -1572 388350
rect -1516 388294 -1448 388350
rect -1392 388294 -1296 388350
rect -1916 388226 -1296 388294
rect -1916 388170 -1820 388226
rect -1764 388170 -1696 388226
rect -1640 388170 -1572 388226
rect -1516 388170 -1448 388226
rect -1392 388170 -1296 388226
rect -1916 388102 -1296 388170
rect -1916 388046 -1820 388102
rect -1764 388046 -1696 388102
rect -1640 388046 -1572 388102
rect -1516 388046 -1448 388102
rect -1392 388046 -1296 388102
rect -1916 387978 -1296 388046
rect -1916 387922 -1820 387978
rect -1764 387922 -1696 387978
rect -1640 387922 -1572 387978
rect -1516 387922 -1448 387978
rect -1392 387922 -1296 387978
rect -1916 370350 -1296 387922
rect -1916 370294 -1820 370350
rect -1764 370294 -1696 370350
rect -1640 370294 -1572 370350
rect -1516 370294 -1448 370350
rect -1392 370294 -1296 370350
rect -1916 370226 -1296 370294
rect -1916 370170 -1820 370226
rect -1764 370170 -1696 370226
rect -1640 370170 -1572 370226
rect -1516 370170 -1448 370226
rect -1392 370170 -1296 370226
rect -1916 370102 -1296 370170
rect -1916 370046 -1820 370102
rect -1764 370046 -1696 370102
rect -1640 370046 -1572 370102
rect -1516 370046 -1448 370102
rect -1392 370046 -1296 370102
rect -1916 369978 -1296 370046
rect -1916 369922 -1820 369978
rect -1764 369922 -1696 369978
rect -1640 369922 -1572 369978
rect -1516 369922 -1448 369978
rect -1392 369922 -1296 369978
rect -1916 352350 -1296 369922
rect -1916 352294 -1820 352350
rect -1764 352294 -1696 352350
rect -1640 352294 -1572 352350
rect -1516 352294 -1448 352350
rect -1392 352294 -1296 352350
rect -1916 352226 -1296 352294
rect -1916 352170 -1820 352226
rect -1764 352170 -1696 352226
rect -1640 352170 -1572 352226
rect -1516 352170 -1448 352226
rect -1392 352170 -1296 352226
rect -1916 352102 -1296 352170
rect -1916 352046 -1820 352102
rect -1764 352046 -1696 352102
rect -1640 352046 -1572 352102
rect -1516 352046 -1448 352102
rect -1392 352046 -1296 352102
rect -1916 351978 -1296 352046
rect -1916 351922 -1820 351978
rect -1764 351922 -1696 351978
rect -1640 351922 -1572 351978
rect -1516 351922 -1448 351978
rect -1392 351922 -1296 351978
rect -1916 334350 -1296 351922
rect -1916 334294 -1820 334350
rect -1764 334294 -1696 334350
rect -1640 334294 -1572 334350
rect -1516 334294 -1448 334350
rect -1392 334294 -1296 334350
rect -1916 334226 -1296 334294
rect -1916 334170 -1820 334226
rect -1764 334170 -1696 334226
rect -1640 334170 -1572 334226
rect -1516 334170 -1448 334226
rect -1392 334170 -1296 334226
rect -1916 334102 -1296 334170
rect -1916 334046 -1820 334102
rect -1764 334046 -1696 334102
rect -1640 334046 -1572 334102
rect -1516 334046 -1448 334102
rect -1392 334046 -1296 334102
rect -1916 333978 -1296 334046
rect -1916 333922 -1820 333978
rect -1764 333922 -1696 333978
rect -1640 333922 -1572 333978
rect -1516 333922 -1448 333978
rect -1392 333922 -1296 333978
rect -1916 316350 -1296 333922
rect -1916 316294 -1820 316350
rect -1764 316294 -1696 316350
rect -1640 316294 -1572 316350
rect -1516 316294 -1448 316350
rect -1392 316294 -1296 316350
rect -1916 316226 -1296 316294
rect -1916 316170 -1820 316226
rect -1764 316170 -1696 316226
rect -1640 316170 -1572 316226
rect -1516 316170 -1448 316226
rect -1392 316170 -1296 316226
rect -1916 316102 -1296 316170
rect -1916 316046 -1820 316102
rect -1764 316046 -1696 316102
rect -1640 316046 -1572 316102
rect -1516 316046 -1448 316102
rect -1392 316046 -1296 316102
rect -1916 315978 -1296 316046
rect -1916 315922 -1820 315978
rect -1764 315922 -1696 315978
rect -1640 315922 -1572 315978
rect -1516 315922 -1448 315978
rect -1392 315922 -1296 315978
rect -1916 298350 -1296 315922
rect -1916 298294 -1820 298350
rect -1764 298294 -1696 298350
rect -1640 298294 -1572 298350
rect -1516 298294 -1448 298350
rect -1392 298294 -1296 298350
rect -1916 298226 -1296 298294
rect -1916 298170 -1820 298226
rect -1764 298170 -1696 298226
rect -1640 298170 -1572 298226
rect -1516 298170 -1448 298226
rect -1392 298170 -1296 298226
rect -1916 298102 -1296 298170
rect -1916 298046 -1820 298102
rect -1764 298046 -1696 298102
rect -1640 298046 -1572 298102
rect -1516 298046 -1448 298102
rect -1392 298046 -1296 298102
rect -1916 297978 -1296 298046
rect -1916 297922 -1820 297978
rect -1764 297922 -1696 297978
rect -1640 297922 -1572 297978
rect -1516 297922 -1448 297978
rect -1392 297922 -1296 297978
rect -1916 280350 -1296 297922
rect -1916 280294 -1820 280350
rect -1764 280294 -1696 280350
rect -1640 280294 -1572 280350
rect -1516 280294 -1448 280350
rect -1392 280294 -1296 280350
rect -1916 280226 -1296 280294
rect -1916 280170 -1820 280226
rect -1764 280170 -1696 280226
rect -1640 280170 -1572 280226
rect -1516 280170 -1448 280226
rect -1392 280170 -1296 280226
rect -1916 280102 -1296 280170
rect -1916 280046 -1820 280102
rect -1764 280046 -1696 280102
rect -1640 280046 -1572 280102
rect -1516 280046 -1448 280102
rect -1392 280046 -1296 280102
rect -1916 279978 -1296 280046
rect -1916 279922 -1820 279978
rect -1764 279922 -1696 279978
rect -1640 279922 -1572 279978
rect -1516 279922 -1448 279978
rect -1392 279922 -1296 279978
rect -1916 262350 -1296 279922
rect -1916 262294 -1820 262350
rect -1764 262294 -1696 262350
rect -1640 262294 -1572 262350
rect -1516 262294 -1448 262350
rect -1392 262294 -1296 262350
rect -1916 262226 -1296 262294
rect -1916 262170 -1820 262226
rect -1764 262170 -1696 262226
rect -1640 262170 -1572 262226
rect -1516 262170 -1448 262226
rect -1392 262170 -1296 262226
rect -1916 262102 -1296 262170
rect -1916 262046 -1820 262102
rect -1764 262046 -1696 262102
rect -1640 262046 -1572 262102
rect -1516 262046 -1448 262102
rect -1392 262046 -1296 262102
rect -1916 261978 -1296 262046
rect -1916 261922 -1820 261978
rect -1764 261922 -1696 261978
rect -1640 261922 -1572 261978
rect -1516 261922 -1448 261978
rect -1392 261922 -1296 261978
rect -1916 244350 -1296 261922
rect -1916 244294 -1820 244350
rect -1764 244294 -1696 244350
rect -1640 244294 -1572 244350
rect -1516 244294 -1448 244350
rect -1392 244294 -1296 244350
rect -1916 244226 -1296 244294
rect -1916 244170 -1820 244226
rect -1764 244170 -1696 244226
rect -1640 244170 -1572 244226
rect -1516 244170 -1448 244226
rect -1392 244170 -1296 244226
rect -1916 244102 -1296 244170
rect -1916 244046 -1820 244102
rect -1764 244046 -1696 244102
rect -1640 244046 -1572 244102
rect -1516 244046 -1448 244102
rect -1392 244046 -1296 244102
rect -1916 243978 -1296 244046
rect -1916 243922 -1820 243978
rect -1764 243922 -1696 243978
rect -1640 243922 -1572 243978
rect -1516 243922 -1448 243978
rect -1392 243922 -1296 243978
rect -1916 226350 -1296 243922
rect -1916 226294 -1820 226350
rect -1764 226294 -1696 226350
rect -1640 226294 -1572 226350
rect -1516 226294 -1448 226350
rect -1392 226294 -1296 226350
rect -1916 226226 -1296 226294
rect -1916 226170 -1820 226226
rect -1764 226170 -1696 226226
rect -1640 226170 -1572 226226
rect -1516 226170 -1448 226226
rect -1392 226170 -1296 226226
rect -1916 226102 -1296 226170
rect -1916 226046 -1820 226102
rect -1764 226046 -1696 226102
rect -1640 226046 -1572 226102
rect -1516 226046 -1448 226102
rect -1392 226046 -1296 226102
rect -1916 225978 -1296 226046
rect -1916 225922 -1820 225978
rect -1764 225922 -1696 225978
rect -1640 225922 -1572 225978
rect -1516 225922 -1448 225978
rect -1392 225922 -1296 225978
rect -1916 208350 -1296 225922
rect -1916 208294 -1820 208350
rect -1764 208294 -1696 208350
rect -1640 208294 -1572 208350
rect -1516 208294 -1448 208350
rect -1392 208294 -1296 208350
rect -1916 208226 -1296 208294
rect -1916 208170 -1820 208226
rect -1764 208170 -1696 208226
rect -1640 208170 -1572 208226
rect -1516 208170 -1448 208226
rect -1392 208170 -1296 208226
rect -1916 208102 -1296 208170
rect -1916 208046 -1820 208102
rect -1764 208046 -1696 208102
rect -1640 208046 -1572 208102
rect -1516 208046 -1448 208102
rect -1392 208046 -1296 208102
rect -1916 207978 -1296 208046
rect -1916 207922 -1820 207978
rect -1764 207922 -1696 207978
rect -1640 207922 -1572 207978
rect -1516 207922 -1448 207978
rect -1392 207922 -1296 207978
rect -1916 190350 -1296 207922
rect -1916 190294 -1820 190350
rect -1764 190294 -1696 190350
rect -1640 190294 -1572 190350
rect -1516 190294 -1448 190350
rect -1392 190294 -1296 190350
rect -1916 190226 -1296 190294
rect -1916 190170 -1820 190226
rect -1764 190170 -1696 190226
rect -1640 190170 -1572 190226
rect -1516 190170 -1448 190226
rect -1392 190170 -1296 190226
rect -1916 190102 -1296 190170
rect -1916 190046 -1820 190102
rect -1764 190046 -1696 190102
rect -1640 190046 -1572 190102
rect -1516 190046 -1448 190102
rect -1392 190046 -1296 190102
rect -1916 189978 -1296 190046
rect -1916 189922 -1820 189978
rect -1764 189922 -1696 189978
rect -1640 189922 -1572 189978
rect -1516 189922 -1448 189978
rect -1392 189922 -1296 189978
rect -1916 172350 -1296 189922
rect -1916 172294 -1820 172350
rect -1764 172294 -1696 172350
rect -1640 172294 -1572 172350
rect -1516 172294 -1448 172350
rect -1392 172294 -1296 172350
rect -1916 172226 -1296 172294
rect -1916 172170 -1820 172226
rect -1764 172170 -1696 172226
rect -1640 172170 -1572 172226
rect -1516 172170 -1448 172226
rect -1392 172170 -1296 172226
rect -1916 172102 -1296 172170
rect -1916 172046 -1820 172102
rect -1764 172046 -1696 172102
rect -1640 172046 -1572 172102
rect -1516 172046 -1448 172102
rect -1392 172046 -1296 172102
rect -1916 171978 -1296 172046
rect -1916 171922 -1820 171978
rect -1764 171922 -1696 171978
rect -1640 171922 -1572 171978
rect -1516 171922 -1448 171978
rect -1392 171922 -1296 171978
rect -1916 154350 -1296 171922
rect -1916 154294 -1820 154350
rect -1764 154294 -1696 154350
rect -1640 154294 -1572 154350
rect -1516 154294 -1448 154350
rect -1392 154294 -1296 154350
rect -1916 154226 -1296 154294
rect -1916 154170 -1820 154226
rect -1764 154170 -1696 154226
rect -1640 154170 -1572 154226
rect -1516 154170 -1448 154226
rect -1392 154170 -1296 154226
rect -1916 154102 -1296 154170
rect -1916 154046 -1820 154102
rect -1764 154046 -1696 154102
rect -1640 154046 -1572 154102
rect -1516 154046 -1448 154102
rect -1392 154046 -1296 154102
rect -1916 153978 -1296 154046
rect -1916 153922 -1820 153978
rect -1764 153922 -1696 153978
rect -1640 153922 -1572 153978
rect -1516 153922 -1448 153978
rect -1392 153922 -1296 153978
rect -1916 136350 -1296 153922
rect -1916 136294 -1820 136350
rect -1764 136294 -1696 136350
rect -1640 136294 -1572 136350
rect -1516 136294 -1448 136350
rect -1392 136294 -1296 136350
rect -1916 136226 -1296 136294
rect -1916 136170 -1820 136226
rect -1764 136170 -1696 136226
rect -1640 136170 -1572 136226
rect -1516 136170 -1448 136226
rect -1392 136170 -1296 136226
rect -1916 136102 -1296 136170
rect -1916 136046 -1820 136102
rect -1764 136046 -1696 136102
rect -1640 136046 -1572 136102
rect -1516 136046 -1448 136102
rect -1392 136046 -1296 136102
rect -1916 135978 -1296 136046
rect -1916 135922 -1820 135978
rect -1764 135922 -1696 135978
rect -1640 135922 -1572 135978
rect -1516 135922 -1448 135978
rect -1392 135922 -1296 135978
rect -1916 118350 -1296 135922
rect -1916 118294 -1820 118350
rect -1764 118294 -1696 118350
rect -1640 118294 -1572 118350
rect -1516 118294 -1448 118350
rect -1392 118294 -1296 118350
rect -1916 118226 -1296 118294
rect -1916 118170 -1820 118226
rect -1764 118170 -1696 118226
rect -1640 118170 -1572 118226
rect -1516 118170 -1448 118226
rect -1392 118170 -1296 118226
rect -1916 118102 -1296 118170
rect -1916 118046 -1820 118102
rect -1764 118046 -1696 118102
rect -1640 118046 -1572 118102
rect -1516 118046 -1448 118102
rect -1392 118046 -1296 118102
rect -1916 117978 -1296 118046
rect -1916 117922 -1820 117978
rect -1764 117922 -1696 117978
rect -1640 117922 -1572 117978
rect -1516 117922 -1448 117978
rect -1392 117922 -1296 117978
rect -1916 100350 -1296 117922
rect -1916 100294 -1820 100350
rect -1764 100294 -1696 100350
rect -1640 100294 -1572 100350
rect -1516 100294 -1448 100350
rect -1392 100294 -1296 100350
rect -1916 100226 -1296 100294
rect -1916 100170 -1820 100226
rect -1764 100170 -1696 100226
rect -1640 100170 -1572 100226
rect -1516 100170 -1448 100226
rect -1392 100170 -1296 100226
rect -1916 100102 -1296 100170
rect -1916 100046 -1820 100102
rect -1764 100046 -1696 100102
rect -1640 100046 -1572 100102
rect -1516 100046 -1448 100102
rect -1392 100046 -1296 100102
rect -1916 99978 -1296 100046
rect -1916 99922 -1820 99978
rect -1764 99922 -1696 99978
rect -1640 99922 -1572 99978
rect -1516 99922 -1448 99978
rect -1392 99922 -1296 99978
rect -1916 82350 -1296 99922
rect -1916 82294 -1820 82350
rect -1764 82294 -1696 82350
rect -1640 82294 -1572 82350
rect -1516 82294 -1448 82350
rect -1392 82294 -1296 82350
rect -1916 82226 -1296 82294
rect -1916 82170 -1820 82226
rect -1764 82170 -1696 82226
rect -1640 82170 -1572 82226
rect -1516 82170 -1448 82226
rect -1392 82170 -1296 82226
rect -1916 82102 -1296 82170
rect -1916 82046 -1820 82102
rect -1764 82046 -1696 82102
rect -1640 82046 -1572 82102
rect -1516 82046 -1448 82102
rect -1392 82046 -1296 82102
rect -1916 81978 -1296 82046
rect -1916 81922 -1820 81978
rect -1764 81922 -1696 81978
rect -1640 81922 -1572 81978
rect -1516 81922 -1448 81978
rect -1392 81922 -1296 81978
rect -1916 64350 -1296 81922
rect -1916 64294 -1820 64350
rect -1764 64294 -1696 64350
rect -1640 64294 -1572 64350
rect -1516 64294 -1448 64350
rect -1392 64294 -1296 64350
rect -1916 64226 -1296 64294
rect -1916 64170 -1820 64226
rect -1764 64170 -1696 64226
rect -1640 64170 -1572 64226
rect -1516 64170 -1448 64226
rect -1392 64170 -1296 64226
rect -1916 64102 -1296 64170
rect -1916 64046 -1820 64102
rect -1764 64046 -1696 64102
rect -1640 64046 -1572 64102
rect -1516 64046 -1448 64102
rect -1392 64046 -1296 64102
rect -1916 63978 -1296 64046
rect -1916 63922 -1820 63978
rect -1764 63922 -1696 63978
rect -1640 63922 -1572 63978
rect -1516 63922 -1448 63978
rect -1392 63922 -1296 63978
rect -1916 46350 -1296 63922
rect -1916 46294 -1820 46350
rect -1764 46294 -1696 46350
rect -1640 46294 -1572 46350
rect -1516 46294 -1448 46350
rect -1392 46294 -1296 46350
rect -1916 46226 -1296 46294
rect -1916 46170 -1820 46226
rect -1764 46170 -1696 46226
rect -1640 46170 -1572 46226
rect -1516 46170 -1448 46226
rect -1392 46170 -1296 46226
rect -1916 46102 -1296 46170
rect -1916 46046 -1820 46102
rect -1764 46046 -1696 46102
rect -1640 46046 -1572 46102
rect -1516 46046 -1448 46102
rect -1392 46046 -1296 46102
rect -1916 45978 -1296 46046
rect -1916 45922 -1820 45978
rect -1764 45922 -1696 45978
rect -1640 45922 -1572 45978
rect -1516 45922 -1448 45978
rect -1392 45922 -1296 45978
rect -1916 28350 -1296 45922
rect -1916 28294 -1820 28350
rect -1764 28294 -1696 28350
rect -1640 28294 -1572 28350
rect -1516 28294 -1448 28350
rect -1392 28294 -1296 28350
rect -1916 28226 -1296 28294
rect -1916 28170 -1820 28226
rect -1764 28170 -1696 28226
rect -1640 28170 -1572 28226
rect -1516 28170 -1448 28226
rect -1392 28170 -1296 28226
rect -1916 28102 -1296 28170
rect -1916 28046 -1820 28102
rect -1764 28046 -1696 28102
rect -1640 28046 -1572 28102
rect -1516 28046 -1448 28102
rect -1392 28046 -1296 28102
rect -1916 27978 -1296 28046
rect -1916 27922 -1820 27978
rect -1764 27922 -1696 27978
rect -1640 27922 -1572 27978
rect -1516 27922 -1448 27978
rect -1392 27922 -1296 27978
rect -1916 10350 -1296 27922
rect -1916 10294 -1820 10350
rect -1764 10294 -1696 10350
rect -1640 10294 -1572 10350
rect -1516 10294 -1448 10350
rect -1392 10294 -1296 10350
rect -1916 10226 -1296 10294
rect -1916 10170 -1820 10226
rect -1764 10170 -1696 10226
rect -1640 10170 -1572 10226
rect -1516 10170 -1448 10226
rect -1392 10170 -1296 10226
rect -1916 10102 -1296 10170
rect -1916 10046 -1820 10102
rect -1764 10046 -1696 10102
rect -1640 10046 -1572 10102
rect -1516 10046 -1448 10102
rect -1392 10046 -1296 10102
rect -1916 9978 -1296 10046
rect -1916 9922 -1820 9978
rect -1764 9922 -1696 9978
rect -1640 9922 -1572 9978
rect -1516 9922 -1448 9978
rect -1392 9922 -1296 9978
rect -1916 -1120 -1296 9922
rect -956 597212 -336 597308
rect -956 597156 -860 597212
rect -804 597156 -736 597212
rect -680 597156 -612 597212
rect -556 597156 -488 597212
rect -432 597156 -336 597212
rect -956 597088 -336 597156
rect -956 597032 -860 597088
rect -804 597032 -736 597088
rect -680 597032 -612 597088
rect -556 597032 -488 597088
rect -432 597032 -336 597088
rect -956 596964 -336 597032
rect -956 596908 -860 596964
rect -804 596908 -736 596964
rect -680 596908 -612 596964
rect -556 596908 -488 596964
rect -432 596908 -336 596964
rect -956 596840 -336 596908
rect -956 596784 -860 596840
rect -804 596784 -736 596840
rect -680 596784 -612 596840
rect -556 596784 -488 596840
rect -432 596784 -336 596840
rect -956 580350 -336 596784
rect -956 580294 -860 580350
rect -804 580294 -736 580350
rect -680 580294 -612 580350
rect -556 580294 -488 580350
rect -432 580294 -336 580350
rect -956 580226 -336 580294
rect -956 580170 -860 580226
rect -804 580170 -736 580226
rect -680 580170 -612 580226
rect -556 580170 -488 580226
rect -432 580170 -336 580226
rect -956 580102 -336 580170
rect -956 580046 -860 580102
rect -804 580046 -736 580102
rect -680 580046 -612 580102
rect -556 580046 -488 580102
rect -432 580046 -336 580102
rect -956 579978 -336 580046
rect -956 579922 -860 579978
rect -804 579922 -736 579978
rect -680 579922 -612 579978
rect -556 579922 -488 579978
rect -432 579922 -336 579978
rect -956 562350 -336 579922
rect -956 562294 -860 562350
rect -804 562294 -736 562350
rect -680 562294 -612 562350
rect -556 562294 -488 562350
rect -432 562294 -336 562350
rect -956 562226 -336 562294
rect -956 562170 -860 562226
rect -804 562170 -736 562226
rect -680 562170 -612 562226
rect -556 562170 -488 562226
rect -432 562170 -336 562226
rect -956 562102 -336 562170
rect -956 562046 -860 562102
rect -804 562046 -736 562102
rect -680 562046 -612 562102
rect -556 562046 -488 562102
rect -432 562046 -336 562102
rect -956 561978 -336 562046
rect -956 561922 -860 561978
rect -804 561922 -736 561978
rect -680 561922 -612 561978
rect -556 561922 -488 561978
rect -432 561922 -336 561978
rect -956 544350 -336 561922
rect -956 544294 -860 544350
rect -804 544294 -736 544350
rect -680 544294 -612 544350
rect -556 544294 -488 544350
rect -432 544294 -336 544350
rect -956 544226 -336 544294
rect -956 544170 -860 544226
rect -804 544170 -736 544226
rect -680 544170 -612 544226
rect -556 544170 -488 544226
rect -432 544170 -336 544226
rect -956 544102 -336 544170
rect -956 544046 -860 544102
rect -804 544046 -736 544102
rect -680 544046 -612 544102
rect -556 544046 -488 544102
rect -432 544046 -336 544102
rect -956 543978 -336 544046
rect -956 543922 -860 543978
rect -804 543922 -736 543978
rect -680 543922 -612 543978
rect -556 543922 -488 543978
rect -432 543922 -336 543978
rect -956 526350 -336 543922
rect -956 526294 -860 526350
rect -804 526294 -736 526350
rect -680 526294 -612 526350
rect -556 526294 -488 526350
rect -432 526294 -336 526350
rect -956 526226 -336 526294
rect -956 526170 -860 526226
rect -804 526170 -736 526226
rect -680 526170 -612 526226
rect -556 526170 -488 526226
rect -432 526170 -336 526226
rect -956 526102 -336 526170
rect -956 526046 -860 526102
rect -804 526046 -736 526102
rect -680 526046 -612 526102
rect -556 526046 -488 526102
rect -432 526046 -336 526102
rect -956 525978 -336 526046
rect -956 525922 -860 525978
rect -804 525922 -736 525978
rect -680 525922 -612 525978
rect -556 525922 -488 525978
rect -432 525922 -336 525978
rect -956 508350 -336 525922
rect -956 508294 -860 508350
rect -804 508294 -736 508350
rect -680 508294 -612 508350
rect -556 508294 -488 508350
rect -432 508294 -336 508350
rect -956 508226 -336 508294
rect -956 508170 -860 508226
rect -804 508170 -736 508226
rect -680 508170 -612 508226
rect -556 508170 -488 508226
rect -432 508170 -336 508226
rect -956 508102 -336 508170
rect -956 508046 -860 508102
rect -804 508046 -736 508102
rect -680 508046 -612 508102
rect -556 508046 -488 508102
rect -432 508046 -336 508102
rect -956 507978 -336 508046
rect -956 507922 -860 507978
rect -804 507922 -736 507978
rect -680 507922 -612 507978
rect -556 507922 -488 507978
rect -432 507922 -336 507978
rect -956 490350 -336 507922
rect -956 490294 -860 490350
rect -804 490294 -736 490350
rect -680 490294 -612 490350
rect -556 490294 -488 490350
rect -432 490294 -336 490350
rect -956 490226 -336 490294
rect -956 490170 -860 490226
rect -804 490170 -736 490226
rect -680 490170 -612 490226
rect -556 490170 -488 490226
rect -432 490170 -336 490226
rect -956 490102 -336 490170
rect -956 490046 -860 490102
rect -804 490046 -736 490102
rect -680 490046 -612 490102
rect -556 490046 -488 490102
rect -432 490046 -336 490102
rect -956 489978 -336 490046
rect -956 489922 -860 489978
rect -804 489922 -736 489978
rect -680 489922 -612 489978
rect -556 489922 -488 489978
rect -432 489922 -336 489978
rect -956 472350 -336 489922
rect -956 472294 -860 472350
rect -804 472294 -736 472350
rect -680 472294 -612 472350
rect -556 472294 -488 472350
rect -432 472294 -336 472350
rect -956 472226 -336 472294
rect -956 472170 -860 472226
rect -804 472170 -736 472226
rect -680 472170 -612 472226
rect -556 472170 -488 472226
rect -432 472170 -336 472226
rect -956 472102 -336 472170
rect -956 472046 -860 472102
rect -804 472046 -736 472102
rect -680 472046 -612 472102
rect -556 472046 -488 472102
rect -432 472046 -336 472102
rect -956 471978 -336 472046
rect -956 471922 -860 471978
rect -804 471922 -736 471978
rect -680 471922 -612 471978
rect -556 471922 -488 471978
rect -432 471922 -336 471978
rect -956 454350 -336 471922
rect -956 454294 -860 454350
rect -804 454294 -736 454350
rect -680 454294 -612 454350
rect -556 454294 -488 454350
rect -432 454294 -336 454350
rect -956 454226 -336 454294
rect -956 454170 -860 454226
rect -804 454170 -736 454226
rect -680 454170 -612 454226
rect -556 454170 -488 454226
rect -432 454170 -336 454226
rect -956 454102 -336 454170
rect -956 454046 -860 454102
rect -804 454046 -736 454102
rect -680 454046 -612 454102
rect -556 454046 -488 454102
rect -432 454046 -336 454102
rect -956 453978 -336 454046
rect -956 453922 -860 453978
rect -804 453922 -736 453978
rect -680 453922 -612 453978
rect -556 453922 -488 453978
rect -432 453922 -336 453978
rect -956 436350 -336 453922
rect -956 436294 -860 436350
rect -804 436294 -736 436350
rect -680 436294 -612 436350
rect -556 436294 -488 436350
rect -432 436294 -336 436350
rect -956 436226 -336 436294
rect -956 436170 -860 436226
rect -804 436170 -736 436226
rect -680 436170 -612 436226
rect -556 436170 -488 436226
rect -432 436170 -336 436226
rect -956 436102 -336 436170
rect -956 436046 -860 436102
rect -804 436046 -736 436102
rect -680 436046 -612 436102
rect -556 436046 -488 436102
rect -432 436046 -336 436102
rect -956 435978 -336 436046
rect -956 435922 -860 435978
rect -804 435922 -736 435978
rect -680 435922 -612 435978
rect -556 435922 -488 435978
rect -432 435922 -336 435978
rect -956 418350 -336 435922
rect -956 418294 -860 418350
rect -804 418294 -736 418350
rect -680 418294 -612 418350
rect -556 418294 -488 418350
rect -432 418294 -336 418350
rect -956 418226 -336 418294
rect -956 418170 -860 418226
rect -804 418170 -736 418226
rect -680 418170 -612 418226
rect -556 418170 -488 418226
rect -432 418170 -336 418226
rect -956 418102 -336 418170
rect -956 418046 -860 418102
rect -804 418046 -736 418102
rect -680 418046 -612 418102
rect -556 418046 -488 418102
rect -432 418046 -336 418102
rect -956 417978 -336 418046
rect -956 417922 -860 417978
rect -804 417922 -736 417978
rect -680 417922 -612 417978
rect -556 417922 -488 417978
rect -432 417922 -336 417978
rect -956 400350 -336 417922
rect -956 400294 -860 400350
rect -804 400294 -736 400350
rect -680 400294 -612 400350
rect -556 400294 -488 400350
rect -432 400294 -336 400350
rect -956 400226 -336 400294
rect -956 400170 -860 400226
rect -804 400170 -736 400226
rect -680 400170 -612 400226
rect -556 400170 -488 400226
rect -432 400170 -336 400226
rect -956 400102 -336 400170
rect -956 400046 -860 400102
rect -804 400046 -736 400102
rect -680 400046 -612 400102
rect -556 400046 -488 400102
rect -432 400046 -336 400102
rect -956 399978 -336 400046
rect -956 399922 -860 399978
rect -804 399922 -736 399978
rect -680 399922 -612 399978
rect -556 399922 -488 399978
rect -432 399922 -336 399978
rect -956 382350 -336 399922
rect -956 382294 -860 382350
rect -804 382294 -736 382350
rect -680 382294 -612 382350
rect -556 382294 -488 382350
rect -432 382294 -336 382350
rect -956 382226 -336 382294
rect -956 382170 -860 382226
rect -804 382170 -736 382226
rect -680 382170 -612 382226
rect -556 382170 -488 382226
rect -432 382170 -336 382226
rect -956 382102 -336 382170
rect -956 382046 -860 382102
rect -804 382046 -736 382102
rect -680 382046 -612 382102
rect -556 382046 -488 382102
rect -432 382046 -336 382102
rect -956 381978 -336 382046
rect -956 381922 -860 381978
rect -804 381922 -736 381978
rect -680 381922 -612 381978
rect -556 381922 -488 381978
rect -432 381922 -336 381978
rect -956 364350 -336 381922
rect -956 364294 -860 364350
rect -804 364294 -736 364350
rect -680 364294 -612 364350
rect -556 364294 -488 364350
rect -432 364294 -336 364350
rect -956 364226 -336 364294
rect -956 364170 -860 364226
rect -804 364170 -736 364226
rect -680 364170 -612 364226
rect -556 364170 -488 364226
rect -432 364170 -336 364226
rect -956 364102 -336 364170
rect -956 364046 -860 364102
rect -804 364046 -736 364102
rect -680 364046 -612 364102
rect -556 364046 -488 364102
rect -432 364046 -336 364102
rect -956 363978 -336 364046
rect -956 363922 -860 363978
rect -804 363922 -736 363978
rect -680 363922 -612 363978
rect -556 363922 -488 363978
rect -432 363922 -336 363978
rect -956 346350 -336 363922
rect -956 346294 -860 346350
rect -804 346294 -736 346350
rect -680 346294 -612 346350
rect -556 346294 -488 346350
rect -432 346294 -336 346350
rect -956 346226 -336 346294
rect -956 346170 -860 346226
rect -804 346170 -736 346226
rect -680 346170 -612 346226
rect -556 346170 -488 346226
rect -432 346170 -336 346226
rect -956 346102 -336 346170
rect -956 346046 -860 346102
rect -804 346046 -736 346102
rect -680 346046 -612 346102
rect -556 346046 -488 346102
rect -432 346046 -336 346102
rect -956 345978 -336 346046
rect -956 345922 -860 345978
rect -804 345922 -736 345978
rect -680 345922 -612 345978
rect -556 345922 -488 345978
rect -432 345922 -336 345978
rect -956 328350 -336 345922
rect -956 328294 -860 328350
rect -804 328294 -736 328350
rect -680 328294 -612 328350
rect -556 328294 -488 328350
rect -432 328294 -336 328350
rect -956 328226 -336 328294
rect -956 328170 -860 328226
rect -804 328170 -736 328226
rect -680 328170 -612 328226
rect -556 328170 -488 328226
rect -432 328170 -336 328226
rect -956 328102 -336 328170
rect -956 328046 -860 328102
rect -804 328046 -736 328102
rect -680 328046 -612 328102
rect -556 328046 -488 328102
rect -432 328046 -336 328102
rect -956 327978 -336 328046
rect -956 327922 -860 327978
rect -804 327922 -736 327978
rect -680 327922 -612 327978
rect -556 327922 -488 327978
rect -432 327922 -336 327978
rect -956 310350 -336 327922
rect -956 310294 -860 310350
rect -804 310294 -736 310350
rect -680 310294 -612 310350
rect -556 310294 -488 310350
rect -432 310294 -336 310350
rect -956 310226 -336 310294
rect -956 310170 -860 310226
rect -804 310170 -736 310226
rect -680 310170 -612 310226
rect -556 310170 -488 310226
rect -432 310170 -336 310226
rect -956 310102 -336 310170
rect -956 310046 -860 310102
rect -804 310046 -736 310102
rect -680 310046 -612 310102
rect -556 310046 -488 310102
rect -432 310046 -336 310102
rect -956 309978 -336 310046
rect -956 309922 -860 309978
rect -804 309922 -736 309978
rect -680 309922 -612 309978
rect -556 309922 -488 309978
rect -432 309922 -336 309978
rect -956 292350 -336 309922
rect -956 292294 -860 292350
rect -804 292294 -736 292350
rect -680 292294 -612 292350
rect -556 292294 -488 292350
rect -432 292294 -336 292350
rect -956 292226 -336 292294
rect -956 292170 -860 292226
rect -804 292170 -736 292226
rect -680 292170 -612 292226
rect -556 292170 -488 292226
rect -432 292170 -336 292226
rect -956 292102 -336 292170
rect -956 292046 -860 292102
rect -804 292046 -736 292102
rect -680 292046 -612 292102
rect -556 292046 -488 292102
rect -432 292046 -336 292102
rect -956 291978 -336 292046
rect -956 291922 -860 291978
rect -804 291922 -736 291978
rect -680 291922 -612 291978
rect -556 291922 -488 291978
rect -432 291922 -336 291978
rect -956 274350 -336 291922
rect -956 274294 -860 274350
rect -804 274294 -736 274350
rect -680 274294 -612 274350
rect -556 274294 -488 274350
rect -432 274294 -336 274350
rect -956 274226 -336 274294
rect -956 274170 -860 274226
rect -804 274170 -736 274226
rect -680 274170 -612 274226
rect -556 274170 -488 274226
rect -432 274170 -336 274226
rect -956 274102 -336 274170
rect -956 274046 -860 274102
rect -804 274046 -736 274102
rect -680 274046 -612 274102
rect -556 274046 -488 274102
rect -432 274046 -336 274102
rect -956 273978 -336 274046
rect -956 273922 -860 273978
rect -804 273922 -736 273978
rect -680 273922 -612 273978
rect -556 273922 -488 273978
rect -432 273922 -336 273978
rect -956 256350 -336 273922
rect -956 256294 -860 256350
rect -804 256294 -736 256350
rect -680 256294 -612 256350
rect -556 256294 -488 256350
rect -432 256294 -336 256350
rect -956 256226 -336 256294
rect -956 256170 -860 256226
rect -804 256170 -736 256226
rect -680 256170 -612 256226
rect -556 256170 -488 256226
rect -432 256170 -336 256226
rect -956 256102 -336 256170
rect -956 256046 -860 256102
rect -804 256046 -736 256102
rect -680 256046 -612 256102
rect -556 256046 -488 256102
rect -432 256046 -336 256102
rect -956 255978 -336 256046
rect -956 255922 -860 255978
rect -804 255922 -736 255978
rect -680 255922 -612 255978
rect -556 255922 -488 255978
rect -432 255922 -336 255978
rect -956 238350 -336 255922
rect -956 238294 -860 238350
rect -804 238294 -736 238350
rect -680 238294 -612 238350
rect -556 238294 -488 238350
rect -432 238294 -336 238350
rect -956 238226 -336 238294
rect -956 238170 -860 238226
rect -804 238170 -736 238226
rect -680 238170 -612 238226
rect -556 238170 -488 238226
rect -432 238170 -336 238226
rect -956 238102 -336 238170
rect -956 238046 -860 238102
rect -804 238046 -736 238102
rect -680 238046 -612 238102
rect -556 238046 -488 238102
rect -432 238046 -336 238102
rect -956 237978 -336 238046
rect -956 237922 -860 237978
rect -804 237922 -736 237978
rect -680 237922 -612 237978
rect -556 237922 -488 237978
rect -432 237922 -336 237978
rect -956 220350 -336 237922
rect -956 220294 -860 220350
rect -804 220294 -736 220350
rect -680 220294 -612 220350
rect -556 220294 -488 220350
rect -432 220294 -336 220350
rect -956 220226 -336 220294
rect -956 220170 -860 220226
rect -804 220170 -736 220226
rect -680 220170 -612 220226
rect -556 220170 -488 220226
rect -432 220170 -336 220226
rect -956 220102 -336 220170
rect -956 220046 -860 220102
rect -804 220046 -736 220102
rect -680 220046 -612 220102
rect -556 220046 -488 220102
rect -432 220046 -336 220102
rect -956 219978 -336 220046
rect -956 219922 -860 219978
rect -804 219922 -736 219978
rect -680 219922 -612 219978
rect -556 219922 -488 219978
rect -432 219922 -336 219978
rect -956 202350 -336 219922
rect -956 202294 -860 202350
rect -804 202294 -736 202350
rect -680 202294 -612 202350
rect -556 202294 -488 202350
rect -432 202294 -336 202350
rect -956 202226 -336 202294
rect -956 202170 -860 202226
rect -804 202170 -736 202226
rect -680 202170 -612 202226
rect -556 202170 -488 202226
rect -432 202170 -336 202226
rect -956 202102 -336 202170
rect -956 202046 -860 202102
rect -804 202046 -736 202102
rect -680 202046 -612 202102
rect -556 202046 -488 202102
rect -432 202046 -336 202102
rect -956 201978 -336 202046
rect -956 201922 -860 201978
rect -804 201922 -736 201978
rect -680 201922 -612 201978
rect -556 201922 -488 201978
rect -432 201922 -336 201978
rect -956 184350 -336 201922
rect -956 184294 -860 184350
rect -804 184294 -736 184350
rect -680 184294 -612 184350
rect -556 184294 -488 184350
rect -432 184294 -336 184350
rect -956 184226 -336 184294
rect -956 184170 -860 184226
rect -804 184170 -736 184226
rect -680 184170 -612 184226
rect -556 184170 -488 184226
rect -432 184170 -336 184226
rect -956 184102 -336 184170
rect -956 184046 -860 184102
rect -804 184046 -736 184102
rect -680 184046 -612 184102
rect -556 184046 -488 184102
rect -432 184046 -336 184102
rect -956 183978 -336 184046
rect -956 183922 -860 183978
rect -804 183922 -736 183978
rect -680 183922 -612 183978
rect -556 183922 -488 183978
rect -432 183922 -336 183978
rect -956 166350 -336 183922
rect -956 166294 -860 166350
rect -804 166294 -736 166350
rect -680 166294 -612 166350
rect -556 166294 -488 166350
rect -432 166294 -336 166350
rect -956 166226 -336 166294
rect -956 166170 -860 166226
rect -804 166170 -736 166226
rect -680 166170 -612 166226
rect -556 166170 -488 166226
rect -432 166170 -336 166226
rect -956 166102 -336 166170
rect -956 166046 -860 166102
rect -804 166046 -736 166102
rect -680 166046 -612 166102
rect -556 166046 -488 166102
rect -432 166046 -336 166102
rect -956 165978 -336 166046
rect -956 165922 -860 165978
rect -804 165922 -736 165978
rect -680 165922 -612 165978
rect -556 165922 -488 165978
rect -432 165922 -336 165978
rect -956 148350 -336 165922
rect -956 148294 -860 148350
rect -804 148294 -736 148350
rect -680 148294 -612 148350
rect -556 148294 -488 148350
rect -432 148294 -336 148350
rect -956 148226 -336 148294
rect -956 148170 -860 148226
rect -804 148170 -736 148226
rect -680 148170 -612 148226
rect -556 148170 -488 148226
rect -432 148170 -336 148226
rect -956 148102 -336 148170
rect -956 148046 -860 148102
rect -804 148046 -736 148102
rect -680 148046 -612 148102
rect -556 148046 -488 148102
rect -432 148046 -336 148102
rect -956 147978 -336 148046
rect -956 147922 -860 147978
rect -804 147922 -736 147978
rect -680 147922 -612 147978
rect -556 147922 -488 147978
rect -432 147922 -336 147978
rect -956 130350 -336 147922
rect -956 130294 -860 130350
rect -804 130294 -736 130350
rect -680 130294 -612 130350
rect -556 130294 -488 130350
rect -432 130294 -336 130350
rect -956 130226 -336 130294
rect -956 130170 -860 130226
rect -804 130170 -736 130226
rect -680 130170 -612 130226
rect -556 130170 -488 130226
rect -432 130170 -336 130226
rect -956 130102 -336 130170
rect -956 130046 -860 130102
rect -804 130046 -736 130102
rect -680 130046 -612 130102
rect -556 130046 -488 130102
rect -432 130046 -336 130102
rect -956 129978 -336 130046
rect -956 129922 -860 129978
rect -804 129922 -736 129978
rect -680 129922 -612 129978
rect -556 129922 -488 129978
rect -432 129922 -336 129978
rect -956 112350 -336 129922
rect -956 112294 -860 112350
rect -804 112294 -736 112350
rect -680 112294 -612 112350
rect -556 112294 -488 112350
rect -432 112294 -336 112350
rect -956 112226 -336 112294
rect -956 112170 -860 112226
rect -804 112170 -736 112226
rect -680 112170 -612 112226
rect -556 112170 -488 112226
rect -432 112170 -336 112226
rect -956 112102 -336 112170
rect -956 112046 -860 112102
rect -804 112046 -736 112102
rect -680 112046 -612 112102
rect -556 112046 -488 112102
rect -432 112046 -336 112102
rect -956 111978 -336 112046
rect -956 111922 -860 111978
rect -804 111922 -736 111978
rect -680 111922 -612 111978
rect -556 111922 -488 111978
rect -432 111922 -336 111978
rect -956 94350 -336 111922
rect -956 94294 -860 94350
rect -804 94294 -736 94350
rect -680 94294 -612 94350
rect -556 94294 -488 94350
rect -432 94294 -336 94350
rect -956 94226 -336 94294
rect -956 94170 -860 94226
rect -804 94170 -736 94226
rect -680 94170 -612 94226
rect -556 94170 -488 94226
rect -432 94170 -336 94226
rect -956 94102 -336 94170
rect -956 94046 -860 94102
rect -804 94046 -736 94102
rect -680 94046 -612 94102
rect -556 94046 -488 94102
rect -432 94046 -336 94102
rect -956 93978 -336 94046
rect -956 93922 -860 93978
rect -804 93922 -736 93978
rect -680 93922 -612 93978
rect -556 93922 -488 93978
rect -432 93922 -336 93978
rect -956 76350 -336 93922
rect -956 76294 -860 76350
rect -804 76294 -736 76350
rect -680 76294 -612 76350
rect -556 76294 -488 76350
rect -432 76294 -336 76350
rect -956 76226 -336 76294
rect -956 76170 -860 76226
rect -804 76170 -736 76226
rect -680 76170 -612 76226
rect -556 76170 -488 76226
rect -432 76170 -336 76226
rect -956 76102 -336 76170
rect -956 76046 -860 76102
rect -804 76046 -736 76102
rect -680 76046 -612 76102
rect -556 76046 -488 76102
rect -432 76046 -336 76102
rect -956 75978 -336 76046
rect -956 75922 -860 75978
rect -804 75922 -736 75978
rect -680 75922 -612 75978
rect -556 75922 -488 75978
rect -432 75922 -336 75978
rect -956 58350 -336 75922
rect -956 58294 -860 58350
rect -804 58294 -736 58350
rect -680 58294 -612 58350
rect -556 58294 -488 58350
rect -432 58294 -336 58350
rect -956 58226 -336 58294
rect -956 58170 -860 58226
rect -804 58170 -736 58226
rect -680 58170 -612 58226
rect -556 58170 -488 58226
rect -432 58170 -336 58226
rect -956 58102 -336 58170
rect -956 58046 -860 58102
rect -804 58046 -736 58102
rect -680 58046 -612 58102
rect -556 58046 -488 58102
rect -432 58046 -336 58102
rect -956 57978 -336 58046
rect -956 57922 -860 57978
rect -804 57922 -736 57978
rect -680 57922 -612 57978
rect -556 57922 -488 57978
rect -432 57922 -336 57978
rect -956 40350 -336 57922
rect -956 40294 -860 40350
rect -804 40294 -736 40350
rect -680 40294 -612 40350
rect -556 40294 -488 40350
rect -432 40294 -336 40350
rect -956 40226 -336 40294
rect -956 40170 -860 40226
rect -804 40170 -736 40226
rect -680 40170 -612 40226
rect -556 40170 -488 40226
rect -432 40170 -336 40226
rect -956 40102 -336 40170
rect -956 40046 -860 40102
rect -804 40046 -736 40102
rect -680 40046 -612 40102
rect -556 40046 -488 40102
rect -432 40046 -336 40102
rect -956 39978 -336 40046
rect -956 39922 -860 39978
rect -804 39922 -736 39978
rect -680 39922 -612 39978
rect -556 39922 -488 39978
rect -432 39922 -336 39978
rect -956 22350 -336 39922
rect -956 22294 -860 22350
rect -804 22294 -736 22350
rect -680 22294 -612 22350
rect -556 22294 -488 22350
rect -432 22294 -336 22350
rect -956 22226 -336 22294
rect -956 22170 -860 22226
rect -804 22170 -736 22226
rect -680 22170 -612 22226
rect -556 22170 -488 22226
rect -432 22170 -336 22226
rect -956 22102 -336 22170
rect -956 22046 -860 22102
rect -804 22046 -736 22102
rect -680 22046 -612 22102
rect -556 22046 -488 22102
rect -432 22046 -336 22102
rect -956 21978 -336 22046
rect -956 21922 -860 21978
rect -804 21922 -736 21978
rect -680 21922 -612 21978
rect -556 21922 -488 21978
rect -432 21922 -336 21978
rect -956 4350 -336 21922
rect -956 4294 -860 4350
rect -804 4294 -736 4350
rect -680 4294 -612 4350
rect -556 4294 -488 4350
rect -432 4294 -336 4350
rect -956 4226 -336 4294
rect -956 4170 -860 4226
rect -804 4170 -736 4226
rect -680 4170 -612 4226
rect -556 4170 -488 4226
rect -432 4170 -336 4226
rect -956 4102 -336 4170
rect -956 4046 -860 4102
rect -804 4046 -736 4102
rect -680 4046 -612 4102
rect -556 4046 -488 4102
rect -432 4046 -336 4102
rect -956 3978 -336 4046
rect -956 3922 -860 3978
rect -804 3922 -736 3978
rect -680 3922 -612 3978
rect -556 3922 -488 3978
rect -432 3922 -336 3978
rect -956 -160 -336 3922
rect -956 -216 -860 -160
rect -804 -216 -736 -160
rect -680 -216 -612 -160
rect -556 -216 -488 -160
rect -432 -216 -336 -160
rect -956 -284 -336 -216
rect -956 -340 -860 -284
rect -804 -340 -736 -284
rect -680 -340 -612 -284
rect -556 -340 -488 -284
rect -432 -340 -336 -284
rect -956 -408 -336 -340
rect -956 -464 -860 -408
rect -804 -464 -736 -408
rect -680 -464 -612 -408
rect -556 -464 -488 -408
rect -432 -464 -336 -408
rect -956 -532 -336 -464
rect -956 -588 -860 -532
rect -804 -588 -736 -532
rect -680 -588 -612 -532
rect -556 -588 -488 -532
rect -432 -588 -336 -532
rect -956 -684 -336 -588
rect 5418 597212 6038 598268
rect 5418 597156 5514 597212
rect 5570 597156 5638 597212
rect 5694 597156 5762 597212
rect 5818 597156 5886 597212
rect 5942 597156 6038 597212
rect 5418 597088 6038 597156
rect 5418 597032 5514 597088
rect 5570 597032 5638 597088
rect 5694 597032 5762 597088
rect 5818 597032 5886 597088
rect 5942 597032 6038 597088
rect 5418 596964 6038 597032
rect 5418 596908 5514 596964
rect 5570 596908 5638 596964
rect 5694 596908 5762 596964
rect 5818 596908 5886 596964
rect 5942 596908 6038 596964
rect 5418 596840 6038 596908
rect 5418 596784 5514 596840
rect 5570 596784 5638 596840
rect 5694 596784 5762 596840
rect 5818 596784 5886 596840
rect 5942 596784 6038 596840
rect 5418 580350 6038 596784
rect 5418 580294 5514 580350
rect 5570 580294 5638 580350
rect 5694 580294 5762 580350
rect 5818 580294 5886 580350
rect 5942 580294 6038 580350
rect 5418 580226 6038 580294
rect 5418 580170 5514 580226
rect 5570 580170 5638 580226
rect 5694 580170 5762 580226
rect 5818 580170 5886 580226
rect 5942 580170 6038 580226
rect 5418 580102 6038 580170
rect 5418 580046 5514 580102
rect 5570 580046 5638 580102
rect 5694 580046 5762 580102
rect 5818 580046 5886 580102
rect 5942 580046 6038 580102
rect 5418 579978 6038 580046
rect 5418 579922 5514 579978
rect 5570 579922 5638 579978
rect 5694 579922 5762 579978
rect 5818 579922 5886 579978
rect 5942 579922 6038 579978
rect 5418 562350 6038 579922
rect 5418 562294 5514 562350
rect 5570 562294 5638 562350
rect 5694 562294 5762 562350
rect 5818 562294 5886 562350
rect 5942 562294 6038 562350
rect 5418 562226 6038 562294
rect 5418 562170 5514 562226
rect 5570 562170 5638 562226
rect 5694 562170 5762 562226
rect 5818 562170 5886 562226
rect 5942 562170 6038 562226
rect 5418 562102 6038 562170
rect 5418 562046 5514 562102
rect 5570 562046 5638 562102
rect 5694 562046 5762 562102
rect 5818 562046 5886 562102
rect 5942 562046 6038 562102
rect 5418 561978 6038 562046
rect 5418 561922 5514 561978
rect 5570 561922 5638 561978
rect 5694 561922 5762 561978
rect 5818 561922 5886 561978
rect 5942 561922 6038 561978
rect 5418 544350 6038 561922
rect 5418 544294 5514 544350
rect 5570 544294 5638 544350
rect 5694 544294 5762 544350
rect 5818 544294 5886 544350
rect 5942 544294 6038 544350
rect 5418 544226 6038 544294
rect 5418 544170 5514 544226
rect 5570 544170 5638 544226
rect 5694 544170 5762 544226
rect 5818 544170 5886 544226
rect 5942 544170 6038 544226
rect 5418 544102 6038 544170
rect 5418 544046 5514 544102
rect 5570 544046 5638 544102
rect 5694 544046 5762 544102
rect 5818 544046 5886 544102
rect 5942 544046 6038 544102
rect 5418 543978 6038 544046
rect 5418 543922 5514 543978
rect 5570 543922 5638 543978
rect 5694 543922 5762 543978
rect 5818 543922 5886 543978
rect 5942 543922 6038 543978
rect 5418 526350 6038 543922
rect 5418 526294 5514 526350
rect 5570 526294 5638 526350
rect 5694 526294 5762 526350
rect 5818 526294 5886 526350
rect 5942 526294 6038 526350
rect 5418 526226 6038 526294
rect 5418 526170 5514 526226
rect 5570 526170 5638 526226
rect 5694 526170 5762 526226
rect 5818 526170 5886 526226
rect 5942 526170 6038 526226
rect 5418 526102 6038 526170
rect 5418 526046 5514 526102
rect 5570 526046 5638 526102
rect 5694 526046 5762 526102
rect 5818 526046 5886 526102
rect 5942 526046 6038 526102
rect 5418 525978 6038 526046
rect 5418 525922 5514 525978
rect 5570 525922 5638 525978
rect 5694 525922 5762 525978
rect 5818 525922 5886 525978
rect 5942 525922 6038 525978
rect 5418 508350 6038 525922
rect 5418 508294 5514 508350
rect 5570 508294 5638 508350
rect 5694 508294 5762 508350
rect 5818 508294 5886 508350
rect 5942 508294 6038 508350
rect 5418 508226 6038 508294
rect 5418 508170 5514 508226
rect 5570 508170 5638 508226
rect 5694 508170 5762 508226
rect 5818 508170 5886 508226
rect 5942 508170 6038 508226
rect 5418 508102 6038 508170
rect 5418 508046 5514 508102
rect 5570 508046 5638 508102
rect 5694 508046 5762 508102
rect 5818 508046 5886 508102
rect 5942 508046 6038 508102
rect 5418 507978 6038 508046
rect 5418 507922 5514 507978
rect 5570 507922 5638 507978
rect 5694 507922 5762 507978
rect 5818 507922 5886 507978
rect 5942 507922 6038 507978
rect 5418 490350 6038 507922
rect 5418 490294 5514 490350
rect 5570 490294 5638 490350
rect 5694 490294 5762 490350
rect 5818 490294 5886 490350
rect 5942 490294 6038 490350
rect 5418 490226 6038 490294
rect 5418 490170 5514 490226
rect 5570 490170 5638 490226
rect 5694 490170 5762 490226
rect 5818 490170 5886 490226
rect 5942 490170 6038 490226
rect 5418 490102 6038 490170
rect 5418 490046 5514 490102
rect 5570 490046 5638 490102
rect 5694 490046 5762 490102
rect 5818 490046 5886 490102
rect 5942 490046 6038 490102
rect 5418 489978 6038 490046
rect 5418 489922 5514 489978
rect 5570 489922 5638 489978
rect 5694 489922 5762 489978
rect 5818 489922 5886 489978
rect 5942 489922 6038 489978
rect 5418 472350 6038 489922
rect 5418 472294 5514 472350
rect 5570 472294 5638 472350
rect 5694 472294 5762 472350
rect 5818 472294 5886 472350
rect 5942 472294 6038 472350
rect 5418 472226 6038 472294
rect 5418 472170 5514 472226
rect 5570 472170 5638 472226
rect 5694 472170 5762 472226
rect 5818 472170 5886 472226
rect 5942 472170 6038 472226
rect 5418 472102 6038 472170
rect 5418 472046 5514 472102
rect 5570 472046 5638 472102
rect 5694 472046 5762 472102
rect 5818 472046 5886 472102
rect 5942 472046 6038 472102
rect 5418 471978 6038 472046
rect 5418 471922 5514 471978
rect 5570 471922 5638 471978
rect 5694 471922 5762 471978
rect 5818 471922 5886 471978
rect 5942 471922 6038 471978
rect 5418 454350 6038 471922
rect 5418 454294 5514 454350
rect 5570 454294 5638 454350
rect 5694 454294 5762 454350
rect 5818 454294 5886 454350
rect 5942 454294 6038 454350
rect 5418 454226 6038 454294
rect 5418 454170 5514 454226
rect 5570 454170 5638 454226
rect 5694 454170 5762 454226
rect 5818 454170 5886 454226
rect 5942 454170 6038 454226
rect 5418 454102 6038 454170
rect 5418 454046 5514 454102
rect 5570 454046 5638 454102
rect 5694 454046 5762 454102
rect 5818 454046 5886 454102
rect 5942 454046 6038 454102
rect 5418 453978 6038 454046
rect 5418 453922 5514 453978
rect 5570 453922 5638 453978
rect 5694 453922 5762 453978
rect 5818 453922 5886 453978
rect 5942 453922 6038 453978
rect 5418 436350 6038 453922
rect 5418 436294 5514 436350
rect 5570 436294 5638 436350
rect 5694 436294 5762 436350
rect 5818 436294 5886 436350
rect 5942 436294 6038 436350
rect 5418 436226 6038 436294
rect 5418 436170 5514 436226
rect 5570 436170 5638 436226
rect 5694 436170 5762 436226
rect 5818 436170 5886 436226
rect 5942 436170 6038 436226
rect 5418 436102 6038 436170
rect 5418 436046 5514 436102
rect 5570 436046 5638 436102
rect 5694 436046 5762 436102
rect 5818 436046 5886 436102
rect 5942 436046 6038 436102
rect 5418 435978 6038 436046
rect 5418 435922 5514 435978
rect 5570 435922 5638 435978
rect 5694 435922 5762 435978
rect 5818 435922 5886 435978
rect 5942 435922 6038 435978
rect 5418 418350 6038 435922
rect 5418 418294 5514 418350
rect 5570 418294 5638 418350
rect 5694 418294 5762 418350
rect 5818 418294 5886 418350
rect 5942 418294 6038 418350
rect 5418 418226 6038 418294
rect 5418 418170 5514 418226
rect 5570 418170 5638 418226
rect 5694 418170 5762 418226
rect 5818 418170 5886 418226
rect 5942 418170 6038 418226
rect 5418 418102 6038 418170
rect 5418 418046 5514 418102
rect 5570 418046 5638 418102
rect 5694 418046 5762 418102
rect 5818 418046 5886 418102
rect 5942 418046 6038 418102
rect 5418 417978 6038 418046
rect 5418 417922 5514 417978
rect 5570 417922 5638 417978
rect 5694 417922 5762 417978
rect 5818 417922 5886 417978
rect 5942 417922 6038 417978
rect 5418 400350 6038 417922
rect 5418 400294 5514 400350
rect 5570 400294 5638 400350
rect 5694 400294 5762 400350
rect 5818 400294 5886 400350
rect 5942 400294 6038 400350
rect 5418 400226 6038 400294
rect 5418 400170 5514 400226
rect 5570 400170 5638 400226
rect 5694 400170 5762 400226
rect 5818 400170 5886 400226
rect 5942 400170 6038 400226
rect 5418 400102 6038 400170
rect 5418 400046 5514 400102
rect 5570 400046 5638 400102
rect 5694 400046 5762 400102
rect 5818 400046 5886 400102
rect 5942 400046 6038 400102
rect 5418 399978 6038 400046
rect 5418 399922 5514 399978
rect 5570 399922 5638 399978
rect 5694 399922 5762 399978
rect 5818 399922 5886 399978
rect 5942 399922 6038 399978
rect 5418 382350 6038 399922
rect 5418 382294 5514 382350
rect 5570 382294 5638 382350
rect 5694 382294 5762 382350
rect 5818 382294 5886 382350
rect 5942 382294 6038 382350
rect 5418 382226 6038 382294
rect 5418 382170 5514 382226
rect 5570 382170 5638 382226
rect 5694 382170 5762 382226
rect 5818 382170 5886 382226
rect 5942 382170 6038 382226
rect 5418 382102 6038 382170
rect 5418 382046 5514 382102
rect 5570 382046 5638 382102
rect 5694 382046 5762 382102
rect 5818 382046 5886 382102
rect 5942 382046 6038 382102
rect 5418 381978 6038 382046
rect 5418 381922 5514 381978
rect 5570 381922 5638 381978
rect 5694 381922 5762 381978
rect 5818 381922 5886 381978
rect 5942 381922 6038 381978
rect 5418 364350 6038 381922
rect 5418 364294 5514 364350
rect 5570 364294 5638 364350
rect 5694 364294 5762 364350
rect 5818 364294 5886 364350
rect 5942 364294 6038 364350
rect 5418 364226 6038 364294
rect 5418 364170 5514 364226
rect 5570 364170 5638 364226
rect 5694 364170 5762 364226
rect 5818 364170 5886 364226
rect 5942 364170 6038 364226
rect 5418 364102 6038 364170
rect 5418 364046 5514 364102
rect 5570 364046 5638 364102
rect 5694 364046 5762 364102
rect 5818 364046 5886 364102
rect 5942 364046 6038 364102
rect 5418 363978 6038 364046
rect 5418 363922 5514 363978
rect 5570 363922 5638 363978
rect 5694 363922 5762 363978
rect 5818 363922 5886 363978
rect 5942 363922 6038 363978
rect 5418 346350 6038 363922
rect 5418 346294 5514 346350
rect 5570 346294 5638 346350
rect 5694 346294 5762 346350
rect 5818 346294 5886 346350
rect 5942 346294 6038 346350
rect 5418 346226 6038 346294
rect 5418 346170 5514 346226
rect 5570 346170 5638 346226
rect 5694 346170 5762 346226
rect 5818 346170 5886 346226
rect 5942 346170 6038 346226
rect 5418 346102 6038 346170
rect 5418 346046 5514 346102
rect 5570 346046 5638 346102
rect 5694 346046 5762 346102
rect 5818 346046 5886 346102
rect 5942 346046 6038 346102
rect 5418 345978 6038 346046
rect 5418 345922 5514 345978
rect 5570 345922 5638 345978
rect 5694 345922 5762 345978
rect 5818 345922 5886 345978
rect 5942 345922 6038 345978
rect 5418 328350 6038 345922
rect 5418 328294 5514 328350
rect 5570 328294 5638 328350
rect 5694 328294 5762 328350
rect 5818 328294 5886 328350
rect 5942 328294 6038 328350
rect 5418 328226 6038 328294
rect 5418 328170 5514 328226
rect 5570 328170 5638 328226
rect 5694 328170 5762 328226
rect 5818 328170 5886 328226
rect 5942 328170 6038 328226
rect 5418 328102 6038 328170
rect 5418 328046 5514 328102
rect 5570 328046 5638 328102
rect 5694 328046 5762 328102
rect 5818 328046 5886 328102
rect 5942 328046 6038 328102
rect 5418 327978 6038 328046
rect 5418 327922 5514 327978
rect 5570 327922 5638 327978
rect 5694 327922 5762 327978
rect 5818 327922 5886 327978
rect 5942 327922 6038 327978
rect 5418 310350 6038 327922
rect 5418 310294 5514 310350
rect 5570 310294 5638 310350
rect 5694 310294 5762 310350
rect 5818 310294 5886 310350
rect 5942 310294 6038 310350
rect 5418 310226 6038 310294
rect 5418 310170 5514 310226
rect 5570 310170 5638 310226
rect 5694 310170 5762 310226
rect 5818 310170 5886 310226
rect 5942 310170 6038 310226
rect 5418 310102 6038 310170
rect 5418 310046 5514 310102
rect 5570 310046 5638 310102
rect 5694 310046 5762 310102
rect 5818 310046 5886 310102
rect 5942 310046 6038 310102
rect 5418 309978 6038 310046
rect 5418 309922 5514 309978
rect 5570 309922 5638 309978
rect 5694 309922 5762 309978
rect 5818 309922 5886 309978
rect 5942 309922 6038 309978
rect 5418 292350 6038 309922
rect 5418 292294 5514 292350
rect 5570 292294 5638 292350
rect 5694 292294 5762 292350
rect 5818 292294 5886 292350
rect 5942 292294 6038 292350
rect 5418 292226 6038 292294
rect 5418 292170 5514 292226
rect 5570 292170 5638 292226
rect 5694 292170 5762 292226
rect 5818 292170 5886 292226
rect 5942 292170 6038 292226
rect 5418 292102 6038 292170
rect 5418 292046 5514 292102
rect 5570 292046 5638 292102
rect 5694 292046 5762 292102
rect 5818 292046 5886 292102
rect 5942 292046 6038 292102
rect 5418 291978 6038 292046
rect 5418 291922 5514 291978
rect 5570 291922 5638 291978
rect 5694 291922 5762 291978
rect 5818 291922 5886 291978
rect 5942 291922 6038 291978
rect 5418 274350 6038 291922
rect 5418 274294 5514 274350
rect 5570 274294 5638 274350
rect 5694 274294 5762 274350
rect 5818 274294 5886 274350
rect 5942 274294 6038 274350
rect 5418 274226 6038 274294
rect 5418 274170 5514 274226
rect 5570 274170 5638 274226
rect 5694 274170 5762 274226
rect 5818 274170 5886 274226
rect 5942 274170 6038 274226
rect 5418 274102 6038 274170
rect 5418 274046 5514 274102
rect 5570 274046 5638 274102
rect 5694 274046 5762 274102
rect 5818 274046 5886 274102
rect 5942 274046 6038 274102
rect 5418 273978 6038 274046
rect 5418 273922 5514 273978
rect 5570 273922 5638 273978
rect 5694 273922 5762 273978
rect 5818 273922 5886 273978
rect 5942 273922 6038 273978
rect 5418 256350 6038 273922
rect 5418 256294 5514 256350
rect 5570 256294 5638 256350
rect 5694 256294 5762 256350
rect 5818 256294 5886 256350
rect 5942 256294 6038 256350
rect 5418 256226 6038 256294
rect 5418 256170 5514 256226
rect 5570 256170 5638 256226
rect 5694 256170 5762 256226
rect 5818 256170 5886 256226
rect 5942 256170 6038 256226
rect 5418 256102 6038 256170
rect 5418 256046 5514 256102
rect 5570 256046 5638 256102
rect 5694 256046 5762 256102
rect 5818 256046 5886 256102
rect 5942 256046 6038 256102
rect 5418 255978 6038 256046
rect 5418 255922 5514 255978
rect 5570 255922 5638 255978
rect 5694 255922 5762 255978
rect 5818 255922 5886 255978
rect 5942 255922 6038 255978
rect 5418 238350 6038 255922
rect 5418 238294 5514 238350
rect 5570 238294 5638 238350
rect 5694 238294 5762 238350
rect 5818 238294 5886 238350
rect 5942 238294 6038 238350
rect 5418 238226 6038 238294
rect 5418 238170 5514 238226
rect 5570 238170 5638 238226
rect 5694 238170 5762 238226
rect 5818 238170 5886 238226
rect 5942 238170 6038 238226
rect 5418 238102 6038 238170
rect 5418 238046 5514 238102
rect 5570 238046 5638 238102
rect 5694 238046 5762 238102
rect 5818 238046 5886 238102
rect 5942 238046 6038 238102
rect 5418 237978 6038 238046
rect 5418 237922 5514 237978
rect 5570 237922 5638 237978
rect 5694 237922 5762 237978
rect 5818 237922 5886 237978
rect 5942 237922 6038 237978
rect 5418 220350 6038 237922
rect 5418 220294 5514 220350
rect 5570 220294 5638 220350
rect 5694 220294 5762 220350
rect 5818 220294 5886 220350
rect 5942 220294 6038 220350
rect 5418 220226 6038 220294
rect 5418 220170 5514 220226
rect 5570 220170 5638 220226
rect 5694 220170 5762 220226
rect 5818 220170 5886 220226
rect 5942 220170 6038 220226
rect 5418 220102 6038 220170
rect 5418 220046 5514 220102
rect 5570 220046 5638 220102
rect 5694 220046 5762 220102
rect 5818 220046 5886 220102
rect 5942 220046 6038 220102
rect 5418 219978 6038 220046
rect 5418 219922 5514 219978
rect 5570 219922 5638 219978
rect 5694 219922 5762 219978
rect 5818 219922 5886 219978
rect 5942 219922 6038 219978
rect 5418 202350 6038 219922
rect 5418 202294 5514 202350
rect 5570 202294 5638 202350
rect 5694 202294 5762 202350
rect 5818 202294 5886 202350
rect 5942 202294 6038 202350
rect 5418 202226 6038 202294
rect 5418 202170 5514 202226
rect 5570 202170 5638 202226
rect 5694 202170 5762 202226
rect 5818 202170 5886 202226
rect 5942 202170 6038 202226
rect 5418 202102 6038 202170
rect 5418 202046 5514 202102
rect 5570 202046 5638 202102
rect 5694 202046 5762 202102
rect 5818 202046 5886 202102
rect 5942 202046 6038 202102
rect 5418 201978 6038 202046
rect 5418 201922 5514 201978
rect 5570 201922 5638 201978
rect 5694 201922 5762 201978
rect 5818 201922 5886 201978
rect 5942 201922 6038 201978
rect 5418 184350 6038 201922
rect 5418 184294 5514 184350
rect 5570 184294 5638 184350
rect 5694 184294 5762 184350
rect 5818 184294 5886 184350
rect 5942 184294 6038 184350
rect 5418 184226 6038 184294
rect 5418 184170 5514 184226
rect 5570 184170 5638 184226
rect 5694 184170 5762 184226
rect 5818 184170 5886 184226
rect 5942 184170 6038 184226
rect 5418 184102 6038 184170
rect 5418 184046 5514 184102
rect 5570 184046 5638 184102
rect 5694 184046 5762 184102
rect 5818 184046 5886 184102
rect 5942 184046 6038 184102
rect 5418 183978 6038 184046
rect 5418 183922 5514 183978
rect 5570 183922 5638 183978
rect 5694 183922 5762 183978
rect 5818 183922 5886 183978
rect 5942 183922 6038 183978
rect 5418 166350 6038 183922
rect 5418 166294 5514 166350
rect 5570 166294 5638 166350
rect 5694 166294 5762 166350
rect 5818 166294 5886 166350
rect 5942 166294 6038 166350
rect 5418 166226 6038 166294
rect 5418 166170 5514 166226
rect 5570 166170 5638 166226
rect 5694 166170 5762 166226
rect 5818 166170 5886 166226
rect 5942 166170 6038 166226
rect 5418 166102 6038 166170
rect 5418 166046 5514 166102
rect 5570 166046 5638 166102
rect 5694 166046 5762 166102
rect 5818 166046 5886 166102
rect 5942 166046 6038 166102
rect 5418 165978 6038 166046
rect 5418 165922 5514 165978
rect 5570 165922 5638 165978
rect 5694 165922 5762 165978
rect 5818 165922 5886 165978
rect 5942 165922 6038 165978
rect 5418 148350 6038 165922
rect 5418 148294 5514 148350
rect 5570 148294 5638 148350
rect 5694 148294 5762 148350
rect 5818 148294 5886 148350
rect 5942 148294 6038 148350
rect 5418 148226 6038 148294
rect 5418 148170 5514 148226
rect 5570 148170 5638 148226
rect 5694 148170 5762 148226
rect 5818 148170 5886 148226
rect 5942 148170 6038 148226
rect 5418 148102 6038 148170
rect 5418 148046 5514 148102
rect 5570 148046 5638 148102
rect 5694 148046 5762 148102
rect 5818 148046 5886 148102
rect 5942 148046 6038 148102
rect 5418 147978 6038 148046
rect 5418 147922 5514 147978
rect 5570 147922 5638 147978
rect 5694 147922 5762 147978
rect 5818 147922 5886 147978
rect 5942 147922 6038 147978
rect 5418 130350 6038 147922
rect 5418 130294 5514 130350
rect 5570 130294 5638 130350
rect 5694 130294 5762 130350
rect 5818 130294 5886 130350
rect 5942 130294 6038 130350
rect 5418 130226 6038 130294
rect 5418 130170 5514 130226
rect 5570 130170 5638 130226
rect 5694 130170 5762 130226
rect 5818 130170 5886 130226
rect 5942 130170 6038 130226
rect 5418 130102 6038 130170
rect 5418 130046 5514 130102
rect 5570 130046 5638 130102
rect 5694 130046 5762 130102
rect 5818 130046 5886 130102
rect 5942 130046 6038 130102
rect 5418 129978 6038 130046
rect 5418 129922 5514 129978
rect 5570 129922 5638 129978
rect 5694 129922 5762 129978
rect 5818 129922 5886 129978
rect 5942 129922 6038 129978
rect 5418 112350 6038 129922
rect 5418 112294 5514 112350
rect 5570 112294 5638 112350
rect 5694 112294 5762 112350
rect 5818 112294 5886 112350
rect 5942 112294 6038 112350
rect 5418 112226 6038 112294
rect 5418 112170 5514 112226
rect 5570 112170 5638 112226
rect 5694 112170 5762 112226
rect 5818 112170 5886 112226
rect 5942 112170 6038 112226
rect 5418 112102 6038 112170
rect 5418 112046 5514 112102
rect 5570 112046 5638 112102
rect 5694 112046 5762 112102
rect 5818 112046 5886 112102
rect 5942 112046 6038 112102
rect 5418 111978 6038 112046
rect 5418 111922 5514 111978
rect 5570 111922 5638 111978
rect 5694 111922 5762 111978
rect 5818 111922 5886 111978
rect 5942 111922 6038 111978
rect 5418 94350 6038 111922
rect 5418 94294 5514 94350
rect 5570 94294 5638 94350
rect 5694 94294 5762 94350
rect 5818 94294 5886 94350
rect 5942 94294 6038 94350
rect 5418 94226 6038 94294
rect 5418 94170 5514 94226
rect 5570 94170 5638 94226
rect 5694 94170 5762 94226
rect 5818 94170 5886 94226
rect 5942 94170 6038 94226
rect 5418 94102 6038 94170
rect 5418 94046 5514 94102
rect 5570 94046 5638 94102
rect 5694 94046 5762 94102
rect 5818 94046 5886 94102
rect 5942 94046 6038 94102
rect 5418 93978 6038 94046
rect 5418 93922 5514 93978
rect 5570 93922 5638 93978
rect 5694 93922 5762 93978
rect 5818 93922 5886 93978
rect 5942 93922 6038 93978
rect 5418 76350 6038 93922
rect 5418 76294 5514 76350
rect 5570 76294 5638 76350
rect 5694 76294 5762 76350
rect 5818 76294 5886 76350
rect 5942 76294 6038 76350
rect 5418 76226 6038 76294
rect 5418 76170 5514 76226
rect 5570 76170 5638 76226
rect 5694 76170 5762 76226
rect 5818 76170 5886 76226
rect 5942 76170 6038 76226
rect 5418 76102 6038 76170
rect 5418 76046 5514 76102
rect 5570 76046 5638 76102
rect 5694 76046 5762 76102
rect 5818 76046 5886 76102
rect 5942 76046 6038 76102
rect 5418 75978 6038 76046
rect 5418 75922 5514 75978
rect 5570 75922 5638 75978
rect 5694 75922 5762 75978
rect 5818 75922 5886 75978
rect 5942 75922 6038 75978
rect 5418 58350 6038 75922
rect 5418 58294 5514 58350
rect 5570 58294 5638 58350
rect 5694 58294 5762 58350
rect 5818 58294 5886 58350
rect 5942 58294 6038 58350
rect 5418 58226 6038 58294
rect 5418 58170 5514 58226
rect 5570 58170 5638 58226
rect 5694 58170 5762 58226
rect 5818 58170 5886 58226
rect 5942 58170 6038 58226
rect 5418 58102 6038 58170
rect 5418 58046 5514 58102
rect 5570 58046 5638 58102
rect 5694 58046 5762 58102
rect 5818 58046 5886 58102
rect 5942 58046 6038 58102
rect 5418 57978 6038 58046
rect 5418 57922 5514 57978
rect 5570 57922 5638 57978
rect 5694 57922 5762 57978
rect 5818 57922 5886 57978
rect 5942 57922 6038 57978
rect 5418 40350 6038 57922
rect 5418 40294 5514 40350
rect 5570 40294 5638 40350
rect 5694 40294 5762 40350
rect 5818 40294 5886 40350
rect 5942 40294 6038 40350
rect 5418 40226 6038 40294
rect 5418 40170 5514 40226
rect 5570 40170 5638 40226
rect 5694 40170 5762 40226
rect 5818 40170 5886 40226
rect 5942 40170 6038 40226
rect 5418 40102 6038 40170
rect 5418 40046 5514 40102
rect 5570 40046 5638 40102
rect 5694 40046 5762 40102
rect 5818 40046 5886 40102
rect 5942 40046 6038 40102
rect 5418 39978 6038 40046
rect 5418 39922 5514 39978
rect 5570 39922 5638 39978
rect 5694 39922 5762 39978
rect 5818 39922 5886 39978
rect 5942 39922 6038 39978
rect 5418 22350 6038 39922
rect 5418 22294 5514 22350
rect 5570 22294 5638 22350
rect 5694 22294 5762 22350
rect 5818 22294 5886 22350
rect 5942 22294 6038 22350
rect 5418 22226 6038 22294
rect 5418 22170 5514 22226
rect 5570 22170 5638 22226
rect 5694 22170 5762 22226
rect 5818 22170 5886 22226
rect 5942 22170 6038 22226
rect 5418 22102 6038 22170
rect 5418 22046 5514 22102
rect 5570 22046 5638 22102
rect 5694 22046 5762 22102
rect 5818 22046 5886 22102
rect 5942 22046 6038 22102
rect 5418 21978 6038 22046
rect 5418 21922 5514 21978
rect 5570 21922 5638 21978
rect 5694 21922 5762 21978
rect 5818 21922 5886 21978
rect 5942 21922 6038 21978
rect 5418 4350 6038 21922
rect 5418 4294 5514 4350
rect 5570 4294 5638 4350
rect 5694 4294 5762 4350
rect 5818 4294 5886 4350
rect 5942 4294 6038 4350
rect 5418 4226 6038 4294
rect 5418 4170 5514 4226
rect 5570 4170 5638 4226
rect 5694 4170 5762 4226
rect 5818 4170 5886 4226
rect 5942 4170 6038 4226
rect 5418 4102 6038 4170
rect 5418 4046 5514 4102
rect 5570 4046 5638 4102
rect 5694 4046 5762 4102
rect 5818 4046 5886 4102
rect 5942 4046 6038 4102
rect 5418 3978 6038 4046
rect 5418 3922 5514 3978
rect 5570 3922 5638 3978
rect 5694 3922 5762 3978
rect 5818 3922 5886 3978
rect 5942 3922 6038 3978
rect 5418 -160 6038 3922
rect 5418 -216 5514 -160
rect 5570 -216 5638 -160
rect 5694 -216 5762 -160
rect 5818 -216 5886 -160
rect 5942 -216 6038 -160
rect 5418 -284 6038 -216
rect 5418 -340 5514 -284
rect 5570 -340 5638 -284
rect 5694 -340 5762 -284
rect 5818 -340 5886 -284
rect 5942 -340 6038 -284
rect 5418 -408 6038 -340
rect 5418 -464 5514 -408
rect 5570 -464 5638 -408
rect 5694 -464 5762 -408
rect 5818 -464 5886 -408
rect 5942 -464 6038 -408
rect 5418 -532 6038 -464
rect 5418 -588 5514 -532
rect 5570 -588 5638 -532
rect 5694 -588 5762 -532
rect 5818 -588 5886 -532
rect 5942 -588 6038 -532
rect -1916 -1176 -1820 -1120
rect -1764 -1176 -1696 -1120
rect -1640 -1176 -1572 -1120
rect -1516 -1176 -1448 -1120
rect -1392 -1176 -1296 -1120
rect -1916 -1244 -1296 -1176
rect -1916 -1300 -1820 -1244
rect -1764 -1300 -1696 -1244
rect -1640 -1300 -1572 -1244
rect -1516 -1300 -1448 -1244
rect -1392 -1300 -1296 -1244
rect -1916 -1368 -1296 -1300
rect -1916 -1424 -1820 -1368
rect -1764 -1424 -1696 -1368
rect -1640 -1424 -1572 -1368
rect -1516 -1424 -1448 -1368
rect -1392 -1424 -1296 -1368
rect -1916 -1492 -1296 -1424
rect -1916 -1548 -1820 -1492
rect -1764 -1548 -1696 -1492
rect -1640 -1548 -1572 -1492
rect -1516 -1548 -1448 -1492
rect -1392 -1548 -1296 -1492
rect -1916 -1644 -1296 -1548
rect 5418 -1644 6038 -588
rect 9138 598172 9758 598268
rect 9138 598116 9234 598172
rect 9290 598116 9358 598172
rect 9414 598116 9482 598172
rect 9538 598116 9606 598172
rect 9662 598116 9758 598172
rect 9138 598048 9758 598116
rect 9138 597992 9234 598048
rect 9290 597992 9358 598048
rect 9414 597992 9482 598048
rect 9538 597992 9606 598048
rect 9662 597992 9758 598048
rect 9138 597924 9758 597992
rect 9138 597868 9234 597924
rect 9290 597868 9358 597924
rect 9414 597868 9482 597924
rect 9538 597868 9606 597924
rect 9662 597868 9758 597924
rect 9138 597800 9758 597868
rect 9138 597744 9234 597800
rect 9290 597744 9358 597800
rect 9414 597744 9482 597800
rect 9538 597744 9606 597800
rect 9662 597744 9758 597800
rect 9138 586350 9758 597744
rect 9138 586294 9234 586350
rect 9290 586294 9358 586350
rect 9414 586294 9482 586350
rect 9538 586294 9606 586350
rect 9662 586294 9758 586350
rect 9138 586226 9758 586294
rect 9138 586170 9234 586226
rect 9290 586170 9358 586226
rect 9414 586170 9482 586226
rect 9538 586170 9606 586226
rect 9662 586170 9758 586226
rect 9138 586102 9758 586170
rect 9138 586046 9234 586102
rect 9290 586046 9358 586102
rect 9414 586046 9482 586102
rect 9538 586046 9606 586102
rect 9662 586046 9758 586102
rect 9138 585978 9758 586046
rect 9138 585922 9234 585978
rect 9290 585922 9358 585978
rect 9414 585922 9482 585978
rect 9538 585922 9606 585978
rect 9662 585922 9758 585978
rect 9138 568350 9758 585922
rect 9138 568294 9234 568350
rect 9290 568294 9358 568350
rect 9414 568294 9482 568350
rect 9538 568294 9606 568350
rect 9662 568294 9758 568350
rect 9138 568226 9758 568294
rect 9138 568170 9234 568226
rect 9290 568170 9358 568226
rect 9414 568170 9482 568226
rect 9538 568170 9606 568226
rect 9662 568170 9758 568226
rect 9138 568102 9758 568170
rect 9138 568046 9234 568102
rect 9290 568046 9358 568102
rect 9414 568046 9482 568102
rect 9538 568046 9606 568102
rect 9662 568046 9758 568102
rect 9138 567978 9758 568046
rect 9138 567922 9234 567978
rect 9290 567922 9358 567978
rect 9414 567922 9482 567978
rect 9538 567922 9606 567978
rect 9662 567922 9758 567978
rect 9138 550350 9758 567922
rect 36138 597212 36758 598268
rect 36138 597156 36234 597212
rect 36290 597156 36358 597212
rect 36414 597156 36482 597212
rect 36538 597156 36606 597212
rect 36662 597156 36758 597212
rect 36138 597088 36758 597156
rect 36138 597032 36234 597088
rect 36290 597032 36358 597088
rect 36414 597032 36482 597088
rect 36538 597032 36606 597088
rect 36662 597032 36758 597088
rect 36138 596964 36758 597032
rect 36138 596908 36234 596964
rect 36290 596908 36358 596964
rect 36414 596908 36482 596964
rect 36538 596908 36606 596964
rect 36662 596908 36758 596964
rect 36138 596840 36758 596908
rect 36138 596784 36234 596840
rect 36290 596784 36358 596840
rect 36414 596784 36482 596840
rect 36538 596784 36606 596840
rect 36662 596784 36758 596840
rect 36138 580350 36758 596784
rect 36138 580294 36234 580350
rect 36290 580294 36358 580350
rect 36414 580294 36482 580350
rect 36538 580294 36606 580350
rect 36662 580294 36758 580350
rect 36138 580226 36758 580294
rect 36138 580170 36234 580226
rect 36290 580170 36358 580226
rect 36414 580170 36482 580226
rect 36538 580170 36606 580226
rect 36662 580170 36758 580226
rect 36138 580102 36758 580170
rect 36138 580046 36234 580102
rect 36290 580046 36358 580102
rect 36414 580046 36482 580102
rect 36538 580046 36606 580102
rect 36662 580046 36758 580102
rect 36138 579978 36758 580046
rect 36138 579922 36234 579978
rect 36290 579922 36358 579978
rect 36414 579922 36482 579978
rect 36538 579922 36606 579978
rect 36662 579922 36758 579978
rect 24448 562350 24768 562384
rect 24448 562294 24518 562350
rect 24574 562294 24642 562350
rect 24698 562294 24768 562350
rect 24448 562226 24768 562294
rect 24448 562170 24518 562226
rect 24574 562170 24642 562226
rect 24698 562170 24768 562226
rect 24448 562102 24768 562170
rect 24448 562046 24518 562102
rect 24574 562046 24642 562102
rect 24698 562046 24768 562102
rect 24448 561978 24768 562046
rect 24448 561922 24518 561978
rect 24574 561922 24642 561978
rect 24698 561922 24768 561978
rect 24448 561888 24768 561922
rect 36138 562350 36758 579922
rect 39858 598172 40478 598268
rect 39858 598116 39954 598172
rect 40010 598116 40078 598172
rect 40134 598116 40202 598172
rect 40258 598116 40326 598172
rect 40382 598116 40478 598172
rect 39858 598048 40478 598116
rect 39858 597992 39954 598048
rect 40010 597992 40078 598048
rect 40134 597992 40202 598048
rect 40258 597992 40326 598048
rect 40382 597992 40478 598048
rect 39858 597924 40478 597992
rect 39858 597868 39954 597924
rect 40010 597868 40078 597924
rect 40134 597868 40202 597924
rect 40258 597868 40326 597924
rect 40382 597868 40478 597924
rect 39858 597800 40478 597868
rect 39858 597744 39954 597800
rect 40010 597744 40078 597800
rect 40134 597744 40202 597800
rect 40258 597744 40326 597800
rect 40382 597744 40478 597800
rect 39858 586350 40478 597744
rect 39858 586294 39954 586350
rect 40010 586294 40078 586350
rect 40134 586294 40202 586350
rect 40258 586294 40326 586350
rect 40382 586294 40478 586350
rect 39858 586226 40478 586294
rect 39858 586170 39954 586226
rect 40010 586170 40078 586226
rect 40134 586170 40202 586226
rect 40258 586170 40326 586226
rect 40382 586170 40478 586226
rect 39858 586102 40478 586170
rect 39858 586046 39954 586102
rect 40010 586046 40078 586102
rect 40134 586046 40202 586102
rect 40258 586046 40326 586102
rect 40382 586046 40478 586102
rect 39858 585978 40478 586046
rect 39858 585922 39954 585978
rect 40010 585922 40078 585978
rect 40134 585922 40202 585978
rect 40258 585922 40326 585978
rect 40382 585922 40478 585978
rect 39858 568407 40478 585922
rect 39858 568351 39954 568407
rect 40010 568351 40078 568407
rect 40134 568351 40202 568407
rect 40258 568351 40326 568407
rect 40382 568351 40478 568407
rect 39858 568283 40478 568351
rect 39858 568227 39954 568283
rect 40010 568227 40078 568283
rect 40134 568227 40202 568283
rect 40258 568227 40326 568283
rect 40382 568227 40478 568283
rect 39858 568188 40478 568227
rect 66858 597212 67478 598268
rect 66858 597156 66954 597212
rect 67010 597156 67078 597212
rect 67134 597156 67202 597212
rect 67258 597156 67326 597212
rect 67382 597156 67478 597212
rect 66858 597088 67478 597156
rect 66858 597032 66954 597088
rect 67010 597032 67078 597088
rect 67134 597032 67202 597088
rect 67258 597032 67326 597088
rect 67382 597032 67478 597088
rect 66858 596964 67478 597032
rect 66858 596908 66954 596964
rect 67010 596908 67078 596964
rect 67134 596908 67202 596964
rect 67258 596908 67326 596964
rect 67382 596908 67478 596964
rect 66858 596840 67478 596908
rect 66858 596784 66954 596840
rect 67010 596784 67078 596840
rect 67134 596784 67202 596840
rect 67258 596784 67326 596840
rect 67382 596784 67478 596840
rect 66858 580350 67478 596784
rect 66858 580294 66954 580350
rect 67010 580294 67078 580350
rect 67134 580294 67202 580350
rect 67258 580294 67326 580350
rect 67382 580294 67478 580350
rect 66858 580226 67478 580294
rect 66858 580170 66954 580226
rect 67010 580170 67078 580226
rect 67134 580170 67202 580226
rect 67258 580170 67326 580226
rect 67382 580170 67478 580226
rect 66858 580102 67478 580170
rect 66858 580046 66954 580102
rect 67010 580046 67078 580102
rect 67134 580046 67202 580102
rect 67258 580046 67326 580102
rect 67382 580046 67478 580102
rect 66858 579978 67478 580046
rect 66858 579922 66954 579978
rect 67010 579922 67078 579978
rect 67134 579922 67202 579978
rect 67258 579922 67326 579978
rect 67382 579922 67478 579978
rect 36138 562294 36234 562350
rect 36290 562294 36358 562350
rect 36414 562294 36482 562350
rect 36538 562294 36606 562350
rect 36662 562294 36758 562350
rect 36138 562226 36758 562294
rect 36138 562170 36234 562226
rect 36290 562170 36358 562226
rect 36414 562170 36482 562226
rect 36538 562170 36606 562226
rect 36662 562170 36758 562226
rect 36138 562102 36758 562170
rect 36138 562046 36234 562102
rect 36290 562046 36358 562102
rect 36414 562046 36482 562102
rect 36538 562046 36606 562102
rect 36662 562046 36758 562102
rect 36138 561978 36758 562046
rect 36138 561922 36234 561978
rect 36290 561922 36358 561978
rect 36414 561922 36482 561978
rect 36538 561922 36606 561978
rect 36662 561922 36758 561978
rect 18396 555940 18452 555950
rect 18396 554518 18452 555884
rect 18396 554418 18452 554428
rect 9138 550294 9234 550350
rect 9290 550294 9358 550350
rect 9414 550294 9482 550350
rect 9538 550294 9606 550350
rect 9662 550294 9758 550350
rect 9138 550226 9758 550294
rect 9138 550170 9234 550226
rect 9290 550170 9358 550226
rect 9414 550170 9482 550226
rect 9538 550170 9606 550226
rect 9662 550170 9758 550226
rect 9138 550102 9758 550170
rect 9138 550046 9234 550102
rect 9290 550046 9358 550102
rect 9414 550046 9482 550102
rect 9538 550046 9606 550102
rect 9662 550046 9758 550102
rect 9138 549978 9758 550046
rect 9138 549922 9234 549978
rect 9290 549922 9358 549978
rect 9414 549922 9482 549978
rect 9538 549922 9606 549978
rect 9662 549922 9758 549978
rect 9138 532350 9758 549922
rect 18284 553252 18340 553262
rect 18172 545188 18228 545198
rect 9138 532294 9234 532350
rect 9290 532294 9358 532350
rect 9414 532294 9482 532350
rect 9538 532294 9606 532350
rect 9662 532294 9758 532350
rect 9138 532226 9758 532294
rect 9138 532170 9234 532226
rect 9290 532170 9358 532226
rect 9414 532170 9482 532226
rect 9538 532170 9606 532226
rect 9662 532170 9758 532226
rect 9138 532102 9758 532170
rect 9138 532046 9234 532102
rect 9290 532046 9358 532102
rect 9414 532046 9482 532102
rect 9538 532046 9606 532102
rect 9662 532046 9758 532102
rect 9138 531978 9758 532046
rect 9138 531922 9234 531978
rect 9290 531922 9358 531978
rect 9414 531922 9482 531978
rect 9538 531922 9606 531978
rect 9662 531922 9758 531978
rect 9138 514350 9758 531922
rect 18060 543844 18116 543854
rect 18060 528276 18116 543788
rect 18172 530068 18228 545132
rect 18172 530002 18228 530012
rect 18060 528210 18116 528220
rect 18284 521668 18340 553196
rect 18284 521602 18340 521612
rect 18396 551908 18452 551918
rect 9138 514294 9234 514350
rect 9290 514294 9358 514350
rect 9414 514294 9482 514350
rect 9538 514294 9606 514350
rect 9662 514294 9758 514350
rect 9138 514226 9758 514294
rect 9138 514170 9234 514226
rect 9290 514170 9358 514226
rect 9414 514170 9482 514226
rect 9538 514170 9606 514226
rect 9662 514170 9758 514226
rect 9138 514102 9758 514170
rect 9138 514046 9234 514102
rect 9290 514046 9358 514102
rect 9414 514046 9482 514102
rect 9538 514046 9606 514102
rect 9662 514046 9758 514102
rect 9138 513978 9758 514046
rect 9138 513922 9234 513978
rect 9290 513922 9358 513978
rect 9414 513922 9482 513978
rect 9538 513922 9606 513978
rect 9662 513922 9758 513978
rect 9138 496350 9758 513922
rect 18396 504196 18452 551852
rect 18396 504130 18452 504140
rect 20076 545860 20132 545870
rect 20076 501956 20132 545804
rect 24448 544350 24768 544384
rect 24448 544294 24518 544350
rect 24574 544294 24642 544350
rect 24698 544294 24768 544350
rect 24448 544226 24768 544294
rect 24448 544170 24518 544226
rect 24574 544170 24642 544226
rect 24698 544170 24768 544226
rect 24448 544102 24768 544170
rect 24448 544046 24518 544102
rect 24574 544046 24642 544102
rect 24698 544046 24768 544102
rect 24448 543978 24768 544046
rect 24448 543922 24518 543978
rect 24574 543922 24642 543978
rect 24698 543922 24768 543978
rect 24448 543888 24768 543922
rect 36138 544350 36758 561922
rect 55168 562350 55488 562384
rect 55168 562294 55238 562350
rect 55294 562294 55362 562350
rect 55418 562294 55488 562350
rect 55168 562226 55488 562294
rect 55168 562170 55238 562226
rect 55294 562170 55362 562226
rect 55418 562170 55488 562226
rect 55168 562102 55488 562170
rect 55168 562046 55238 562102
rect 55294 562046 55362 562102
rect 55418 562046 55488 562102
rect 55168 561978 55488 562046
rect 55168 561922 55238 561978
rect 55294 561922 55362 561978
rect 55418 561922 55488 561978
rect 55168 561888 55488 561922
rect 66858 562350 67478 579922
rect 66858 562294 66954 562350
rect 67010 562294 67078 562350
rect 67134 562294 67202 562350
rect 67258 562294 67326 562350
rect 67382 562294 67478 562350
rect 66858 562226 67478 562294
rect 66858 562170 66954 562226
rect 67010 562170 67078 562226
rect 67134 562170 67202 562226
rect 67258 562170 67326 562226
rect 67382 562170 67478 562226
rect 66858 562102 67478 562170
rect 66858 562046 66954 562102
rect 67010 562046 67078 562102
rect 67134 562046 67202 562102
rect 67258 562046 67326 562102
rect 67382 562046 67478 562102
rect 66858 561978 67478 562046
rect 66858 561922 66954 561978
rect 67010 561922 67078 561978
rect 67134 561922 67202 561978
rect 67258 561922 67326 561978
rect 67382 561922 67478 561978
rect 65100 552580 65156 552590
rect 39808 550350 40128 550384
rect 39808 550294 39878 550350
rect 39934 550294 40002 550350
rect 40058 550294 40128 550350
rect 39808 550226 40128 550294
rect 39808 550170 39878 550226
rect 39934 550170 40002 550226
rect 40058 550170 40128 550226
rect 39808 550102 40128 550170
rect 39808 550046 39878 550102
rect 39934 550046 40002 550102
rect 40058 550046 40128 550102
rect 39808 549978 40128 550046
rect 39808 549922 39878 549978
rect 39934 549922 40002 549978
rect 40058 549922 40128 549978
rect 39808 549888 40128 549922
rect 64652 548548 64708 548558
rect 36138 544294 36234 544350
rect 36290 544294 36358 544350
rect 36414 544294 36482 544350
rect 36538 544294 36606 544350
rect 36662 544294 36758 544350
rect 36138 544226 36758 544294
rect 36138 544170 36234 544226
rect 36290 544170 36358 544226
rect 36414 544170 36482 544226
rect 36538 544170 36606 544226
rect 36662 544170 36758 544226
rect 36138 544102 36758 544170
rect 36138 544046 36234 544102
rect 36290 544046 36358 544102
rect 36414 544046 36482 544102
rect 36538 544046 36606 544102
rect 36662 544046 36758 544102
rect 36138 543978 36758 544046
rect 36138 543922 36234 543978
rect 36290 543922 36358 543978
rect 36414 543922 36482 543978
rect 36538 543922 36606 543978
rect 36662 543922 36758 543978
rect 20076 501890 20132 501900
rect 36138 526350 36758 543922
rect 55168 544350 55488 544384
rect 55168 544294 55238 544350
rect 55294 544294 55362 544350
rect 55418 544294 55488 544350
rect 55168 544226 55488 544294
rect 55168 544170 55238 544226
rect 55294 544170 55362 544226
rect 55418 544170 55488 544226
rect 55168 544102 55488 544170
rect 55168 544046 55238 544102
rect 55294 544046 55362 544102
rect 55418 544046 55488 544102
rect 55168 543978 55488 544046
rect 55168 543922 55238 543978
rect 55294 543922 55362 543978
rect 55418 543922 55488 543978
rect 55168 543888 55488 543922
rect 39808 532350 40128 532384
rect 39808 532294 39878 532350
rect 39934 532294 40002 532350
rect 40058 532294 40128 532350
rect 39808 532226 40128 532294
rect 39808 532170 39878 532226
rect 39934 532170 40002 532226
rect 40058 532170 40128 532226
rect 39808 532102 40128 532170
rect 39808 532046 39878 532102
rect 39934 532046 40002 532102
rect 40058 532046 40128 532102
rect 39808 531978 40128 532046
rect 39808 531922 39878 531978
rect 39934 531922 40002 531978
rect 40058 531922 40128 531978
rect 39808 531888 40128 531922
rect 36138 526294 36234 526350
rect 36290 526294 36358 526350
rect 36414 526294 36482 526350
rect 36538 526294 36606 526350
rect 36662 526294 36758 526350
rect 36138 526226 36758 526294
rect 36138 526170 36234 526226
rect 36290 526170 36358 526226
rect 36414 526170 36482 526226
rect 36538 526170 36606 526226
rect 36662 526170 36758 526226
rect 36138 526102 36758 526170
rect 36138 526046 36234 526102
rect 36290 526046 36358 526102
rect 36414 526046 36482 526102
rect 36538 526046 36606 526102
rect 36662 526046 36758 526102
rect 36138 525978 36758 526046
rect 36138 525922 36234 525978
rect 36290 525922 36358 525978
rect 36414 525922 36482 525978
rect 36538 525922 36606 525978
rect 36662 525922 36758 525978
rect 36138 508350 36758 525922
rect 36138 508294 36234 508350
rect 36290 508294 36358 508350
rect 36414 508294 36482 508350
rect 36538 508294 36606 508350
rect 36662 508294 36758 508350
rect 36138 508226 36758 508294
rect 36138 508170 36234 508226
rect 36290 508170 36358 508226
rect 36414 508170 36482 508226
rect 36538 508170 36606 508226
rect 36662 508170 36758 508226
rect 36138 508102 36758 508170
rect 36138 508046 36234 508102
rect 36290 508046 36358 508102
rect 36414 508046 36482 508102
rect 36538 508046 36606 508102
rect 36662 508046 36758 508102
rect 36138 507978 36758 508046
rect 36138 507922 36234 507978
rect 36290 507922 36358 507978
rect 36414 507922 36482 507978
rect 36538 507922 36606 507978
rect 36662 507922 36758 507978
rect 9138 496294 9234 496350
rect 9290 496294 9358 496350
rect 9414 496294 9482 496350
rect 9538 496294 9606 496350
rect 9662 496294 9758 496350
rect 9138 496226 9758 496294
rect 9138 496170 9234 496226
rect 9290 496170 9358 496226
rect 9414 496170 9482 496226
rect 9538 496170 9606 496226
rect 9662 496170 9758 496226
rect 9138 496102 9758 496170
rect 9138 496046 9234 496102
rect 9290 496046 9358 496102
rect 9414 496046 9482 496102
rect 9538 496046 9606 496102
rect 9662 496046 9758 496102
rect 9138 495978 9758 496046
rect 9138 495922 9234 495978
rect 9290 495922 9358 495978
rect 9414 495922 9482 495978
rect 9538 495922 9606 495978
rect 9662 495922 9758 495978
rect 9138 478350 9758 495922
rect 24448 490350 24768 490384
rect 24448 490294 24518 490350
rect 24574 490294 24642 490350
rect 24698 490294 24768 490350
rect 24448 490226 24768 490294
rect 24448 490170 24518 490226
rect 24574 490170 24642 490226
rect 24698 490170 24768 490226
rect 24448 490102 24768 490170
rect 24448 490046 24518 490102
rect 24574 490046 24642 490102
rect 24698 490046 24768 490102
rect 24448 489978 24768 490046
rect 24448 489922 24518 489978
rect 24574 489922 24642 489978
rect 24698 489922 24768 489978
rect 24448 489888 24768 489922
rect 36138 490350 36758 507922
rect 64652 506436 64708 548492
rect 64652 506370 64708 506380
rect 64764 545860 64820 545870
rect 64764 505316 64820 545804
rect 64988 544516 65044 544526
rect 64764 505250 64820 505260
rect 64876 538468 64932 538478
rect 64876 502516 64932 538412
rect 64988 504756 65044 544460
rect 65100 530180 65156 552524
rect 65100 530114 65156 530124
rect 66858 544350 67478 561922
rect 66858 544294 66954 544350
rect 67010 544294 67078 544350
rect 67134 544294 67202 544350
rect 67258 544294 67326 544350
rect 67382 544294 67478 544350
rect 66858 544226 67478 544294
rect 66858 544170 66954 544226
rect 67010 544170 67078 544226
rect 67134 544170 67202 544226
rect 67258 544170 67326 544226
rect 67382 544170 67478 544226
rect 66858 544102 67478 544170
rect 66858 544046 66954 544102
rect 67010 544046 67078 544102
rect 67134 544046 67202 544102
rect 67258 544046 67326 544102
rect 67382 544046 67478 544102
rect 66858 543978 67478 544046
rect 66858 543922 66954 543978
rect 67010 543922 67078 543978
rect 67134 543922 67202 543978
rect 67258 543922 67326 543978
rect 67382 543922 67478 543978
rect 64988 504690 65044 504700
rect 66858 526350 67478 543922
rect 66858 526294 66954 526350
rect 67010 526294 67078 526350
rect 67134 526294 67202 526350
rect 67258 526294 67326 526350
rect 67382 526294 67478 526350
rect 66858 526226 67478 526294
rect 66858 526170 66954 526226
rect 67010 526170 67078 526226
rect 67134 526170 67202 526226
rect 67258 526170 67326 526226
rect 67382 526170 67478 526226
rect 66858 526102 67478 526170
rect 66858 526046 66954 526102
rect 67010 526046 67078 526102
rect 67134 526046 67202 526102
rect 67258 526046 67326 526102
rect 67382 526046 67478 526102
rect 66858 525978 67478 526046
rect 66858 525922 66954 525978
rect 67010 525922 67078 525978
rect 67134 525922 67202 525978
rect 67258 525922 67326 525978
rect 67382 525922 67478 525978
rect 66858 508350 67478 525922
rect 66858 508294 66954 508350
rect 67010 508294 67078 508350
rect 67134 508294 67202 508350
rect 67258 508294 67326 508350
rect 67382 508294 67478 508350
rect 66858 508226 67478 508294
rect 66858 508170 66954 508226
rect 67010 508170 67078 508226
rect 67134 508170 67202 508226
rect 67258 508170 67326 508226
rect 67382 508170 67478 508226
rect 66858 508102 67478 508170
rect 66858 508046 66954 508102
rect 67010 508046 67078 508102
rect 67134 508046 67202 508102
rect 67258 508046 67326 508102
rect 67382 508046 67478 508102
rect 66858 507978 67478 508046
rect 66858 507922 66954 507978
rect 67010 507922 67078 507978
rect 67134 507922 67202 507978
rect 67258 507922 67326 507978
rect 67382 507922 67478 507978
rect 64876 502450 64932 502460
rect 36138 490294 36234 490350
rect 36290 490294 36358 490350
rect 36414 490294 36482 490350
rect 36538 490294 36606 490350
rect 36662 490294 36758 490350
rect 36138 490226 36758 490294
rect 36138 490170 36234 490226
rect 36290 490170 36358 490226
rect 36414 490170 36482 490226
rect 36538 490170 36606 490226
rect 36662 490170 36758 490226
rect 36138 490102 36758 490170
rect 36138 490046 36234 490102
rect 36290 490046 36358 490102
rect 36414 490046 36482 490102
rect 36538 490046 36606 490102
rect 36662 490046 36758 490102
rect 36138 489978 36758 490046
rect 36138 489922 36234 489978
rect 36290 489922 36358 489978
rect 36414 489922 36482 489978
rect 36538 489922 36606 489978
rect 36662 489922 36758 489978
rect 18396 484036 18452 484046
rect 9138 478294 9234 478350
rect 9290 478294 9358 478350
rect 9414 478294 9482 478350
rect 9538 478294 9606 478350
rect 9662 478294 9758 478350
rect 9138 478226 9758 478294
rect 9138 478170 9234 478226
rect 9290 478170 9358 478226
rect 9414 478170 9482 478226
rect 9538 478170 9606 478226
rect 9662 478170 9758 478226
rect 9138 478102 9758 478170
rect 9138 478046 9234 478102
rect 9290 478046 9358 478102
rect 9414 478046 9482 478102
rect 9538 478046 9606 478102
rect 9662 478046 9758 478102
rect 9138 477978 9758 478046
rect 9138 477922 9234 477978
rect 9290 477922 9358 477978
rect 9414 477922 9482 477978
rect 9538 477922 9606 477978
rect 9662 477922 9758 477978
rect 9138 460350 9758 477922
rect 18172 480676 18228 480686
rect 9138 460294 9234 460350
rect 9290 460294 9358 460350
rect 9414 460294 9482 460350
rect 9538 460294 9606 460350
rect 9662 460294 9758 460350
rect 9138 460226 9758 460294
rect 9138 460170 9234 460226
rect 9290 460170 9358 460226
rect 9414 460170 9482 460226
rect 9538 460170 9606 460226
rect 9662 460170 9758 460226
rect 9138 460102 9758 460170
rect 9138 460046 9234 460102
rect 9290 460046 9358 460102
rect 9414 460046 9482 460102
rect 9538 460046 9606 460102
rect 9662 460046 9758 460102
rect 9138 459978 9758 460046
rect 9138 459922 9234 459978
rect 9290 459922 9358 459978
rect 9414 459922 9482 459978
rect 9538 459922 9606 459978
rect 9662 459922 9758 459978
rect 9138 442350 9758 459922
rect 17948 477316 18004 477326
rect 17948 449428 18004 477260
rect 17948 449362 18004 449372
rect 18060 475972 18116 475982
rect 18060 444836 18116 475916
rect 18172 448196 18228 480620
rect 18172 448130 18228 448140
rect 18284 480004 18340 480014
rect 18060 444770 18116 444780
rect 9138 442294 9234 442350
rect 9290 442294 9358 442350
rect 9414 442294 9482 442350
rect 9538 442294 9606 442350
rect 9662 442294 9758 442350
rect 9138 442226 9758 442294
rect 9138 442170 9234 442226
rect 9290 442170 9358 442226
rect 9414 442170 9482 442226
rect 9538 442170 9606 442226
rect 9662 442170 9758 442226
rect 9138 442102 9758 442170
rect 9138 442046 9234 442102
rect 9290 442046 9358 442102
rect 9414 442046 9482 442102
rect 9538 442046 9606 442102
rect 9662 442046 9758 442102
rect 9138 441978 9758 442046
rect 9138 441922 9234 441978
rect 9290 441922 9358 441978
rect 9414 441922 9482 441978
rect 9538 441922 9606 441978
rect 9662 441922 9758 441978
rect 9138 424350 9758 441922
rect 18284 437668 18340 479948
rect 18284 437602 18340 437612
rect 9138 424294 9234 424350
rect 9290 424294 9358 424350
rect 9414 424294 9482 424350
rect 9538 424294 9606 424350
rect 9662 424294 9758 424350
rect 9138 424226 9758 424294
rect 9138 424170 9234 424226
rect 9290 424170 9358 424226
rect 9414 424170 9482 424226
rect 9538 424170 9606 424226
rect 9662 424170 9758 424226
rect 9138 424102 9758 424170
rect 9138 424046 9234 424102
rect 9290 424046 9358 424102
rect 9414 424046 9482 424102
rect 9538 424046 9606 424102
rect 9662 424046 9758 424102
rect 9138 423978 9758 424046
rect 9138 423922 9234 423978
rect 9290 423922 9358 423978
rect 9414 423922 9482 423978
rect 9538 423922 9606 423978
rect 9662 423922 9758 423978
rect 9138 406350 9758 423922
rect 18396 413218 18452 483980
rect 20076 484036 20132 484046
rect 20076 482878 20132 483980
rect 20076 482812 20132 482822
rect 20076 475300 20132 475310
rect 20076 451108 20132 475244
rect 24448 472350 24768 472384
rect 24448 472294 24518 472350
rect 24574 472294 24642 472350
rect 24698 472294 24768 472350
rect 24448 472226 24768 472294
rect 24448 472170 24518 472226
rect 24574 472170 24642 472226
rect 24698 472170 24768 472226
rect 24448 472102 24768 472170
rect 24448 472046 24518 472102
rect 24574 472046 24642 472102
rect 24698 472046 24768 472102
rect 24448 471978 24768 472046
rect 24448 471922 24518 471978
rect 24574 471922 24642 471978
rect 24698 471922 24768 471978
rect 24448 471888 24768 471922
rect 36138 472350 36758 489922
rect 55168 490350 55488 490384
rect 55168 490294 55238 490350
rect 55294 490294 55362 490350
rect 55418 490294 55488 490350
rect 55168 490226 55488 490294
rect 55168 490170 55238 490226
rect 55294 490170 55362 490226
rect 55418 490170 55488 490226
rect 55168 490102 55488 490170
rect 55168 490046 55238 490102
rect 55294 490046 55362 490102
rect 55418 490046 55488 490102
rect 55168 489978 55488 490046
rect 55168 489922 55238 489978
rect 55294 489922 55362 489978
rect 55418 489922 55488 489978
rect 55168 489888 55488 489922
rect 66858 490350 67478 507922
rect 70578 598172 71198 598268
rect 70578 598116 70674 598172
rect 70730 598116 70798 598172
rect 70854 598116 70922 598172
rect 70978 598116 71046 598172
rect 71102 598116 71198 598172
rect 70578 598048 71198 598116
rect 70578 597992 70674 598048
rect 70730 597992 70798 598048
rect 70854 597992 70922 598048
rect 70978 597992 71046 598048
rect 71102 597992 71198 598048
rect 70578 597924 71198 597992
rect 70578 597868 70674 597924
rect 70730 597868 70798 597924
rect 70854 597868 70922 597924
rect 70978 597868 71046 597924
rect 71102 597868 71198 597924
rect 70578 597800 71198 597868
rect 70578 597744 70674 597800
rect 70730 597744 70798 597800
rect 70854 597744 70922 597800
rect 70978 597744 71046 597800
rect 71102 597744 71198 597800
rect 70578 586350 71198 597744
rect 70578 586294 70674 586350
rect 70730 586294 70798 586350
rect 70854 586294 70922 586350
rect 70978 586294 71046 586350
rect 71102 586294 71198 586350
rect 70578 586226 71198 586294
rect 70578 586170 70674 586226
rect 70730 586170 70798 586226
rect 70854 586170 70922 586226
rect 70978 586170 71046 586226
rect 71102 586170 71198 586226
rect 70578 586102 71198 586170
rect 70578 586046 70674 586102
rect 70730 586046 70798 586102
rect 70854 586046 70922 586102
rect 70978 586046 71046 586102
rect 71102 586046 71198 586102
rect 70578 585978 71198 586046
rect 70578 585922 70674 585978
rect 70730 585922 70798 585978
rect 70854 585922 70922 585978
rect 70978 585922 71046 585978
rect 71102 585922 71198 585978
rect 70578 568350 71198 585922
rect 70578 568294 70674 568350
rect 70730 568294 70798 568350
rect 70854 568294 70922 568350
rect 70978 568294 71046 568350
rect 71102 568294 71198 568350
rect 70578 568226 71198 568294
rect 70578 568170 70674 568226
rect 70730 568170 70798 568226
rect 70854 568170 70922 568226
rect 70978 568170 71046 568226
rect 71102 568170 71198 568226
rect 70578 568102 71198 568170
rect 70578 568046 70674 568102
rect 70730 568046 70798 568102
rect 70854 568046 70922 568102
rect 70978 568046 71046 568102
rect 71102 568046 71198 568102
rect 70578 567978 71198 568046
rect 70578 567922 70674 567978
rect 70730 567922 70798 567978
rect 70854 567922 70922 567978
rect 70978 567922 71046 567978
rect 71102 567922 71198 567978
rect 70578 550350 71198 567922
rect 97578 597212 98198 598268
rect 97578 597156 97674 597212
rect 97730 597156 97798 597212
rect 97854 597156 97922 597212
rect 97978 597156 98046 597212
rect 98102 597156 98198 597212
rect 97578 597088 98198 597156
rect 97578 597032 97674 597088
rect 97730 597032 97798 597088
rect 97854 597032 97922 597088
rect 97978 597032 98046 597088
rect 98102 597032 98198 597088
rect 97578 596964 98198 597032
rect 97578 596908 97674 596964
rect 97730 596908 97798 596964
rect 97854 596908 97922 596964
rect 97978 596908 98046 596964
rect 98102 596908 98198 596964
rect 97578 596840 98198 596908
rect 97578 596784 97674 596840
rect 97730 596784 97798 596840
rect 97854 596784 97922 596840
rect 97978 596784 98046 596840
rect 98102 596784 98198 596840
rect 97578 580350 98198 596784
rect 97578 580294 97674 580350
rect 97730 580294 97798 580350
rect 97854 580294 97922 580350
rect 97978 580294 98046 580350
rect 98102 580294 98198 580350
rect 97578 580226 98198 580294
rect 97578 580170 97674 580226
rect 97730 580170 97798 580226
rect 97854 580170 97922 580226
rect 97978 580170 98046 580226
rect 98102 580170 98198 580226
rect 97578 580102 98198 580170
rect 97578 580046 97674 580102
rect 97730 580046 97798 580102
rect 97854 580046 97922 580102
rect 97978 580046 98046 580102
rect 98102 580046 98198 580102
rect 97578 579978 98198 580046
rect 97578 579922 97674 579978
rect 97730 579922 97798 579978
rect 97854 579922 97922 579978
rect 97978 579922 98046 579978
rect 98102 579922 98198 579978
rect 86448 562350 86768 562384
rect 86448 562294 86518 562350
rect 86574 562294 86642 562350
rect 86698 562294 86768 562350
rect 86448 562226 86768 562294
rect 86448 562170 86518 562226
rect 86574 562170 86642 562226
rect 86698 562170 86768 562226
rect 86448 562102 86768 562170
rect 86448 562046 86518 562102
rect 86574 562046 86642 562102
rect 86698 562046 86768 562102
rect 86448 561978 86768 562046
rect 86448 561922 86518 561978
rect 86574 561922 86642 561978
rect 86698 561922 86768 561978
rect 86448 561888 86768 561922
rect 97578 562350 98198 579922
rect 101298 598172 101918 598268
rect 101298 598116 101394 598172
rect 101450 598116 101518 598172
rect 101574 598116 101642 598172
rect 101698 598116 101766 598172
rect 101822 598116 101918 598172
rect 101298 598048 101918 598116
rect 101298 597992 101394 598048
rect 101450 597992 101518 598048
rect 101574 597992 101642 598048
rect 101698 597992 101766 598048
rect 101822 597992 101918 598048
rect 101298 597924 101918 597992
rect 101298 597868 101394 597924
rect 101450 597868 101518 597924
rect 101574 597868 101642 597924
rect 101698 597868 101766 597924
rect 101822 597868 101918 597924
rect 101298 597800 101918 597868
rect 101298 597744 101394 597800
rect 101450 597744 101518 597800
rect 101574 597744 101642 597800
rect 101698 597744 101766 597800
rect 101822 597744 101918 597800
rect 101298 586350 101918 597744
rect 101298 586294 101394 586350
rect 101450 586294 101518 586350
rect 101574 586294 101642 586350
rect 101698 586294 101766 586350
rect 101822 586294 101918 586350
rect 101298 586226 101918 586294
rect 101298 586170 101394 586226
rect 101450 586170 101518 586226
rect 101574 586170 101642 586226
rect 101698 586170 101766 586226
rect 101822 586170 101918 586226
rect 101298 586102 101918 586170
rect 101298 586046 101394 586102
rect 101450 586046 101518 586102
rect 101574 586046 101642 586102
rect 101698 586046 101766 586102
rect 101822 586046 101918 586102
rect 101298 585978 101918 586046
rect 101298 585922 101394 585978
rect 101450 585922 101518 585978
rect 101574 585922 101642 585978
rect 101698 585922 101766 585978
rect 101822 585922 101918 585978
rect 101298 568407 101918 585922
rect 101298 568351 101394 568407
rect 101450 568351 101518 568407
rect 101574 568351 101642 568407
rect 101698 568351 101766 568407
rect 101822 568351 101918 568407
rect 101298 568283 101918 568351
rect 101298 568227 101394 568283
rect 101450 568227 101518 568283
rect 101574 568227 101642 568283
rect 101698 568227 101766 568283
rect 101822 568227 101918 568283
rect 101298 568188 101918 568227
rect 128298 597212 128918 598268
rect 128298 597156 128394 597212
rect 128450 597156 128518 597212
rect 128574 597156 128642 597212
rect 128698 597156 128766 597212
rect 128822 597156 128918 597212
rect 128298 597088 128918 597156
rect 128298 597032 128394 597088
rect 128450 597032 128518 597088
rect 128574 597032 128642 597088
rect 128698 597032 128766 597088
rect 128822 597032 128918 597088
rect 128298 596964 128918 597032
rect 128298 596908 128394 596964
rect 128450 596908 128518 596964
rect 128574 596908 128642 596964
rect 128698 596908 128766 596964
rect 128822 596908 128918 596964
rect 128298 596840 128918 596908
rect 128298 596784 128394 596840
rect 128450 596784 128518 596840
rect 128574 596784 128642 596840
rect 128698 596784 128766 596840
rect 128822 596784 128918 596840
rect 128298 580350 128918 596784
rect 128298 580294 128394 580350
rect 128450 580294 128518 580350
rect 128574 580294 128642 580350
rect 128698 580294 128766 580350
rect 128822 580294 128918 580350
rect 128298 580226 128918 580294
rect 128298 580170 128394 580226
rect 128450 580170 128518 580226
rect 128574 580170 128642 580226
rect 128698 580170 128766 580226
rect 128822 580170 128918 580226
rect 128298 580102 128918 580170
rect 128298 580046 128394 580102
rect 128450 580046 128518 580102
rect 128574 580046 128642 580102
rect 128698 580046 128766 580102
rect 128822 580046 128918 580102
rect 128298 579978 128918 580046
rect 128298 579922 128394 579978
rect 128450 579922 128518 579978
rect 128574 579922 128642 579978
rect 128698 579922 128766 579978
rect 128822 579922 128918 579978
rect 97578 562294 97674 562350
rect 97730 562294 97798 562350
rect 97854 562294 97922 562350
rect 97978 562294 98046 562350
rect 98102 562294 98198 562350
rect 97578 562226 98198 562294
rect 97578 562170 97674 562226
rect 97730 562170 97798 562226
rect 97854 562170 97922 562226
rect 97978 562170 98046 562226
rect 98102 562170 98198 562226
rect 97578 562102 98198 562170
rect 97578 562046 97674 562102
rect 97730 562046 97798 562102
rect 97854 562046 97922 562102
rect 97978 562046 98046 562102
rect 98102 562046 98198 562102
rect 97578 561978 98198 562046
rect 97578 561922 97674 561978
rect 97730 561922 97798 561978
rect 97854 561922 97922 561978
rect 97978 561922 98046 561978
rect 98102 561922 98198 561978
rect 70578 550294 70674 550350
rect 70730 550294 70798 550350
rect 70854 550294 70922 550350
rect 70978 550294 71046 550350
rect 71102 550294 71198 550350
rect 70578 550226 71198 550294
rect 70578 550170 70674 550226
rect 70730 550170 70798 550226
rect 70854 550170 70922 550226
rect 70978 550170 71046 550226
rect 71102 550170 71198 550226
rect 70578 550102 71198 550170
rect 70578 550046 70674 550102
rect 70730 550046 70798 550102
rect 70854 550046 70922 550102
rect 70978 550046 71046 550102
rect 71102 550046 71198 550102
rect 70578 549978 71198 550046
rect 70578 549922 70674 549978
rect 70730 549922 70798 549978
rect 70854 549922 70922 549978
rect 70978 549922 71046 549978
rect 71102 549922 71198 549978
rect 70578 532350 71198 549922
rect 80108 555268 80164 555278
rect 70578 532294 70674 532350
rect 70730 532294 70798 532350
rect 70854 532294 70922 532350
rect 70978 532294 71046 532350
rect 71102 532294 71198 532350
rect 70578 532226 71198 532294
rect 70578 532170 70674 532226
rect 70730 532170 70798 532226
rect 70854 532170 70922 532226
rect 70978 532170 71046 532226
rect 71102 532170 71198 532226
rect 70578 532102 71198 532170
rect 70578 532046 70674 532102
rect 70730 532046 70798 532102
rect 70854 532046 70922 532102
rect 70978 532046 71046 532102
rect 71102 532046 71198 532102
rect 70578 531978 71198 532046
rect 70578 531922 70674 531978
rect 70730 531922 70798 531978
rect 70854 531922 70922 531978
rect 70978 531922 71046 531978
rect 71102 531922 71198 531978
rect 70578 514350 71198 531922
rect 70578 514294 70674 514350
rect 70730 514294 70798 514350
rect 70854 514294 70922 514350
rect 70978 514294 71046 514350
rect 71102 514294 71198 514350
rect 70578 514226 71198 514294
rect 70578 514170 70674 514226
rect 70730 514170 70798 514226
rect 70854 514170 70922 514226
rect 70978 514170 71046 514226
rect 71102 514170 71198 514226
rect 70578 514102 71198 514170
rect 70578 514046 70674 514102
rect 70730 514046 70798 514102
rect 70854 514046 70922 514102
rect 70978 514046 71046 514102
rect 71102 514046 71198 514102
rect 70578 513978 71198 514046
rect 70578 513922 70674 513978
rect 70730 513922 70798 513978
rect 70854 513922 70922 513978
rect 70978 513922 71046 513978
rect 71102 513922 71198 513978
rect 70578 496350 71198 513922
rect 74732 549892 74788 549902
rect 74732 504868 74788 549836
rect 74844 549220 74900 549230
rect 74844 509908 74900 549164
rect 80108 514948 80164 555212
rect 80444 554596 80500 554606
rect 80332 551236 80388 551246
rect 80220 544516 80276 544526
rect 80220 528052 80276 544460
rect 80220 527986 80276 527996
rect 80332 518308 80388 551180
rect 80444 520100 80500 554540
rect 82684 554518 82740 554528
rect 82684 553924 82740 554462
rect 82684 553858 82740 553868
rect 80444 520034 80500 520044
rect 82012 549220 82068 549230
rect 80332 518242 80388 518252
rect 82012 515956 82068 549164
rect 82236 547204 82292 547214
rect 82124 546532 82180 546542
rect 82124 518420 82180 546476
rect 82236 519988 82292 547148
rect 86448 544350 86768 544384
rect 86448 544294 86518 544350
rect 86574 544294 86642 544350
rect 86698 544294 86768 544350
rect 86448 544226 86768 544294
rect 86448 544170 86518 544226
rect 86574 544170 86642 544226
rect 86698 544170 86768 544226
rect 86448 544102 86768 544170
rect 86448 544046 86518 544102
rect 86574 544046 86642 544102
rect 86698 544046 86768 544102
rect 86448 543978 86768 544046
rect 86448 543922 86518 543978
rect 86574 543922 86642 543978
rect 86698 543922 86768 543978
rect 86448 543888 86768 543922
rect 97578 544350 98198 561922
rect 117168 562350 117488 562384
rect 117168 562294 117238 562350
rect 117294 562294 117362 562350
rect 117418 562294 117488 562350
rect 117168 562226 117488 562294
rect 117168 562170 117238 562226
rect 117294 562170 117362 562226
rect 117418 562170 117488 562226
rect 117168 562102 117488 562170
rect 117168 562046 117238 562102
rect 117294 562046 117362 562102
rect 117418 562046 117488 562102
rect 117168 561978 117488 562046
rect 117168 561922 117238 561978
rect 117294 561922 117362 561978
rect 117418 561922 117488 561978
rect 117168 561888 117488 561922
rect 128298 562350 128918 579922
rect 128298 562294 128394 562350
rect 128450 562294 128518 562350
rect 128574 562294 128642 562350
rect 128698 562294 128766 562350
rect 128822 562294 128918 562350
rect 128298 562226 128918 562294
rect 128298 562170 128394 562226
rect 128450 562170 128518 562226
rect 128574 562170 128642 562226
rect 128698 562170 128766 562226
rect 128822 562170 128918 562226
rect 128298 562102 128918 562170
rect 128298 562046 128394 562102
rect 128450 562046 128518 562102
rect 128574 562046 128642 562102
rect 128698 562046 128766 562102
rect 128822 562046 128918 562102
rect 128298 561978 128918 562046
rect 128298 561922 128394 561978
rect 128450 561922 128518 561978
rect 128574 561922 128642 561978
rect 128698 561922 128766 561978
rect 128822 561922 128918 561978
rect 126924 554596 126980 554606
rect 101808 550350 102128 550384
rect 101808 550294 101878 550350
rect 101934 550294 102002 550350
rect 102058 550294 102128 550350
rect 101808 550226 102128 550294
rect 101808 550170 101878 550226
rect 101934 550170 102002 550226
rect 102058 550170 102128 550226
rect 101808 550102 102128 550170
rect 101808 550046 101878 550102
rect 101934 550046 102002 550102
rect 102058 550046 102128 550102
rect 101808 549978 102128 550046
rect 101808 549922 101878 549978
rect 101934 549922 102002 549978
rect 102058 549922 102128 549978
rect 101808 549888 102128 549922
rect 126812 547876 126868 547886
rect 97578 544294 97674 544350
rect 97730 544294 97798 544350
rect 97854 544294 97922 544350
rect 97978 544294 98046 544350
rect 98102 544294 98198 544350
rect 97578 544226 98198 544294
rect 97578 544170 97674 544226
rect 97730 544170 97798 544226
rect 97854 544170 97922 544226
rect 97978 544170 98046 544226
rect 98102 544170 98198 544226
rect 97578 544102 98198 544170
rect 97578 544046 97674 544102
rect 97730 544046 97798 544102
rect 97854 544046 97922 544102
rect 97978 544046 98046 544102
rect 98102 544046 98198 544102
rect 97578 543978 98198 544046
rect 97578 543922 97674 543978
rect 97730 543922 97798 543978
rect 97854 543922 97922 543978
rect 97978 543922 98046 543978
rect 98102 543922 98198 543978
rect 82236 519922 82292 519932
rect 97578 526350 98198 543922
rect 117168 544350 117488 544384
rect 117168 544294 117238 544350
rect 117294 544294 117362 544350
rect 117418 544294 117488 544350
rect 117168 544226 117488 544294
rect 117168 544170 117238 544226
rect 117294 544170 117362 544226
rect 117418 544170 117488 544226
rect 117168 544102 117488 544170
rect 117168 544046 117238 544102
rect 117294 544046 117362 544102
rect 117418 544046 117488 544102
rect 117168 543978 117488 544046
rect 117168 543922 117238 543978
rect 117294 543922 117362 543978
rect 117418 543922 117488 543978
rect 117168 543888 117488 543922
rect 101808 532350 102128 532384
rect 101808 532294 101878 532350
rect 101934 532294 102002 532350
rect 102058 532294 102128 532350
rect 101808 532226 102128 532294
rect 101808 532170 101878 532226
rect 101934 532170 102002 532226
rect 102058 532170 102128 532226
rect 101808 532102 102128 532170
rect 101808 532046 101878 532102
rect 101934 532046 102002 532102
rect 102058 532046 102128 532102
rect 101808 531978 102128 532046
rect 101808 531922 101878 531978
rect 101934 531922 102002 531978
rect 102058 531922 102128 531978
rect 101808 531888 102128 531922
rect 97578 526294 97674 526350
rect 97730 526294 97798 526350
rect 97854 526294 97922 526350
rect 97978 526294 98046 526350
rect 98102 526294 98198 526350
rect 97578 526226 98198 526294
rect 97578 526170 97674 526226
rect 97730 526170 97798 526226
rect 97854 526170 97922 526226
rect 97978 526170 98046 526226
rect 98102 526170 98198 526226
rect 97578 526102 98198 526170
rect 97578 526046 97674 526102
rect 97730 526046 97798 526102
rect 97854 526046 97922 526102
rect 97978 526046 98046 526102
rect 98102 526046 98198 526102
rect 97578 525978 98198 526046
rect 97578 525922 97674 525978
rect 97730 525922 97798 525978
rect 97854 525922 97922 525978
rect 97978 525922 98046 525978
rect 98102 525922 98198 525978
rect 82124 518354 82180 518364
rect 82012 515890 82068 515900
rect 80108 514882 80164 514892
rect 74844 509842 74900 509852
rect 74732 504802 74788 504812
rect 97578 508350 98198 525922
rect 126812 513156 126868 547820
rect 126924 521780 126980 554540
rect 127260 552580 127316 552590
rect 126924 521714 126980 521724
rect 127036 547204 127092 547214
rect 127036 513716 127092 547148
rect 127036 513650 127092 513660
rect 127148 545860 127204 545870
rect 126812 513090 126868 513100
rect 127148 510916 127204 545804
rect 127260 526708 127316 552524
rect 127260 526642 127316 526652
rect 128298 544350 128918 561922
rect 128298 544294 128394 544350
rect 128450 544294 128518 544350
rect 128574 544294 128642 544350
rect 128698 544294 128766 544350
rect 128822 544294 128918 544350
rect 128298 544226 128918 544294
rect 128298 544170 128394 544226
rect 128450 544170 128518 544226
rect 128574 544170 128642 544226
rect 128698 544170 128766 544226
rect 128822 544170 128918 544226
rect 128298 544102 128918 544170
rect 128298 544046 128394 544102
rect 128450 544046 128518 544102
rect 128574 544046 128642 544102
rect 128698 544046 128766 544102
rect 128822 544046 128918 544102
rect 128298 543978 128918 544046
rect 128298 543922 128394 543978
rect 128450 543922 128518 543978
rect 128574 543922 128642 543978
rect 128698 543922 128766 543978
rect 128822 543922 128918 543978
rect 127148 510850 127204 510860
rect 128298 526350 128918 543922
rect 128298 526294 128394 526350
rect 128450 526294 128518 526350
rect 128574 526294 128642 526350
rect 128698 526294 128766 526350
rect 128822 526294 128918 526350
rect 128298 526226 128918 526294
rect 128298 526170 128394 526226
rect 128450 526170 128518 526226
rect 128574 526170 128642 526226
rect 128698 526170 128766 526226
rect 128822 526170 128918 526226
rect 128298 526102 128918 526170
rect 128298 526046 128394 526102
rect 128450 526046 128518 526102
rect 128574 526046 128642 526102
rect 128698 526046 128766 526102
rect 128822 526046 128918 526102
rect 128298 525978 128918 526046
rect 128298 525922 128394 525978
rect 128450 525922 128518 525978
rect 128574 525922 128642 525978
rect 128698 525922 128766 525978
rect 128822 525922 128918 525978
rect 97578 508294 97674 508350
rect 97730 508294 97798 508350
rect 97854 508294 97922 508350
rect 97978 508294 98046 508350
rect 98102 508294 98198 508350
rect 97578 508226 98198 508294
rect 97578 508170 97674 508226
rect 97730 508170 97798 508226
rect 97854 508170 97922 508226
rect 97978 508170 98046 508226
rect 98102 508170 98198 508226
rect 97578 508102 98198 508170
rect 97578 508046 97674 508102
rect 97730 508046 97798 508102
rect 97854 508046 97922 508102
rect 97978 508046 98046 508102
rect 98102 508046 98198 508102
rect 97578 507978 98198 508046
rect 97578 507922 97674 507978
rect 97730 507922 97798 507978
rect 97854 507922 97922 507978
rect 97978 507922 98046 507978
rect 98102 507922 98198 507978
rect 70578 496294 70674 496350
rect 70730 496294 70798 496350
rect 70854 496294 70922 496350
rect 70978 496294 71046 496350
rect 71102 496294 71198 496350
rect 70578 496226 71198 496294
rect 70578 496170 70674 496226
rect 70730 496170 70798 496226
rect 70854 496170 70922 496226
rect 70978 496170 71046 496226
rect 71102 496170 71198 496226
rect 70578 496102 71198 496170
rect 70578 496046 70674 496102
rect 70730 496046 70798 496102
rect 70854 496046 70922 496102
rect 70978 496046 71046 496102
rect 71102 496046 71198 496102
rect 70578 495978 71198 496046
rect 70578 495922 70674 495978
rect 70730 495922 70798 495978
rect 70854 495922 70922 495978
rect 70978 495922 71046 495978
rect 71102 495922 71198 495978
rect 66858 490294 66954 490350
rect 67010 490294 67078 490350
rect 67134 490294 67202 490350
rect 67258 490294 67326 490350
rect 67382 490294 67478 490350
rect 66858 490226 67478 490294
rect 66858 490170 66954 490226
rect 67010 490170 67078 490226
rect 67134 490170 67202 490226
rect 67258 490170 67326 490226
rect 67382 490170 67478 490226
rect 66858 490102 67478 490170
rect 66858 490046 66954 490102
rect 67010 490046 67078 490102
rect 67134 490046 67202 490102
rect 67258 490046 67326 490102
rect 67382 490046 67478 490102
rect 66858 489978 67478 490046
rect 66858 489922 66954 489978
rect 67010 489922 67078 489978
rect 67134 489922 67202 489978
rect 67258 489922 67326 489978
rect 67382 489922 67478 489978
rect 64764 483364 64820 483374
rect 39808 478350 40128 478384
rect 39808 478294 39878 478350
rect 39934 478294 40002 478350
rect 40058 478294 40128 478350
rect 39808 478226 40128 478294
rect 39808 478170 39878 478226
rect 39934 478170 40002 478226
rect 40058 478170 40128 478226
rect 39808 478102 40128 478170
rect 39808 478046 39878 478102
rect 39934 478046 40002 478102
rect 40058 478046 40128 478102
rect 39808 477978 40128 478046
rect 39808 477922 39878 477978
rect 39934 477922 40002 477978
rect 40058 477922 40128 477978
rect 39808 477888 40128 477922
rect 64652 475972 64708 475982
rect 36138 472294 36234 472350
rect 36290 472294 36358 472350
rect 36414 472294 36482 472350
rect 36538 472294 36606 472350
rect 36662 472294 36758 472350
rect 36138 472226 36758 472294
rect 36138 472170 36234 472226
rect 36290 472170 36358 472226
rect 36414 472170 36482 472226
rect 36538 472170 36606 472226
rect 36662 472170 36758 472226
rect 36138 472102 36758 472170
rect 36138 472046 36234 472102
rect 36290 472046 36358 472102
rect 36414 472046 36482 472102
rect 36538 472046 36606 472102
rect 36662 472046 36758 472102
rect 36138 471978 36758 472046
rect 36138 471922 36234 471978
rect 36290 471922 36358 471978
rect 36414 471922 36482 471978
rect 36538 471922 36606 471978
rect 36662 471922 36758 471978
rect 20076 451042 20132 451052
rect 36138 454350 36758 471922
rect 55168 472350 55488 472384
rect 55168 472294 55238 472350
rect 55294 472294 55362 472350
rect 55418 472294 55488 472350
rect 55168 472226 55488 472294
rect 55168 472170 55238 472226
rect 55294 472170 55362 472226
rect 55418 472170 55488 472226
rect 55168 472102 55488 472170
rect 55168 472046 55238 472102
rect 55294 472046 55362 472102
rect 55418 472046 55488 472102
rect 55168 471978 55488 472046
rect 55168 471922 55238 471978
rect 55294 471922 55362 471978
rect 55418 471922 55488 471978
rect 55168 471888 55488 471922
rect 39808 460350 40128 460384
rect 39808 460294 39878 460350
rect 39934 460294 40002 460350
rect 40058 460294 40128 460350
rect 39808 460226 40128 460294
rect 39808 460170 39878 460226
rect 39934 460170 40002 460226
rect 40058 460170 40128 460226
rect 39808 460102 40128 460170
rect 39808 460046 39878 460102
rect 39934 460046 40002 460102
rect 40058 460046 40128 460102
rect 39808 459978 40128 460046
rect 39808 459922 39878 459978
rect 39934 459922 40002 459978
rect 40058 459922 40128 459978
rect 39808 459888 40128 459922
rect 36138 454294 36234 454350
rect 36290 454294 36358 454350
rect 36414 454294 36482 454350
rect 36538 454294 36606 454350
rect 36662 454294 36758 454350
rect 36138 454226 36758 454294
rect 36138 454170 36234 454226
rect 36290 454170 36358 454226
rect 36414 454170 36482 454226
rect 36538 454170 36606 454226
rect 36662 454170 36758 454226
rect 36138 454102 36758 454170
rect 36138 454046 36234 454102
rect 36290 454046 36358 454102
rect 36414 454046 36482 454102
rect 36538 454046 36606 454102
rect 36662 454046 36758 454102
rect 36138 453978 36758 454046
rect 36138 453922 36234 453978
rect 36290 453922 36358 453978
rect 36414 453922 36482 453978
rect 36538 453922 36606 453978
rect 36662 453922 36758 453978
rect 36138 436350 36758 453922
rect 64652 441028 64708 475916
rect 64764 449316 64820 483308
rect 64764 449250 64820 449260
rect 64876 481348 64932 481358
rect 64876 447636 64932 481292
rect 65100 479332 65156 479342
rect 64876 447570 64932 447580
rect 64988 471268 65044 471278
rect 64988 441140 65044 471212
rect 65100 448756 65156 479276
rect 65100 448690 65156 448700
rect 66858 472350 67478 489922
rect 66858 472294 66954 472350
rect 67010 472294 67078 472350
rect 67134 472294 67202 472350
rect 67258 472294 67326 472350
rect 67382 472294 67478 472350
rect 66858 472226 67478 472294
rect 66858 472170 66954 472226
rect 67010 472170 67078 472226
rect 67134 472170 67202 472226
rect 67258 472170 67326 472226
rect 67382 472170 67478 472226
rect 66858 472102 67478 472170
rect 66858 472046 66954 472102
rect 67010 472046 67078 472102
rect 67134 472046 67202 472102
rect 67258 472046 67326 472102
rect 67382 472046 67478 472102
rect 66858 471978 67478 472046
rect 66858 471922 66954 471978
rect 67010 471922 67078 471978
rect 67134 471922 67202 471978
rect 67258 471922 67326 471978
rect 67382 471922 67478 471978
rect 66858 454350 67478 471922
rect 69692 492772 69748 492782
rect 69692 457828 69748 492716
rect 70578 478350 71198 495922
rect 86448 490350 86768 490384
rect 86448 490294 86518 490350
rect 86574 490294 86642 490350
rect 86698 490294 86768 490350
rect 86448 490226 86768 490294
rect 86448 490170 86518 490226
rect 86574 490170 86642 490226
rect 86698 490170 86768 490226
rect 86448 490102 86768 490170
rect 86448 490046 86518 490102
rect 86574 490046 86642 490102
rect 86698 490046 86768 490102
rect 86448 489978 86768 490046
rect 86448 489922 86518 489978
rect 86574 489922 86642 489978
rect 86698 489922 86768 489978
rect 86448 489888 86768 489922
rect 97578 490350 98198 507922
rect 128298 508350 128918 525922
rect 128298 508294 128394 508350
rect 128450 508294 128518 508350
rect 128574 508294 128642 508350
rect 128698 508294 128766 508350
rect 128822 508294 128918 508350
rect 128298 508226 128918 508294
rect 128298 508170 128394 508226
rect 128450 508170 128518 508226
rect 128574 508170 128642 508226
rect 128698 508170 128766 508226
rect 128822 508170 128918 508226
rect 128298 508102 128918 508170
rect 128298 508046 128394 508102
rect 128450 508046 128518 508102
rect 128574 508046 128642 508102
rect 128698 508046 128766 508102
rect 128822 508046 128918 508102
rect 128298 507978 128918 508046
rect 128298 507922 128394 507978
rect 128450 507922 128518 507978
rect 128574 507922 128642 507978
rect 128698 507922 128766 507978
rect 128822 507922 128918 507978
rect 97578 490294 97674 490350
rect 97730 490294 97798 490350
rect 97854 490294 97922 490350
rect 97978 490294 98046 490350
rect 98102 490294 98198 490350
rect 97578 490226 98198 490294
rect 97578 490170 97674 490226
rect 97730 490170 97798 490226
rect 97854 490170 97922 490226
rect 97978 490170 98046 490226
rect 98102 490170 98198 490226
rect 97578 490102 98198 490170
rect 97578 490046 97674 490102
rect 97730 490046 97798 490102
rect 97854 490046 97922 490102
rect 97978 490046 98046 490102
rect 98102 490046 98198 490102
rect 97578 489978 98198 490046
rect 97578 489922 97674 489978
rect 97730 489922 97798 489978
rect 97854 489922 97922 489978
rect 97978 489922 98046 489978
rect 98102 489922 98198 489978
rect 82684 483364 82740 483374
rect 82684 483058 82740 483308
rect 82684 482992 82740 483002
rect 82236 482020 82292 482030
rect 80556 479332 80612 479342
rect 70578 478294 70674 478350
rect 70730 478294 70798 478350
rect 70854 478294 70922 478350
rect 70978 478294 71046 478350
rect 71102 478294 71198 478350
rect 70578 478226 71198 478294
rect 70578 478170 70674 478226
rect 70730 478170 70798 478226
rect 70854 478170 70922 478226
rect 70978 478170 71046 478226
rect 71102 478170 71198 478226
rect 70578 478102 71198 478170
rect 70578 478046 70674 478102
rect 70730 478046 70798 478102
rect 70854 478046 70922 478102
rect 70978 478046 71046 478102
rect 71102 478046 71198 478102
rect 70578 477978 71198 478046
rect 70578 477922 70674 477978
rect 70730 477922 70798 477978
rect 70854 477922 70922 477978
rect 70978 477922 71046 477978
rect 71102 477922 71198 477978
rect 69692 457762 69748 457772
rect 69804 473284 69860 473294
rect 66858 454294 66954 454350
rect 67010 454294 67078 454350
rect 67134 454294 67202 454350
rect 67258 454294 67326 454350
rect 67382 454294 67478 454350
rect 66858 454226 67478 454294
rect 66858 454170 66954 454226
rect 67010 454170 67078 454226
rect 67134 454170 67202 454226
rect 67258 454170 67326 454226
rect 67382 454170 67478 454226
rect 66858 454102 67478 454170
rect 66858 454046 66954 454102
rect 67010 454046 67078 454102
rect 67134 454046 67202 454102
rect 67258 454046 67326 454102
rect 67382 454046 67478 454102
rect 66858 453978 67478 454046
rect 66858 453922 66954 453978
rect 67010 453922 67078 453978
rect 67134 453922 67202 453978
rect 67258 453922 67326 453978
rect 67382 453922 67478 453978
rect 64988 441074 65044 441084
rect 64652 440962 64708 440972
rect 36138 436294 36234 436350
rect 36290 436294 36358 436350
rect 36414 436294 36482 436350
rect 36538 436294 36606 436350
rect 36662 436294 36758 436350
rect 36138 436226 36758 436294
rect 36138 436170 36234 436226
rect 36290 436170 36358 436226
rect 36414 436170 36482 436226
rect 36538 436170 36606 436226
rect 36662 436170 36758 436226
rect 36138 436102 36758 436170
rect 36138 436046 36234 436102
rect 36290 436046 36358 436102
rect 36414 436046 36482 436102
rect 36538 436046 36606 436102
rect 36662 436046 36758 436102
rect 36138 435978 36758 436046
rect 36138 435922 36234 435978
rect 36290 435922 36358 435978
rect 36414 435922 36482 435978
rect 36538 435922 36606 435978
rect 36662 435922 36758 435978
rect 24448 418350 24768 418384
rect 24448 418294 24518 418350
rect 24574 418294 24642 418350
rect 24698 418294 24768 418350
rect 24448 418226 24768 418294
rect 24448 418170 24518 418226
rect 24574 418170 24642 418226
rect 24698 418170 24768 418226
rect 24448 418102 24768 418170
rect 24448 418046 24518 418102
rect 24574 418046 24642 418102
rect 24698 418046 24768 418102
rect 24448 417978 24768 418046
rect 24448 417922 24518 417978
rect 24574 417922 24642 417978
rect 24698 417922 24768 417978
rect 24448 417888 24768 417922
rect 36138 418350 36758 435922
rect 66858 436350 67478 453922
rect 69804 439572 69860 473228
rect 69804 439506 69860 439516
rect 70578 460350 71198 477922
rect 73164 478660 73220 478670
rect 70578 460294 70674 460350
rect 70730 460294 70798 460350
rect 70854 460294 70922 460350
rect 70978 460294 71046 460350
rect 71102 460294 71198 460350
rect 70578 460226 71198 460294
rect 70578 460170 70674 460226
rect 70730 460170 70798 460226
rect 70854 460170 70922 460226
rect 70978 460170 71046 460226
rect 71102 460170 71198 460226
rect 70578 460102 71198 460170
rect 70578 460046 70674 460102
rect 70730 460046 70798 460102
rect 70854 460046 70922 460102
rect 70978 460046 71046 460102
rect 71102 460046 71198 460102
rect 70578 459978 71198 460046
rect 70578 459922 70674 459978
rect 70730 459922 70798 459978
rect 70854 459922 70922 459978
rect 70978 459922 71046 459978
rect 71102 459922 71198 459978
rect 70578 442350 71198 459922
rect 70578 442294 70674 442350
rect 70730 442294 70798 442350
rect 70854 442294 70922 442350
rect 70978 442294 71046 442350
rect 71102 442294 71198 442350
rect 70578 442226 71198 442294
rect 70578 442170 70674 442226
rect 70730 442170 70798 442226
rect 70854 442170 70922 442226
rect 70978 442170 71046 442226
rect 71102 442170 71198 442226
rect 70578 442102 71198 442170
rect 70578 442046 70674 442102
rect 70730 442046 70798 442102
rect 70854 442046 70922 442102
rect 70978 442046 71046 442102
rect 71102 442046 71198 442102
rect 70578 441978 71198 442046
rect 70578 441922 70674 441978
rect 70730 441922 70798 441978
rect 70854 441922 70922 441978
rect 70978 441922 71046 441978
rect 71102 441922 71198 441978
rect 66858 436294 66954 436350
rect 67010 436294 67078 436350
rect 67134 436294 67202 436350
rect 67258 436294 67326 436350
rect 67382 436294 67478 436350
rect 66858 436226 67478 436294
rect 66858 436170 66954 436226
rect 67010 436170 67078 436226
rect 67134 436170 67202 436226
rect 67258 436170 67326 436226
rect 67382 436170 67478 436226
rect 66858 436102 67478 436170
rect 66858 436046 66954 436102
rect 67010 436046 67078 436102
rect 67134 436046 67202 436102
rect 67258 436046 67326 436102
rect 67382 436046 67478 436102
rect 66858 435978 67478 436046
rect 66858 435922 66954 435978
rect 67010 435922 67078 435978
rect 67134 435922 67202 435978
rect 67258 435922 67326 435978
rect 67382 435922 67478 435978
rect 36138 418294 36234 418350
rect 36290 418294 36358 418350
rect 36414 418294 36482 418350
rect 36538 418294 36606 418350
rect 36662 418294 36758 418350
rect 36138 418226 36758 418294
rect 36138 418170 36234 418226
rect 36290 418170 36358 418226
rect 36414 418170 36482 418226
rect 36538 418170 36606 418226
rect 36662 418170 36758 418226
rect 36138 418102 36758 418170
rect 36138 418046 36234 418102
rect 36290 418046 36358 418102
rect 36414 418046 36482 418102
rect 36538 418046 36606 418102
rect 36662 418046 36758 418102
rect 36138 417978 36758 418046
rect 36138 417922 36234 417978
rect 36290 417922 36358 417978
rect 36414 417922 36482 417978
rect 36538 417922 36606 417978
rect 36662 417922 36758 417978
rect 18396 411796 18452 413162
rect 18396 411730 18452 411740
rect 19964 411684 20020 411694
rect 9138 406294 9234 406350
rect 9290 406294 9358 406350
rect 9414 406294 9482 406350
rect 9538 406294 9606 406350
rect 9662 406294 9758 406350
rect 9138 406226 9758 406294
rect 9138 406170 9234 406226
rect 9290 406170 9358 406226
rect 9414 406170 9482 406226
rect 9538 406170 9606 406226
rect 9662 406170 9758 406226
rect 9138 406102 9758 406170
rect 9138 406046 9234 406102
rect 9290 406046 9358 406102
rect 9414 406046 9482 406102
rect 9538 406046 9606 406102
rect 9662 406046 9758 406102
rect 9138 405978 9758 406046
rect 9138 405922 9234 405978
rect 9290 405922 9358 405978
rect 9414 405922 9482 405978
rect 9538 405922 9606 405978
rect 9662 405922 9758 405978
rect 9138 388350 9758 405922
rect 9138 388294 9234 388350
rect 9290 388294 9358 388350
rect 9414 388294 9482 388350
rect 9538 388294 9606 388350
rect 9662 388294 9758 388350
rect 9138 388226 9758 388294
rect 9138 388170 9234 388226
rect 9290 388170 9358 388226
rect 9414 388170 9482 388226
rect 9538 388170 9606 388226
rect 9662 388170 9758 388226
rect 9138 388102 9758 388170
rect 9138 388046 9234 388102
rect 9290 388046 9358 388102
rect 9414 388046 9482 388102
rect 9538 388046 9606 388102
rect 9662 388046 9758 388102
rect 9138 387978 9758 388046
rect 9138 387922 9234 387978
rect 9290 387922 9358 387978
rect 9414 387922 9482 387978
rect 9538 387922 9606 387978
rect 9662 387922 9758 387978
rect 9138 370350 9758 387922
rect 9138 370294 9234 370350
rect 9290 370294 9358 370350
rect 9414 370294 9482 370350
rect 9538 370294 9606 370350
rect 9662 370294 9758 370350
rect 9138 370226 9758 370294
rect 9138 370170 9234 370226
rect 9290 370170 9358 370226
rect 9414 370170 9482 370226
rect 9538 370170 9606 370226
rect 9662 370170 9758 370226
rect 9138 370102 9758 370170
rect 9138 370046 9234 370102
rect 9290 370046 9358 370102
rect 9414 370046 9482 370102
rect 9538 370046 9606 370102
rect 9662 370046 9758 370102
rect 9138 369978 9758 370046
rect 9138 369922 9234 369978
rect 9290 369922 9358 369978
rect 9414 369922 9482 369978
rect 9538 369922 9606 369978
rect 9662 369922 9758 369978
rect 9138 352350 9758 369922
rect 18060 411460 18116 411470
rect 18060 361956 18116 411404
rect 19852 410788 19908 410798
rect 19740 410116 19796 410126
rect 18284 408100 18340 408110
rect 18172 401380 18228 401390
rect 18172 378980 18228 401324
rect 18172 378914 18228 378924
rect 18284 362516 18340 408044
rect 19740 378868 19796 410060
rect 19852 386596 19908 410732
rect 19852 386530 19908 386540
rect 19964 384916 20020 411628
rect 20636 406756 20692 406776
rect 20636 406672 20692 406682
rect 20076 402724 20132 402734
rect 20076 388052 20132 402668
rect 24448 400350 24768 400384
rect 24448 400294 24518 400350
rect 24574 400294 24642 400350
rect 24698 400294 24768 400350
rect 24448 400226 24768 400294
rect 24448 400170 24518 400226
rect 24574 400170 24642 400226
rect 24698 400170 24768 400226
rect 24448 400102 24768 400170
rect 24448 400046 24518 400102
rect 24574 400046 24642 400102
rect 24698 400046 24768 400102
rect 24448 399978 24768 400046
rect 24448 399922 24518 399978
rect 24574 399922 24642 399978
rect 24698 399922 24768 399978
rect 24448 399888 24768 399922
rect 36138 400350 36758 417922
rect 55168 418350 55488 418384
rect 55168 418294 55238 418350
rect 55294 418294 55362 418350
rect 55418 418294 55488 418350
rect 55168 418226 55488 418294
rect 55168 418170 55238 418226
rect 55294 418170 55362 418226
rect 55418 418170 55488 418226
rect 55168 418102 55488 418170
rect 55168 418046 55238 418102
rect 55294 418046 55362 418102
rect 55418 418046 55488 418102
rect 55168 417978 55488 418046
rect 55168 417922 55238 417978
rect 55294 417922 55362 417978
rect 55418 417922 55488 417978
rect 55168 417888 55488 417922
rect 66858 418350 67478 435922
rect 66858 418294 66954 418350
rect 67010 418294 67078 418350
rect 67134 418294 67202 418350
rect 67258 418294 67326 418350
rect 67382 418294 67478 418350
rect 66858 418226 67478 418294
rect 66858 418170 66954 418226
rect 67010 418170 67078 418226
rect 67134 418170 67202 418226
rect 67258 418170 67326 418226
rect 67382 418170 67478 418226
rect 66858 418102 67478 418170
rect 66858 418046 66954 418102
rect 67010 418046 67078 418102
rect 67134 418046 67202 418102
rect 67258 418046 67326 418102
rect 67382 418046 67478 418102
rect 66858 417978 67478 418046
rect 66858 417922 66954 417978
rect 67010 417922 67078 417978
rect 67134 417922 67202 417978
rect 67258 417922 67326 417978
rect 67382 417922 67478 417978
rect 62972 406738 63028 406748
rect 39808 406350 40128 406384
rect 39808 406294 39878 406350
rect 39934 406294 40002 406350
rect 40058 406294 40128 406350
rect 39808 406226 40128 406294
rect 39808 406170 39878 406226
rect 39934 406170 40002 406226
rect 40058 406170 40128 406226
rect 39808 406102 40128 406170
rect 39808 406046 39878 406102
rect 39934 406046 40002 406102
rect 40058 406046 40128 406102
rect 39808 405978 40128 406046
rect 39808 405922 39878 405978
rect 39934 405922 40002 405978
rect 40058 405922 40128 405978
rect 39808 405888 40128 405922
rect 36138 400294 36234 400350
rect 36290 400294 36358 400350
rect 36414 400294 36482 400350
rect 36538 400294 36606 400350
rect 36662 400294 36758 400350
rect 36138 400226 36758 400294
rect 36138 400170 36234 400226
rect 36290 400170 36358 400226
rect 36414 400170 36482 400226
rect 36538 400170 36606 400226
rect 36662 400170 36758 400226
rect 36138 400102 36758 400170
rect 36138 400046 36234 400102
rect 36290 400046 36358 400102
rect 36414 400046 36482 400102
rect 36538 400046 36606 400102
rect 36662 400046 36758 400102
rect 36138 399978 36758 400046
rect 36138 399922 36234 399978
rect 36290 399922 36358 399978
rect 36414 399922 36482 399978
rect 36538 399922 36606 399978
rect 36662 399922 36758 399978
rect 20076 387986 20132 387996
rect 19964 384850 20020 384860
rect 19740 378802 19796 378812
rect 36138 382350 36758 399922
rect 55168 400350 55488 400384
rect 55168 400294 55238 400350
rect 55294 400294 55362 400350
rect 55418 400294 55488 400350
rect 55168 400226 55488 400294
rect 55168 400170 55238 400226
rect 55294 400170 55362 400226
rect 55418 400170 55488 400226
rect 55168 400102 55488 400170
rect 55168 400046 55238 400102
rect 55294 400046 55362 400102
rect 55418 400046 55488 400102
rect 55168 399978 55488 400046
rect 55168 399922 55238 399978
rect 55294 399922 55362 399978
rect 55418 399922 55488 399978
rect 55168 399888 55488 399922
rect 62972 391438 63028 406682
rect 62972 391372 63028 391382
rect 64652 406084 64708 406094
rect 39808 388389 40128 388446
rect 39808 388333 39836 388389
rect 39892 388333 39940 388389
rect 39996 388333 40044 388389
rect 40100 388333 40128 388389
rect 39808 388276 40128 388333
rect 36138 382294 36234 382350
rect 36290 382294 36358 382350
rect 36414 382294 36482 382350
rect 36538 382294 36606 382350
rect 36662 382294 36758 382350
rect 36138 382226 36758 382294
rect 36138 382170 36234 382226
rect 36290 382170 36358 382226
rect 36414 382170 36482 382226
rect 36538 382170 36606 382226
rect 36662 382170 36758 382226
rect 36138 382102 36758 382170
rect 36138 382046 36234 382102
rect 36290 382046 36358 382102
rect 36414 382046 36482 382102
rect 36538 382046 36606 382102
rect 36662 382046 36758 382102
rect 36138 381978 36758 382046
rect 36138 381922 36234 381978
rect 36290 381922 36358 381978
rect 36414 381922 36482 381978
rect 36538 381922 36606 381978
rect 36662 381922 36758 381978
rect 18284 362450 18340 362460
rect 36138 364350 36758 381922
rect 36138 364294 36234 364350
rect 36290 364294 36358 364350
rect 36414 364294 36482 364350
rect 36538 364294 36606 364350
rect 36662 364294 36758 364350
rect 36138 364226 36758 364294
rect 36138 364170 36234 364226
rect 36290 364170 36358 364226
rect 36414 364170 36482 364226
rect 36538 364170 36606 364226
rect 36662 364170 36758 364226
rect 36138 364102 36758 364170
rect 36138 364046 36234 364102
rect 36290 364046 36358 364102
rect 36414 364046 36482 364102
rect 36538 364046 36606 364102
rect 36662 364046 36758 364102
rect 36138 363978 36758 364046
rect 36138 363922 36234 363978
rect 36290 363922 36358 363978
rect 36414 363922 36482 363978
rect 36538 363922 36606 363978
rect 36662 363922 36758 363978
rect 18060 361890 18116 361900
rect 9138 352294 9234 352350
rect 9290 352294 9358 352350
rect 9414 352294 9482 352350
rect 9538 352294 9606 352350
rect 9662 352294 9758 352350
rect 9138 352226 9758 352294
rect 9138 352170 9234 352226
rect 9290 352170 9358 352226
rect 9414 352170 9482 352226
rect 9538 352170 9606 352226
rect 9662 352170 9758 352226
rect 9138 352102 9758 352170
rect 9138 352046 9234 352102
rect 9290 352046 9358 352102
rect 9414 352046 9482 352102
rect 9538 352046 9606 352102
rect 9662 352046 9758 352102
rect 9138 351978 9758 352046
rect 9138 351922 9234 351978
rect 9290 351922 9358 351978
rect 9414 351922 9482 351978
rect 9538 351922 9606 351978
rect 9662 351922 9758 351978
rect 9138 334350 9758 351922
rect 24448 346350 24768 346384
rect 24448 346294 24518 346350
rect 24574 346294 24642 346350
rect 24698 346294 24768 346350
rect 24448 346226 24768 346294
rect 24448 346170 24518 346226
rect 24574 346170 24642 346226
rect 24698 346170 24768 346226
rect 24448 346102 24768 346170
rect 24448 346046 24518 346102
rect 24574 346046 24642 346102
rect 24698 346046 24768 346102
rect 24448 345978 24768 346046
rect 24448 345922 24518 345978
rect 24574 345922 24642 345978
rect 24698 345922 24768 345978
rect 24448 345888 24768 345922
rect 36138 346350 36758 363922
rect 64652 359716 64708 406028
rect 64876 401380 64932 401390
rect 64876 360276 64932 401324
rect 64876 360210 64932 360220
rect 66858 400350 67478 417922
rect 70578 424350 71198 441922
rect 73052 472612 73108 472622
rect 73052 434308 73108 472556
rect 73164 446516 73220 478604
rect 80332 478660 80388 478670
rect 73164 446450 73220 446460
rect 78316 476644 78372 476654
rect 78316 445956 78372 476588
rect 80332 452900 80388 478604
rect 80332 452834 80388 452844
rect 80444 476644 80500 476654
rect 78316 445890 78372 445900
rect 73052 434242 73108 434252
rect 80444 432628 80500 476588
rect 80556 434420 80612 479276
rect 82124 473956 82180 473966
rect 81452 465220 81508 465230
rect 81452 444276 81508 465164
rect 82012 461188 82068 461198
rect 82012 456148 82068 461132
rect 82012 456082 82068 456092
rect 82124 451556 82180 473900
rect 82124 451490 82180 451500
rect 81452 444210 81508 444220
rect 80556 434354 80612 434364
rect 80444 432562 80500 432572
rect 82236 426580 82292 481964
rect 97578 480894 98198 489922
rect 117168 490350 117488 490384
rect 117168 490294 117238 490350
rect 117294 490294 117362 490350
rect 117418 490294 117488 490350
rect 117168 490226 117488 490294
rect 117168 490170 117238 490226
rect 117294 490170 117362 490226
rect 117418 490170 117488 490226
rect 117168 490102 117488 490170
rect 117168 490046 117238 490102
rect 117294 490046 117362 490102
rect 117418 490046 117488 490102
rect 117168 489978 117488 490046
rect 117168 489922 117238 489978
rect 117294 489922 117362 489978
rect 117418 489922 117488 489978
rect 117168 489888 117488 489922
rect 128298 490350 128918 507922
rect 128298 490294 128394 490350
rect 128450 490294 128518 490350
rect 128574 490294 128642 490350
rect 128698 490294 128766 490350
rect 128822 490294 128918 490350
rect 128298 490226 128918 490294
rect 128298 490170 128394 490226
rect 128450 490170 128518 490226
rect 128574 490170 128642 490226
rect 128698 490170 128766 490226
rect 128822 490170 128918 490226
rect 128298 490102 128918 490170
rect 128298 490046 128394 490102
rect 128450 490046 128518 490102
rect 128574 490046 128642 490102
rect 128698 490046 128766 490102
rect 128822 490046 128918 490102
rect 128298 489978 128918 490046
rect 128298 489922 128394 489978
rect 128450 489922 128518 489978
rect 128574 489922 128642 489978
rect 128698 489922 128766 489978
rect 128822 489922 128918 489978
rect 127596 482020 127652 482030
rect 127596 480452 127652 481964
rect 127596 480386 127652 480396
rect 127596 478660 127652 478670
rect 101808 478350 102128 478384
rect 101808 478294 101878 478350
rect 101934 478294 102002 478350
rect 102058 478294 102128 478350
rect 101808 478226 102128 478294
rect 101808 478170 101878 478226
rect 101934 478170 102002 478226
rect 102058 478170 102128 478226
rect 101808 478102 102128 478170
rect 101808 478046 101878 478102
rect 101934 478046 102002 478102
rect 102058 478046 102128 478102
rect 101808 477978 102128 478046
rect 101808 477922 101878 477978
rect 101934 477922 102002 477978
rect 102058 477922 102128 477978
rect 101808 477888 102128 477922
rect 127596 476308 127652 478604
rect 127596 476242 127652 476252
rect 126812 474628 126868 474638
rect 86448 472350 86768 472384
rect 86448 472294 86518 472350
rect 86574 472294 86642 472350
rect 86698 472294 86768 472350
rect 86448 472226 86768 472294
rect 86448 472170 86518 472226
rect 86574 472170 86642 472226
rect 86698 472170 86768 472226
rect 86448 472102 86768 472170
rect 86448 472046 86518 472102
rect 86574 472046 86642 472102
rect 86698 472046 86768 472102
rect 86448 471978 86768 472046
rect 86448 471922 86518 471978
rect 86574 471922 86642 471978
rect 86698 471922 86768 471978
rect 86448 471888 86768 471922
rect 97578 472350 98198 473234
rect 97578 472294 97674 472350
rect 97730 472294 97798 472350
rect 97854 472294 97922 472350
rect 97978 472294 98046 472350
rect 98102 472294 98198 472350
rect 97578 472226 98198 472294
rect 97578 472170 97674 472226
rect 97730 472170 97798 472226
rect 97854 472170 97922 472226
rect 97978 472170 98046 472226
rect 98102 472170 98198 472226
rect 97578 472102 98198 472170
rect 97578 472046 97674 472102
rect 97730 472046 97798 472102
rect 97854 472046 97922 472102
rect 97978 472046 98046 472102
rect 98102 472046 98198 472102
rect 97578 471978 98198 472046
rect 97578 471922 97674 471978
rect 97730 471922 97798 471978
rect 97854 471922 97922 471978
rect 97978 471922 98046 471978
rect 98102 471922 98198 471978
rect 82236 426514 82292 426524
rect 97578 454350 98198 471922
rect 117168 472350 117488 472384
rect 117168 472294 117238 472350
rect 117294 472294 117362 472350
rect 117418 472294 117488 472350
rect 117168 472226 117488 472294
rect 117168 472170 117238 472226
rect 117294 472170 117362 472226
rect 117418 472170 117488 472226
rect 117168 472102 117488 472170
rect 117168 472046 117238 472102
rect 117294 472046 117362 472102
rect 117418 472046 117488 472102
rect 117168 471978 117488 472046
rect 117168 471922 117238 471978
rect 117294 471922 117362 471978
rect 117418 471922 117488 471978
rect 117168 471888 117488 471922
rect 101808 460350 102128 460384
rect 101808 460294 101878 460350
rect 101934 460294 102002 460350
rect 102058 460294 102128 460350
rect 101808 460226 102128 460294
rect 101808 460170 101878 460226
rect 101934 460170 102002 460226
rect 102058 460170 102128 460226
rect 101808 460102 102128 460170
rect 101808 460046 101878 460102
rect 101934 460046 102002 460102
rect 102058 460046 102128 460102
rect 101808 459978 102128 460046
rect 101808 459922 101878 459978
rect 101934 459922 102002 459978
rect 102058 459922 102128 459978
rect 101808 459888 102128 459922
rect 97578 454294 97674 454350
rect 97730 454294 97798 454350
rect 97854 454294 97922 454350
rect 97978 454294 98046 454350
rect 98102 454294 98198 454350
rect 97578 454226 98198 454294
rect 97578 454170 97674 454226
rect 97730 454170 97798 454226
rect 97854 454170 97922 454226
rect 97978 454170 98046 454226
rect 98102 454170 98198 454226
rect 97578 454102 98198 454170
rect 97578 454046 97674 454102
rect 97730 454046 97798 454102
rect 97854 454046 97922 454102
rect 97978 454046 98046 454102
rect 98102 454046 98198 454102
rect 97578 453978 98198 454046
rect 97578 453922 97674 453978
rect 97730 453922 97798 453978
rect 97854 453922 97922 453978
rect 97978 453922 98046 453978
rect 98102 453922 98198 453978
rect 97578 436350 98198 453922
rect 126812 438004 126868 474572
rect 127036 473956 127092 473966
rect 127036 446068 127092 473900
rect 127036 446002 127092 446012
rect 128298 472350 128918 489922
rect 132018 598172 132638 598268
rect 132018 598116 132114 598172
rect 132170 598116 132238 598172
rect 132294 598116 132362 598172
rect 132418 598116 132486 598172
rect 132542 598116 132638 598172
rect 132018 598048 132638 598116
rect 132018 597992 132114 598048
rect 132170 597992 132238 598048
rect 132294 597992 132362 598048
rect 132418 597992 132486 598048
rect 132542 597992 132638 598048
rect 132018 597924 132638 597992
rect 132018 597868 132114 597924
rect 132170 597868 132238 597924
rect 132294 597868 132362 597924
rect 132418 597868 132486 597924
rect 132542 597868 132638 597924
rect 132018 597800 132638 597868
rect 132018 597744 132114 597800
rect 132170 597744 132238 597800
rect 132294 597744 132362 597800
rect 132418 597744 132486 597800
rect 132542 597744 132638 597800
rect 132018 586350 132638 597744
rect 132018 586294 132114 586350
rect 132170 586294 132238 586350
rect 132294 586294 132362 586350
rect 132418 586294 132486 586350
rect 132542 586294 132638 586350
rect 132018 586226 132638 586294
rect 132018 586170 132114 586226
rect 132170 586170 132238 586226
rect 132294 586170 132362 586226
rect 132418 586170 132486 586226
rect 132542 586170 132638 586226
rect 132018 586102 132638 586170
rect 132018 586046 132114 586102
rect 132170 586046 132238 586102
rect 132294 586046 132362 586102
rect 132418 586046 132486 586102
rect 132542 586046 132638 586102
rect 132018 585978 132638 586046
rect 132018 585922 132114 585978
rect 132170 585922 132238 585978
rect 132294 585922 132362 585978
rect 132418 585922 132486 585978
rect 132542 585922 132638 585978
rect 132018 568350 132638 585922
rect 132018 568294 132114 568350
rect 132170 568294 132238 568350
rect 132294 568294 132362 568350
rect 132418 568294 132486 568350
rect 132542 568294 132638 568350
rect 132018 568226 132638 568294
rect 132018 568170 132114 568226
rect 132170 568170 132238 568226
rect 132294 568170 132362 568226
rect 132418 568170 132486 568226
rect 132542 568170 132638 568226
rect 132018 568102 132638 568170
rect 132018 568046 132114 568102
rect 132170 568046 132238 568102
rect 132294 568046 132362 568102
rect 132418 568046 132486 568102
rect 132542 568046 132638 568102
rect 132018 567978 132638 568046
rect 132018 567922 132114 567978
rect 132170 567922 132238 567978
rect 132294 567922 132362 567978
rect 132418 567922 132486 567978
rect 132542 567922 132638 567978
rect 132018 550350 132638 567922
rect 159018 597212 159638 598268
rect 159018 597156 159114 597212
rect 159170 597156 159238 597212
rect 159294 597156 159362 597212
rect 159418 597156 159486 597212
rect 159542 597156 159638 597212
rect 159018 597088 159638 597156
rect 159018 597032 159114 597088
rect 159170 597032 159238 597088
rect 159294 597032 159362 597088
rect 159418 597032 159486 597088
rect 159542 597032 159638 597088
rect 159018 596964 159638 597032
rect 159018 596908 159114 596964
rect 159170 596908 159238 596964
rect 159294 596908 159362 596964
rect 159418 596908 159486 596964
rect 159542 596908 159638 596964
rect 159018 596840 159638 596908
rect 159018 596784 159114 596840
rect 159170 596784 159238 596840
rect 159294 596784 159362 596840
rect 159418 596784 159486 596840
rect 159542 596784 159638 596840
rect 159018 580350 159638 596784
rect 159018 580294 159114 580350
rect 159170 580294 159238 580350
rect 159294 580294 159362 580350
rect 159418 580294 159486 580350
rect 159542 580294 159638 580350
rect 159018 580226 159638 580294
rect 159018 580170 159114 580226
rect 159170 580170 159238 580226
rect 159294 580170 159362 580226
rect 159418 580170 159486 580226
rect 159542 580170 159638 580226
rect 159018 580102 159638 580170
rect 159018 580046 159114 580102
rect 159170 580046 159238 580102
rect 159294 580046 159362 580102
rect 159418 580046 159486 580102
rect 159542 580046 159638 580102
rect 159018 579978 159638 580046
rect 159018 579922 159114 579978
rect 159170 579922 159238 579978
rect 159294 579922 159362 579978
rect 159418 579922 159486 579978
rect 159542 579922 159638 579978
rect 141036 564004 141092 564014
rect 141036 556164 141092 563948
rect 148448 562350 148768 562384
rect 148448 562294 148518 562350
rect 148574 562294 148642 562350
rect 148698 562294 148768 562350
rect 148448 562226 148768 562294
rect 148448 562170 148518 562226
rect 148574 562170 148642 562226
rect 148698 562170 148768 562226
rect 148448 562102 148768 562170
rect 148448 562046 148518 562102
rect 148574 562046 148642 562102
rect 148698 562046 148768 562102
rect 148448 561978 148768 562046
rect 148448 561922 148518 561978
rect 148574 561922 148642 561978
rect 148698 561922 148768 561978
rect 148448 561888 148768 561922
rect 159018 562350 159638 579922
rect 159018 562294 159114 562350
rect 159170 562294 159238 562350
rect 159294 562294 159362 562350
rect 159418 562294 159486 562350
rect 159542 562294 159638 562350
rect 159018 562226 159638 562294
rect 159018 562170 159114 562226
rect 159170 562170 159238 562226
rect 159294 562170 159362 562226
rect 159418 562170 159486 562226
rect 159542 562170 159638 562226
rect 159018 562102 159638 562170
rect 159018 562046 159114 562102
rect 159170 562046 159238 562102
rect 159294 562046 159362 562102
rect 159418 562046 159486 562102
rect 159542 562046 159638 562102
rect 159018 561978 159638 562046
rect 159018 561922 159114 561978
rect 159170 561922 159238 561978
rect 159294 561922 159362 561978
rect 159418 561922 159486 561978
rect 159542 561922 159638 561978
rect 141036 556098 141092 556108
rect 141932 556164 141988 556174
rect 141036 555940 141092 555950
rect 141036 554518 141092 555884
rect 141036 554452 141092 554462
rect 141036 551908 141092 551918
rect 132018 550294 132114 550350
rect 132170 550294 132238 550350
rect 132294 550294 132362 550350
rect 132418 550294 132486 550350
rect 132542 550294 132638 550350
rect 132018 550226 132638 550294
rect 132018 550170 132114 550226
rect 132170 550170 132238 550226
rect 132294 550170 132362 550226
rect 132418 550170 132486 550226
rect 132542 550170 132638 550226
rect 132018 550102 132638 550170
rect 132018 550046 132114 550102
rect 132170 550046 132238 550102
rect 132294 550046 132362 550102
rect 132418 550046 132486 550102
rect 132542 550046 132638 550102
rect 132018 549978 132638 550046
rect 132018 549922 132114 549978
rect 132170 549922 132238 549978
rect 132294 549922 132362 549978
rect 132418 549922 132486 549978
rect 132542 549922 132638 549978
rect 132018 532350 132638 549922
rect 140924 551236 140980 551246
rect 132018 532294 132114 532350
rect 132170 532294 132238 532350
rect 132294 532294 132362 532350
rect 132418 532294 132486 532350
rect 132542 532294 132638 532350
rect 132018 532226 132638 532294
rect 132018 532170 132114 532226
rect 132170 532170 132238 532226
rect 132294 532170 132362 532226
rect 132418 532170 132486 532226
rect 132542 532170 132638 532226
rect 132018 532102 132638 532170
rect 132018 532046 132114 532102
rect 132170 532046 132238 532102
rect 132294 532046 132362 532102
rect 132418 532046 132486 532102
rect 132542 532046 132638 532102
rect 132018 531978 132638 532046
rect 132018 531922 132114 531978
rect 132170 531922 132238 531978
rect 132294 531922 132362 531978
rect 132418 531922 132486 531978
rect 132542 531922 132638 531978
rect 132018 514350 132638 531922
rect 132018 514294 132114 514350
rect 132170 514294 132238 514350
rect 132294 514294 132362 514350
rect 132418 514294 132486 514350
rect 132542 514294 132638 514350
rect 132018 514226 132638 514294
rect 132018 514170 132114 514226
rect 132170 514170 132238 514226
rect 132294 514170 132362 514226
rect 132418 514170 132486 514226
rect 132542 514170 132638 514226
rect 132018 514102 132638 514170
rect 132018 514046 132114 514102
rect 132170 514046 132238 514102
rect 132294 514046 132362 514102
rect 132418 514046 132486 514102
rect 132542 514046 132638 514102
rect 132018 513978 132638 514046
rect 132018 513922 132114 513978
rect 132170 513922 132238 513978
rect 132294 513922 132362 513978
rect 132418 513922 132486 513978
rect 132542 513922 132638 513978
rect 132018 496350 132638 513922
rect 138572 545188 138628 545198
rect 138572 509236 138628 545132
rect 140812 545188 140868 545198
rect 140812 530292 140868 545132
rect 140812 530226 140868 530236
rect 140924 529172 140980 551180
rect 141036 546084 141092 551852
rect 141036 546018 141092 546028
rect 140924 529106 140980 529116
rect 141036 544516 141092 544526
rect 141036 511700 141092 544460
rect 141932 516516 141988 556108
rect 144060 555268 144116 555278
rect 144060 555172 144116 555182
rect 143612 548548 143668 548558
rect 141932 516450 141988 516460
rect 142044 546532 142100 546542
rect 142044 514836 142100 546476
rect 142716 543172 142772 543182
rect 142716 520436 142772 543116
rect 142716 520370 142772 520380
rect 142044 514770 142100 514780
rect 141036 511634 141092 511644
rect 138572 509170 138628 509180
rect 143612 508676 143668 548492
rect 143724 546084 143780 546094
rect 143724 519876 143780 546028
rect 148448 544350 148768 544384
rect 148448 544294 148518 544350
rect 148574 544294 148642 544350
rect 148698 544294 148768 544350
rect 148448 544226 148768 544294
rect 148448 544170 148518 544226
rect 148574 544170 148642 544226
rect 148698 544170 148768 544226
rect 148448 544102 148768 544170
rect 148448 544046 148518 544102
rect 148574 544046 148642 544102
rect 148698 544046 148768 544102
rect 148448 543978 148768 544046
rect 148448 543922 148518 543978
rect 148574 543922 148642 543978
rect 148698 543922 148768 543978
rect 148448 543888 148768 543922
rect 159018 544350 159638 561922
rect 162738 598172 163358 598268
rect 162738 598116 162834 598172
rect 162890 598116 162958 598172
rect 163014 598116 163082 598172
rect 163138 598116 163206 598172
rect 163262 598116 163358 598172
rect 162738 598048 163358 598116
rect 162738 597992 162834 598048
rect 162890 597992 162958 598048
rect 163014 597992 163082 598048
rect 163138 597992 163206 598048
rect 163262 597992 163358 598048
rect 162738 597924 163358 597992
rect 162738 597868 162834 597924
rect 162890 597868 162958 597924
rect 163014 597868 163082 597924
rect 163138 597868 163206 597924
rect 163262 597868 163358 597924
rect 162738 597800 163358 597868
rect 162738 597744 162834 597800
rect 162890 597744 162958 597800
rect 163014 597744 163082 597800
rect 163138 597744 163206 597800
rect 163262 597744 163358 597800
rect 162738 586350 163358 597744
rect 162738 586294 162834 586350
rect 162890 586294 162958 586350
rect 163014 586294 163082 586350
rect 163138 586294 163206 586350
rect 163262 586294 163358 586350
rect 162738 586226 163358 586294
rect 162738 586170 162834 586226
rect 162890 586170 162958 586226
rect 163014 586170 163082 586226
rect 163138 586170 163206 586226
rect 163262 586170 163358 586226
rect 162738 586102 163358 586170
rect 162738 586046 162834 586102
rect 162890 586046 162958 586102
rect 163014 586046 163082 586102
rect 163138 586046 163206 586102
rect 163262 586046 163358 586102
rect 162738 585978 163358 586046
rect 162738 585922 162834 585978
rect 162890 585922 162958 585978
rect 163014 585922 163082 585978
rect 163138 585922 163206 585978
rect 163262 585922 163358 585978
rect 162738 568350 163358 585922
rect 162738 568294 162834 568350
rect 162890 568294 162958 568350
rect 163014 568294 163082 568350
rect 163138 568294 163206 568350
rect 163262 568294 163358 568350
rect 162738 568226 163358 568294
rect 162738 568170 162834 568226
rect 162890 568170 162958 568226
rect 163014 568170 163082 568226
rect 163138 568170 163206 568226
rect 163262 568170 163358 568226
rect 162738 568102 163358 568170
rect 162738 568046 162834 568102
rect 162890 568046 162958 568102
rect 163014 568046 163082 568102
rect 163138 568046 163206 568102
rect 163262 568046 163358 568102
rect 162738 567978 163358 568046
rect 162738 567922 162834 567978
rect 162890 567922 162958 567978
rect 163014 567922 163082 567978
rect 163138 567922 163206 567978
rect 163262 567922 163358 567978
rect 162738 553886 163358 567922
rect 189738 597212 190358 598268
rect 189738 597156 189834 597212
rect 189890 597156 189958 597212
rect 190014 597156 190082 597212
rect 190138 597156 190206 597212
rect 190262 597156 190358 597212
rect 189738 597088 190358 597156
rect 189738 597032 189834 597088
rect 189890 597032 189958 597088
rect 190014 597032 190082 597088
rect 190138 597032 190206 597088
rect 190262 597032 190358 597088
rect 189738 596964 190358 597032
rect 189738 596908 189834 596964
rect 189890 596908 189958 596964
rect 190014 596908 190082 596964
rect 190138 596908 190206 596964
rect 190262 596908 190358 596964
rect 189738 596840 190358 596908
rect 189738 596784 189834 596840
rect 189890 596784 189958 596840
rect 190014 596784 190082 596840
rect 190138 596784 190206 596840
rect 190262 596784 190358 596840
rect 189738 580350 190358 596784
rect 189738 580294 189834 580350
rect 189890 580294 189958 580350
rect 190014 580294 190082 580350
rect 190138 580294 190206 580350
rect 190262 580294 190358 580350
rect 189738 580226 190358 580294
rect 189738 580170 189834 580226
rect 189890 580170 189958 580226
rect 190014 580170 190082 580226
rect 190138 580170 190206 580226
rect 190262 580170 190358 580226
rect 189738 580102 190358 580170
rect 189738 580046 189834 580102
rect 189890 580046 189958 580102
rect 190014 580046 190082 580102
rect 190138 580046 190206 580102
rect 190262 580046 190358 580102
rect 189738 579978 190358 580046
rect 189738 579922 189834 579978
rect 189890 579922 189958 579978
rect 190014 579922 190082 579978
rect 190138 579922 190206 579978
rect 190262 579922 190358 579978
rect 179168 562350 179488 562384
rect 179168 562294 179238 562350
rect 179294 562294 179362 562350
rect 179418 562294 179488 562350
rect 179168 562226 179488 562294
rect 179168 562170 179238 562226
rect 179294 562170 179362 562226
rect 179418 562170 179488 562226
rect 179168 562102 179488 562170
rect 179168 562046 179238 562102
rect 179294 562046 179362 562102
rect 179418 562046 179488 562102
rect 179168 561978 179488 562046
rect 179168 561922 179238 561978
rect 179294 561922 179362 561978
rect 179418 561922 179488 561978
rect 179168 561888 179488 561922
rect 189738 562350 190358 579922
rect 189738 562294 189834 562350
rect 189890 562294 189958 562350
rect 190014 562294 190082 562350
rect 190138 562294 190206 562350
rect 190262 562294 190358 562350
rect 189738 562226 190358 562294
rect 189738 562170 189834 562226
rect 189890 562170 189958 562226
rect 190014 562170 190082 562226
rect 190138 562170 190206 562226
rect 190262 562170 190358 562226
rect 189738 562102 190358 562170
rect 189738 562046 189834 562102
rect 189890 562046 189958 562102
rect 190014 562046 190082 562102
rect 190138 562046 190206 562102
rect 190262 562046 190358 562102
rect 189738 561978 190358 562046
rect 189738 561922 189834 561978
rect 189890 561922 189958 561978
rect 190014 561922 190082 561978
rect 190138 561922 190206 561978
rect 190262 561922 190358 561978
rect 189084 551236 189140 551246
rect 163808 550350 164128 550384
rect 163808 550294 163878 550350
rect 163934 550294 164002 550350
rect 164058 550294 164128 550350
rect 163808 550226 164128 550294
rect 163808 550170 163878 550226
rect 163934 550170 164002 550226
rect 164058 550170 164128 550226
rect 163808 550102 164128 550170
rect 163808 550046 163878 550102
rect 163934 550046 164002 550102
rect 164058 550046 164128 550102
rect 163808 549978 164128 550046
rect 163808 549922 163878 549978
rect 163934 549922 164002 549978
rect 164058 549922 164128 549978
rect 163808 549888 164128 549922
rect 188972 549892 189028 549902
rect 159018 544294 159114 544350
rect 159170 544294 159238 544350
rect 159294 544294 159362 544350
rect 159418 544294 159486 544350
rect 159542 544294 159638 544350
rect 159018 544226 159638 544294
rect 159018 544170 159114 544226
rect 159170 544170 159238 544226
rect 159294 544170 159362 544226
rect 159418 544170 159486 544226
rect 159542 544170 159638 544226
rect 159018 544102 159638 544170
rect 159018 544046 159114 544102
rect 159170 544046 159238 544102
rect 159294 544046 159362 544102
rect 159418 544046 159486 544102
rect 159542 544046 159638 544102
rect 159018 543978 159638 544046
rect 159018 543922 159114 543978
rect 159170 543922 159238 543978
rect 159294 543922 159362 543978
rect 159418 543922 159486 543978
rect 159542 543922 159638 543978
rect 146076 529172 146132 529182
rect 146076 523236 146132 529116
rect 146076 523170 146132 523180
rect 159018 526350 159638 543922
rect 179168 544350 179488 544384
rect 179168 544294 179238 544350
rect 179294 544294 179362 544350
rect 179418 544294 179488 544350
rect 179168 544226 179488 544294
rect 179168 544170 179238 544226
rect 179294 544170 179362 544226
rect 179418 544170 179488 544226
rect 179168 544102 179488 544170
rect 179168 544046 179238 544102
rect 179294 544046 179362 544102
rect 179418 544046 179488 544102
rect 179168 543978 179488 544046
rect 179168 543922 179238 543978
rect 179294 543922 179362 543978
rect 179418 543922 179488 543978
rect 179168 543888 179488 543922
rect 159018 526294 159114 526350
rect 159170 526294 159238 526350
rect 159294 526294 159362 526350
rect 159418 526294 159486 526350
rect 159542 526294 159638 526350
rect 159018 526226 159638 526294
rect 159018 526170 159114 526226
rect 159170 526170 159238 526226
rect 159294 526170 159362 526226
rect 159418 526170 159486 526226
rect 159542 526170 159638 526226
rect 159018 526102 159638 526170
rect 159018 526046 159114 526102
rect 159170 526046 159238 526102
rect 159294 526046 159362 526102
rect 159418 526046 159486 526102
rect 159542 526046 159638 526102
rect 159018 525978 159638 526046
rect 159018 525922 159114 525978
rect 159170 525922 159238 525978
rect 159294 525922 159362 525978
rect 159418 525922 159486 525978
rect 159542 525922 159638 525978
rect 143724 519810 143780 519820
rect 143612 508610 143668 508620
rect 132018 496294 132114 496350
rect 132170 496294 132238 496350
rect 132294 496294 132362 496350
rect 132418 496294 132486 496350
rect 132542 496294 132638 496350
rect 132018 496226 132638 496294
rect 132018 496170 132114 496226
rect 132170 496170 132238 496226
rect 132294 496170 132362 496226
rect 132418 496170 132486 496226
rect 132542 496170 132638 496226
rect 132018 496102 132638 496170
rect 132018 496046 132114 496102
rect 132170 496046 132238 496102
rect 132294 496046 132362 496102
rect 132418 496046 132486 496102
rect 132542 496046 132638 496102
rect 132018 495978 132638 496046
rect 132018 495922 132114 495978
rect 132170 495922 132238 495978
rect 132294 495922 132362 495978
rect 132418 495922 132486 495978
rect 132542 495922 132638 495978
rect 128298 472294 128394 472350
rect 128450 472294 128518 472350
rect 128574 472294 128642 472350
rect 128698 472294 128766 472350
rect 128822 472294 128918 472350
rect 128298 472226 128918 472294
rect 128298 472170 128394 472226
rect 128450 472170 128518 472226
rect 128574 472170 128642 472226
rect 128698 472170 128766 472226
rect 128822 472170 128918 472226
rect 128298 472102 128918 472170
rect 128298 472046 128394 472102
rect 128450 472046 128518 472102
rect 128574 472046 128642 472102
rect 128698 472046 128766 472102
rect 128822 472046 128918 472102
rect 128298 471978 128918 472046
rect 128298 471922 128394 471978
rect 128450 471922 128518 471978
rect 128574 471922 128642 471978
rect 128698 471922 128766 471978
rect 128822 471922 128918 471978
rect 128298 454350 128918 471922
rect 130172 480452 130228 480462
rect 130172 457716 130228 480396
rect 130172 457650 130228 457660
rect 132018 478350 132638 495922
rect 159018 508350 159638 525922
rect 159018 508294 159114 508350
rect 159170 508294 159238 508350
rect 159294 508294 159362 508350
rect 159418 508294 159486 508350
rect 159542 508294 159638 508350
rect 159018 508226 159638 508294
rect 159018 508170 159114 508226
rect 159170 508170 159238 508226
rect 159294 508170 159362 508226
rect 159418 508170 159486 508226
rect 159542 508170 159638 508226
rect 159018 508102 159638 508170
rect 159018 508046 159114 508102
rect 159170 508046 159238 508102
rect 159294 508046 159362 508102
rect 159418 508046 159486 508102
rect 159542 508046 159638 508102
rect 159018 507978 159638 508046
rect 159018 507922 159114 507978
rect 159170 507922 159238 507978
rect 159294 507922 159362 507978
rect 159418 507922 159486 507978
rect 159542 507922 159638 507978
rect 143612 493444 143668 493454
rect 140924 492772 140980 492782
rect 136892 482132 136948 482142
rect 132018 478294 132114 478350
rect 132170 478294 132238 478350
rect 132294 478294 132362 478350
rect 132418 478294 132486 478350
rect 132542 478294 132638 478350
rect 132018 478226 132638 478294
rect 132018 478170 132114 478226
rect 132170 478170 132238 478226
rect 132294 478170 132362 478226
rect 132418 478170 132486 478226
rect 132542 478170 132638 478226
rect 132018 478102 132638 478170
rect 132018 478046 132114 478102
rect 132170 478046 132238 478102
rect 132294 478046 132362 478102
rect 132418 478046 132486 478102
rect 132542 478046 132638 478102
rect 132018 477978 132638 478046
rect 132018 477922 132114 477978
rect 132170 477922 132238 477978
rect 132294 477922 132362 477978
rect 132418 477922 132486 477978
rect 132542 477922 132638 477978
rect 132018 460350 132638 477922
rect 132018 460294 132114 460350
rect 132170 460294 132238 460350
rect 132294 460294 132362 460350
rect 132418 460294 132486 460350
rect 132542 460294 132638 460350
rect 132018 460226 132638 460294
rect 132018 460170 132114 460226
rect 132170 460170 132238 460226
rect 132294 460170 132362 460226
rect 132418 460170 132486 460226
rect 132542 460170 132638 460226
rect 132018 460102 132638 460170
rect 132018 460046 132114 460102
rect 132170 460046 132238 460102
rect 132294 460046 132362 460102
rect 132418 460046 132486 460102
rect 132542 460046 132638 460102
rect 132018 459978 132638 460046
rect 132018 459922 132114 459978
rect 132170 459922 132238 459978
rect 132294 459922 132362 459978
rect 132418 459922 132486 459978
rect 132542 459922 132638 459978
rect 128298 454294 128394 454350
rect 128450 454294 128518 454350
rect 128574 454294 128642 454350
rect 128698 454294 128766 454350
rect 128822 454294 128918 454350
rect 128298 454226 128918 454294
rect 128298 454170 128394 454226
rect 128450 454170 128518 454226
rect 128574 454170 128642 454226
rect 128698 454170 128766 454226
rect 128822 454170 128918 454226
rect 128298 454102 128918 454170
rect 128298 454046 128394 454102
rect 128450 454046 128518 454102
rect 128574 454046 128642 454102
rect 128698 454046 128766 454102
rect 128822 454046 128918 454102
rect 128298 453978 128918 454046
rect 128298 453922 128394 453978
rect 128450 453922 128518 453978
rect 128574 453922 128642 453978
rect 128698 453922 128766 453978
rect 128822 453922 128918 453978
rect 126812 437938 126868 437948
rect 97578 436294 97674 436350
rect 97730 436294 97798 436350
rect 97854 436294 97922 436350
rect 97978 436294 98046 436350
rect 98102 436294 98198 436350
rect 97578 436226 98198 436294
rect 97578 436170 97674 436226
rect 97730 436170 97798 436226
rect 97854 436170 97922 436226
rect 97978 436170 98046 436226
rect 98102 436170 98198 436226
rect 97578 436102 98198 436170
rect 97578 436046 97674 436102
rect 97730 436046 97798 436102
rect 97854 436046 97922 436102
rect 97978 436046 98046 436102
rect 98102 436046 98198 436102
rect 97578 435978 98198 436046
rect 97578 435922 97674 435978
rect 97730 435922 97798 435978
rect 97854 435922 97922 435978
rect 97978 435922 98046 435978
rect 98102 435922 98198 435978
rect 70578 424294 70674 424350
rect 70730 424294 70798 424350
rect 70854 424294 70922 424350
rect 70978 424294 71046 424350
rect 71102 424294 71198 424350
rect 70578 424226 71198 424294
rect 70578 424170 70674 424226
rect 70730 424170 70798 424226
rect 70854 424170 70922 424226
rect 70978 424170 71046 424226
rect 71102 424170 71198 424226
rect 70578 424102 71198 424170
rect 70578 424046 70674 424102
rect 70730 424046 70798 424102
rect 70854 424046 70922 424102
rect 70978 424046 71046 424102
rect 71102 424046 71198 424102
rect 70578 423978 71198 424046
rect 70578 423922 70674 423978
rect 70730 423922 70798 423978
rect 70854 423922 70922 423978
rect 70978 423922 71046 423978
rect 71102 423922 71198 423978
rect 66858 400294 66954 400350
rect 67010 400294 67078 400350
rect 67134 400294 67202 400350
rect 67258 400294 67326 400350
rect 67382 400294 67478 400350
rect 66858 400226 67478 400294
rect 66858 400170 66954 400226
rect 67010 400170 67078 400226
rect 67134 400170 67202 400226
rect 67258 400170 67326 400226
rect 67382 400170 67478 400226
rect 66858 400102 67478 400170
rect 66858 400046 66954 400102
rect 67010 400046 67078 400102
rect 67134 400046 67202 400102
rect 67258 400046 67326 400102
rect 67382 400046 67478 400102
rect 66858 399978 67478 400046
rect 66858 399922 66954 399978
rect 67010 399922 67078 399978
rect 67134 399922 67202 399978
rect 67258 399922 67326 399978
rect 67382 399922 67478 399978
rect 66858 382350 67478 399922
rect 66858 382294 66954 382350
rect 67010 382294 67078 382350
rect 67134 382294 67202 382350
rect 67258 382294 67326 382350
rect 67382 382294 67478 382350
rect 66858 382226 67478 382294
rect 66858 382170 66954 382226
rect 67010 382170 67078 382226
rect 67134 382170 67202 382226
rect 67258 382170 67326 382226
rect 67382 382170 67478 382226
rect 66858 382102 67478 382170
rect 66858 382046 66954 382102
rect 67010 382046 67078 382102
rect 67134 382046 67202 382102
rect 67258 382046 67326 382102
rect 67382 382046 67478 382102
rect 66858 381978 67478 382046
rect 66858 381922 66954 381978
rect 67010 381922 67078 381978
rect 67134 381922 67202 381978
rect 67258 381922 67326 381978
rect 67382 381922 67478 381978
rect 66858 364350 67478 381922
rect 69692 410788 69748 410798
rect 69692 377188 69748 410732
rect 69692 377122 69748 377132
rect 70578 406350 71198 423922
rect 86448 418350 86768 418384
rect 86448 418294 86518 418350
rect 86574 418294 86642 418350
rect 86698 418294 86768 418350
rect 86448 418226 86768 418294
rect 86448 418170 86518 418226
rect 86574 418170 86642 418226
rect 86698 418170 86768 418226
rect 86448 418102 86768 418170
rect 86448 418046 86518 418102
rect 86574 418046 86642 418102
rect 86698 418046 86768 418102
rect 86448 417978 86768 418046
rect 86448 417922 86518 417978
rect 86574 417922 86642 417978
rect 86698 417922 86768 417978
rect 86448 417888 86768 417922
rect 97578 418350 98198 435922
rect 128298 436350 128918 453922
rect 128298 436294 128394 436350
rect 128450 436294 128518 436350
rect 128574 436294 128642 436350
rect 128698 436294 128766 436350
rect 128822 436294 128918 436350
rect 128298 436226 128918 436294
rect 128298 436170 128394 436226
rect 128450 436170 128518 436226
rect 128574 436170 128642 436226
rect 128698 436170 128766 436226
rect 128822 436170 128918 436226
rect 128298 436102 128918 436170
rect 128298 436046 128394 436102
rect 128450 436046 128518 436102
rect 128574 436046 128642 436102
rect 128698 436046 128766 436102
rect 128822 436046 128918 436102
rect 128298 435978 128918 436046
rect 128298 435922 128394 435978
rect 128450 435922 128518 435978
rect 128574 435922 128642 435978
rect 128698 435922 128766 435978
rect 128822 435922 128918 435978
rect 97578 418294 97674 418350
rect 97730 418294 97798 418350
rect 97854 418294 97922 418350
rect 97978 418294 98046 418350
rect 98102 418294 98198 418350
rect 97578 418226 98198 418294
rect 97578 418170 97674 418226
rect 97730 418170 97798 418226
rect 97854 418170 97922 418226
rect 97978 418170 98046 418226
rect 98102 418170 98198 418226
rect 97578 418102 98198 418170
rect 97578 418046 97674 418102
rect 97730 418046 97798 418102
rect 97854 418046 97922 418102
rect 97978 418046 98046 418102
rect 98102 418046 98198 418102
rect 97578 417978 98198 418046
rect 97578 417922 97674 417978
rect 97730 417922 97798 417978
rect 97854 417922 97922 417978
rect 97978 417922 98046 417978
rect 98102 417922 98198 417978
rect 82684 412804 82740 412814
rect 82684 412498 82740 412748
rect 82684 412432 82740 412442
rect 70578 406294 70674 406350
rect 70730 406294 70798 406350
rect 70854 406294 70922 406350
rect 70978 406294 71046 406350
rect 71102 406294 71198 406350
rect 70578 406226 71198 406294
rect 70578 406170 70674 406226
rect 70730 406170 70798 406226
rect 70854 406170 70922 406226
rect 70978 406170 71046 406226
rect 71102 406170 71198 406226
rect 70578 406102 71198 406170
rect 70578 406046 70674 406102
rect 70730 406046 70798 406102
rect 70854 406046 70922 406102
rect 70978 406046 71046 406102
rect 71102 406046 71198 406102
rect 70578 405978 71198 406046
rect 70578 405922 70674 405978
rect 70730 405922 70798 405978
rect 70854 405922 70922 405978
rect 70978 405922 71046 405978
rect 71102 405922 71198 405978
rect 70578 388350 71198 405922
rect 74732 410116 74788 410126
rect 70578 388294 70674 388350
rect 70730 388294 70798 388350
rect 70854 388294 70922 388350
rect 70978 388294 71046 388350
rect 71102 388294 71198 388350
rect 70578 388226 71198 388294
rect 70578 388170 70674 388226
rect 70730 388170 70798 388226
rect 70854 388170 70922 388226
rect 70978 388170 71046 388226
rect 71102 388170 71198 388226
rect 70578 388102 71198 388170
rect 70578 388046 70674 388102
rect 70730 388046 70798 388102
rect 70854 388046 70922 388102
rect 70978 388046 71046 388102
rect 71102 388046 71198 388102
rect 70578 387978 71198 388046
rect 70578 387922 70674 387978
rect 70730 387922 70798 387978
rect 70854 387922 70922 387978
rect 70978 387922 71046 387978
rect 71102 387922 71198 387978
rect 66858 364294 66954 364350
rect 67010 364294 67078 364350
rect 67134 364294 67202 364350
rect 67258 364294 67326 364350
rect 67382 364294 67478 364350
rect 66858 364226 67478 364294
rect 66858 364170 66954 364226
rect 67010 364170 67078 364226
rect 67134 364170 67202 364226
rect 67258 364170 67326 364226
rect 67382 364170 67478 364226
rect 66858 364102 67478 364170
rect 66858 364046 66954 364102
rect 67010 364046 67078 364102
rect 67134 364046 67202 364102
rect 67258 364046 67326 364102
rect 67382 364046 67478 364102
rect 66858 363978 67478 364046
rect 66858 363922 66954 363978
rect 67010 363922 67078 363978
rect 67134 363922 67202 363978
rect 67258 363922 67326 363978
rect 67382 363922 67478 363978
rect 64652 359650 64708 359660
rect 39808 352350 40128 352384
rect 39808 352294 39878 352350
rect 39934 352294 40002 352350
rect 40058 352294 40128 352350
rect 39808 352226 40128 352294
rect 39808 352170 39878 352226
rect 39934 352170 40002 352226
rect 40058 352170 40128 352226
rect 39808 352102 40128 352170
rect 39808 352046 39878 352102
rect 39934 352046 40002 352102
rect 40058 352046 40128 352102
rect 39808 351978 40128 352046
rect 39808 351922 39878 351978
rect 39934 351922 40002 351978
rect 40058 351922 40128 351978
rect 39808 351888 40128 351922
rect 36138 346294 36234 346350
rect 36290 346294 36358 346350
rect 36414 346294 36482 346350
rect 36538 346294 36606 346350
rect 36662 346294 36758 346350
rect 36138 346226 36758 346294
rect 36138 346170 36234 346226
rect 36290 346170 36358 346226
rect 36414 346170 36482 346226
rect 36538 346170 36606 346226
rect 36662 346170 36758 346226
rect 36138 346102 36758 346170
rect 36138 346046 36234 346102
rect 36290 346046 36358 346102
rect 36414 346046 36482 346102
rect 36538 346046 36606 346102
rect 36662 346046 36758 346102
rect 36138 345978 36758 346046
rect 36138 345922 36234 345978
rect 36290 345922 36358 345978
rect 36414 345922 36482 345978
rect 36538 345922 36606 345978
rect 36662 345922 36758 345978
rect 20076 341758 20132 341768
rect 20076 341684 20132 341702
rect 20076 341618 20132 341628
rect 9138 334294 9234 334350
rect 9290 334294 9358 334350
rect 9414 334294 9482 334350
rect 9538 334294 9606 334350
rect 9662 334294 9758 334350
rect 9138 334226 9758 334294
rect 9138 334170 9234 334226
rect 9290 334170 9358 334226
rect 9414 334170 9482 334226
rect 9538 334170 9606 334226
rect 9662 334170 9758 334226
rect 9138 334102 9758 334170
rect 9138 334046 9234 334102
rect 9290 334046 9358 334102
rect 9414 334046 9482 334102
rect 9538 334046 9606 334102
rect 9662 334046 9758 334102
rect 9138 333978 9758 334046
rect 9138 333922 9234 333978
rect 9290 333922 9358 333978
rect 9414 333922 9482 333978
rect 9538 333922 9606 333978
rect 9662 333922 9758 333978
rect 9138 316350 9758 333922
rect 18060 338996 18116 339006
rect 18060 331858 18116 338940
rect 20636 336420 20692 336430
rect 18284 336308 18340 336318
rect 18060 331792 18116 331802
rect 18172 332276 18228 332286
rect 9138 316294 9234 316350
rect 9290 316294 9358 316350
rect 9414 316294 9482 316350
rect 9538 316294 9606 316350
rect 9662 316294 9758 316350
rect 9138 316226 9758 316294
rect 9138 316170 9234 316226
rect 9290 316170 9358 316226
rect 9414 316170 9482 316226
rect 9538 316170 9606 316226
rect 9662 316170 9758 316226
rect 9138 316102 9758 316170
rect 9138 316046 9234 316102
rect 9290 316046 9358 316102
rect 9414 316046 9482 316102
rect 9538 316046 9606 316102
rect 9662 316046 9758 316102
rect 9138 315978 9758 316046
rect 9138 315922 9234 315978
rect 9290 315922 9358 315978
rect 9414 315922 9482 315978
rect 9538 315922 9606 315978
rect 9662 315922 9758 315978
rect 9138 298350 9758 315922
rect 18172 299796 18228 332220
rect 18284 302036 18340 336252
rect 20636 336178 20692 336364
rect 20636 336112 20692 336122
rect 18284 301970 18340 301980
rect 18396 334964 18452 334974
rect 18172 299730 18228 299740
rect 18396 299236 18452 334908
rect 20076 332948 20132 332958
rect 20076 327538 20132 332892
rect 24448 328350 24768 328384
rect 24448 328294 24518 328350
rect 24574 328294 24642 328350
rect 24698 328294 24768 328350
rect 24448 328226 24768 328294
rect 24448 328170 24518 328226
rect 24574 328170 24642 328226
rect 24698 328170 24768 328226
rect 24448 328102 24768 328170
rect 24448 328046 24518 328102
rect 24574 328046 24642 328102
rect 24698 328046 24768 328102
rect 24448 327978 24768 328046
rect 24448 327922 24518 327978
rect 24574 327922 24642 327978
rect 24698 327922 24768 327978
rect 24448 327888 24768 327922
rect 36138 328350 36758 345922
rect 55168 346350 55488 346384
rect 55168 346294 55238 346350
rect 55294 346294 55362 346350
rect 55418 346294 55488 346350
rect 55168 346226 55488 346294
rect 55168 346170 55238 346226
rect 55294 346170 55362 346226
rect 55418 346170 55488 346226
rect 55168 346102 55488 346170
rect 55168 346046 55238 346102
rect 55294 346046 55362 346102
rect 55418 346046 55488 346102
rect 55168 345978 55488 346046
rect 55168 345922 55238 345978
rect 55294 345922 55362 345978
rect 55418 345922 55488 345978
rect 55168 345888 55488 345922
rect 66858 346350 67478 363922
rect 66858 346294 66954 346350
rect 67010 346294 67078 346350
rect 67134 346294 67202 346350
rect 67258 346294 67326 346350
rect 67382 346294 67478 346350
rect 66858 346226 67478 346294
rect 66858 346170 66954 346226
rect 67010 346170 67078 346226
rect 67134 346170 67202 346226
rect 67258 346170 67326 346226
rect 67382 346170 67478 346226
rect 66858 346102 67478 346170
rect 66858 346046 66954 346102
rect 67010 346046 67078 346102
rect 67134 346046 67202 346102
rect 67258 346046 67326 346102
rect 67382 346046 67478 346102
rect 66858 345978 67478 346046
rect 66858 345922 66954 345978
rect 67010 345922 67078 345978
rect 67134 345922 67202 345978
rect 67258 345922 67326 345978
rect 67382 345922 67478 345978
rect 65212 339668 65268 339678
rect 64204 337618 64260 337628
rect 64092 336980 64148 336990
rect 39808 334350 40128 334384
rect 39808 334294 39878 334350
rect 39934 334294 40002 334350
rect 40058 334294 40128 334350
rect 39808 334226 40128 334294
rect 39808 334170 39878 334226
rect 39934 334170 40002 334226
rect 40058 334170 40128 334226
rect 39808 334102 40128 334170
rect 39808 334046 39878 334102
rect 39934 334046 40002 334102
rect 40058 334046 40128 334102
rect 39808 333978 40128 334046
rect 39808 333922 39878 333978
rect 39934 333922 40002 333978
rect 40058 333922 40128 333978
rect 39808 333888 40128 333922
rect 64092 330418 64148 336924
rect 64204 336308 64260 337562
rect 64204 336242 64260 336252
rect 64764 335636 64820 335646
rect 64652 332948 64708 332958
rect 64204 331604 64260 331614
rect 64204 331498 64260 331548
rect 64204 331432 64260 331442
rect 64204 330418 64260 330428
rect 64092 330362 64204 330418
rect 64204 330352 64260 330362
rect 36138 328294 36234 328350
rect 36290 328294 36358 328350
rect 36414 328294 36482 328350
rect 36538 328294 36606 328350
rect 36662 328294 36758 328350
rect 36138 328226 36758 328294
rect 36138 328170 36234 328226
rect 36290 328170 36358 328226
rect 36414 328170 36482 328226
rect 36538 328170 36606 328226
rect 36662 328170 36758 328226
rect 36138 328102 36758 328170
rect 36138 328046 36234 328102
rect 36290 328046 36358 328102
rect 36414 328046 36482 328102
rect 36538 328046 36606 328102
rect 36662 328046 36758 328102
rect 36138 327978 36758 328046
rect 36138 327922 36234 327978
rect 36290 327922 36358 327978
rect 36414 327922 36482 327978
rect 36538 327922 36606 327978
rect 36662 327922 36758 327978
rect 20076 327472 20132 327482
rect 18396 299170 18452 299180
rect 36138 310350 36758 327922
rect 55168 328350 55488 328384
rect 55168 328294 55238 328350
rect 55294 328294 55362 328350
rect 55418 328294 55488 328350
rect 55168 328226 55488 328294
rect 55168 328170 55238 328226
rect 55294 328170 55362 328226
rect 55418 328170 55488 328226
rect 55168 328102 55488 328170
rect 55168 328046 55238 328102
rect 55294 328046 55362 328102
rect 55418 328046 55488 328102
rect 55168 327978 55488 328046
rect 55168 327922 55238 327978
rect 55294 327922 55362 327978
rect 55418 327922 55488 327978
rect 55168 327888 55488 327922
rect 36138 310294 36234 310350
rect 36290 310294 36358 310350
rect 36414 310294 36482 310350
rect 36538 310294 36606 310350
rect 36662 310294 36758 310350
rect 36138 310226 36758 310294
rect 36138 310170 36234 310226
rect 36290 310170 36358 310226
rect 36414 310170 36482 310226
rect 36538 310170 36606 310226
rect 36662 310170 36758 310226
rect 36138 310102 36758 310170
rect 36138 310046 36234 310102
rect 36290 310046 36358 310102
rect 36414 310046 36482 310102
rect 36538 310046 36606 310102
rect 36662 310046 36758 310102
rect 36138 309978 36758 310046
rect 36138 309922 36234 309978
rect 36290 309922 36358 309978
rect 36414 309922 36482 309978
rect 36538 309922 36606 309978
rect 36662 309922 36758 309978
rect 9138 298294 9234 298350
rect 9290 298294 9358 298350
rect 9414 298294 9482 298350
rect 9538 298294 9606 298350
rect 9662 298294 9758 298350
rect 9138 298226 9758 298294
rect 9138 298170 9234 298226
rect 9290 298170 9358 298226
rect 9414 298170 9482 298226
rect 9538 298170 9606 298226
rect 9662 298170 9758 298226
rect 9138 298102 9758 298170
rect 9138 298046 9234 298102
rect 9290 298046 9358 298102
rect 9414 298046 9482 298102
rect 9538 298046 9606 298102
rect 9662 298046 9758 298102
rect 9138 297978 9758 298046
rect 9138 297922 9234 297978
rect 9290 297922 9358 297978
rect 9414 297922 9482 297978
rect 9538 297922 9606 297978
rect 9662 297922 9758 297978
rect 9138 280350 9758 297922
rect 9138 280294 9234 280350
rect 9290 280294 9358 280350
rect 9414 280294 9482 280350
rect 9538 280294 9606 280350
rect 9662 280294 9758 280350
rect 9138 280226 9758 280294
rect 9138 280170 9234 280226
rect 9290 280170 9358 280226
rect 9414 280170 9482 280226
rect 9538 280170 9606 280226
rect 9662 280170 9758 280226
rect 9138 280102 9758 280170
rect 9138 280046 9234 280102
rect 9290 280046 9358 280102
rect 9414 280046 9482 280102
rect 9538 280046 9606 280102
rect 9662 280046 9758 280102
rect 9138 279978 9758 280046
rect 9138 279922 9234 279978
rect 9290 279922 9358 279978
rect 9414 279922 9482 279978
rect 9538 279922 9606 279978
rect 9662 279922 9758 279978
rect 9138 262350 9758 279922
rect 36138 292350 36758 309922
rect 64652 303716 64708 332892
rect 64764 304836 64820 335580
rect 65212 330958 65268 339612
rect 65212 330892 65268 330902
rect 64764 304770 64820 304780
rect 66858 328350 67478 345922
rect 70578 370350 71198 387922
rect 73052 405412 73108 405422
rect 73052 387156 73108 405356
rect 74732 387716 74788 410060
rect 82684 410116 82740 410126
rect 79772 409444 79828 409454
rect 76412 407428 76468 407438
rect 74732 387650 74788 387660
rect 74844 395332 74900 395342
rect 73052 387090 73108 387100
rect 74844 384356 74900 395276
rect 74844 384290 74900 384300
rect 76412 372148 76468 407372
rect 79772 379092 79828 409388
rect 82684 409078 82740 410060
rect 82684 409012 82740 409022
rect 82348 407316 82404 407326
rect 81452 406756 81508 406766
rect 81452 385476 81508 406700
rect 82348 406738 82404 407260
rect 97578 406894 98198 417922
rect 117168 418350 117488 418384
rect 117168 418294 117238 418350
rect 117294 418294 117362 418350
rect 117418 418294 117488 418350
rect 117168 418226 117488 418294
rect 117168 418170 117238 418226
rect 117294 418170 117362 418226
rect 117418 418170 117488 418226
rect 117168 418102 117488 418170
rect 117168 418046 117238 418102
rect 117294 418046 117362 418102
rect 117418 418046 117488 418102
rect 117168 417978 117488 418046
rect 117168 417922 117238 417978
rect 117294 417922 117362 417978
rect 117418 417922 117488 417978
rect 117168 417888 117488 417922
rect 128298 418350 128918 435922
rect 128298 418294 128394 418350
rect 128450 418294 128518 418350
rect 128574 418294 128642 418350
rect 128698 418294 128766 418350
rect 128822 418294 128918 418350
rect 128298 418226 128918 418294
rect 128298 418170 128394 418226
rect 128450 418170 128518 418226
rect 128574 418170 128642 418226
rect 128698 418170 128766 418226
rect 128822 418170 128918 418226
rect 128298 418102 128918 418170
rect 128298 418046 128394 418102
rect 128450 418046 128518 418102
rect 128574 418046 128642 418102
rect 128698 418046 128766 418102
rect 128822 418046 128918 418102
rect 128298 417978 128918 418046
rect 128298 417922 128394 417978
rect 128450 417922 128518 417978
rect 128574 417922 128642 417978
rect 128698 417922 128766 417978
rect 128822 417922 128918 417978
rect 127036 410788 127092 410798
rect 126812 410116 126868 410126
rect 126252 409444 126308 409454
rect 82348 406672 82404 406682
rect 125132 406738 125188 406748
rect 101808 406350 102128 406384
rect 101808 406294 101878 406350
rect 101934 406294 102002 406350
rect 102058 406294 102128 406350
rect 101808 406226 102128 406294
rect 101808 406170 101878 406226
rect 101934 406170 102002 406226
rect 102058 406170 102128 406226
rect 101808 406102 102128 406170
rect 101808 406046 101878 406102
rect 101934 406046 102002 406102
rect 102058 406046 102128 406102
rect 101808 405978 102128 406046
rect 101808 405922 101878 405978
rect 101934 405922 102002 405978
rect 102058 405922 102128 405978
rect 101808 405888 102128 405922
rect 81564 404740 81620 404750
rect 81564 387940 81620 404684
rect 82348 400708 82404 400718
rect 82348 398098 82404 400652
rect 86448 400350 86768 400384
rect 86448 400294 86518 400350
rect 86574 400294 86642 400350
rect 86698 400294 86768 400350
rect 86448 400226 86768 400294
rect 86448 400170 86518 400226
rect 86574 400170 86642 400226
rect 86698 400170 86768 400226
rect 86448 400102 86768 400170
rect 86448 400046 86518 400102
rect 86574 400046 86642 400102
rect 86698 400046 86768 400102
rect 86448 399978 86768 400046
rect 86448 399922 86518 399978
rect 86574 399922 86642 399978
rect 86698 399922 86768 399978
rect 86448 399888 86768 399922
rect 117168 400350 117488 400384
rect 117168 400294 117238 400350
rect 117294 400294 117362 400350
rect 117418 400294 117488 400350
rect 117168 400226 117488 400294
rect 117168 400170 117238 400226
rect 117294 400170 117362 400226
rect 117418 400170 117488 400226
rect 117168 400102 117488 400170
rect 117168 400046 117238 400102
rect 117294 400046 117362 400102
rect 117418 400046 117488 400102
rect 117168 399978 117488 400046
rect 117168 399922 117238 399978
rect 117294 399922 117362 399978
rect 117418 399922 117488 399978
rect 117168 399888 117488 399922
rect 82348 398032 82404 398042
rect 81564 387874 81620 387884
rect 81452 385410 81508 385420
rect 79772 379026 79828 379036
rect 97578 382350 98198 399122
rect 125132 396478 125188 406682
rect 126252 402418 126308 409388
rect 126252 402352 126308 402362
rect 125132 396412 125188 396422
rect 101808 388389 102128 388446
rect 101808 388333 101836 388389
rect 101892 388333 101940 388389
rect 101996 388333 102044 388389
rect 102100 388333 102128 388389
rect 101808 388276 102128 388333
rect 97578 382294 97674 382350
rect 97730 382294 97798 382350
rect 97854 382294 97922 382350
rect 97978 382294 98046 382350
rect 98102 382294 98198 382350
rect 97578 382226 98198 382294
rect 97578 382170 97674 382226
rect 97730 382170 97798 382226
rect 97854 382170 97922 382226
rect 97978 382170 98046 382226
rect 98102 382170 98198 382226
rect 97578 382102 98198 382170
rect 97578 382046 97674 382102
rect 97730 382046 97798 382102
rect 97854 382046 97922 382102
rect 97978 382046 98046 382102
rect 98102 382046 98198 382102
rect 97578 381978 98198 382046
rect 97578 381922 97674 381978
rect 97730 381922 97798 381978
rect 97854 381922 97922 381978
rect 97978 381922 98046 381978
rect 98102 381922 98198 381978
rect 76412 372082 76468 372092
rect 70578 370294 70674 370350
rect 70730 370294 70798 370350
rect 70854 370294 70922 370350
rect 70978 370294 71046 370350
rect 71102 370294 71198 370350
rect 70578 370226 71198 370294
rect 70578 370170 70674 370226
rect 70730 370170 70798 370226
rect 70854 370170 70922 370226
rect 70978 370170 71046 370226
rect 71102 370170 71198 370226
rect 70578 370102 71198 370170
rect 70578 370046 70674 370102
rect 70730 370046 70798 370102
rect 70854 370046 70922 370102
rect 70978 370046 71046 370102
rect 71102 370046 71198 370102
rect 70578 369978 71198 370046
rect 70578 369922 70674 369978
rect 70730 369922 70798 369978
rect 70854 369922 70922 369978
rect 70978 369922 71046 369978
rect 71102 369922 71198 369978
rect 70578 352350 71198 369922
rect 70578 352294 70674 352350
rect 70730 352294 70798 352350
rect 70854 352294 70922 352350
rect 70978 352294 71046 352350
rect 71102 352294 71198 352350
rect 70578 352226 71198 352294
rect 70578 352170 70674 352226
rect 70730 352170 70798 352226
rect 70854 352170 70922 352226
rect 70978 352170 71046 352226
rect 71102 352170 71198 352226
rect 70578 352102 71198 352170
rect 70578 352046 70674 352102
rect 70730 352046 70798 352102
rect 70854 352046 70922 352102
rect 70978 352046 71046 352102
rect 71102 352046 71198 352102
rect 70578 351978 71198 352046
rect 70578 351922 70674 351978
rect 70730 351922 70798 351978
rect 70854 351922 70922 351978
rect 70978 351922 71046 351978
rect 71102 351922 71198 351978
rect 70578 334350 71198 351922
rect 97578 364350 98198 381922
rect 126812 365316 126868 410060
rect 126924 404068 126980 404078
rect 126924 366436 126980 404012
rect 127036 369236 127092 410732
rect 127260 408772 127316 408782
rect 127036 369170 127092 369180
rect 127148 406084 127204 406094
rect 126924 366370 126980 366380
rect 126812 365250 126868 365260
rect 127148 364756 127204 406028
rect 127260 368116 127316 408716
rect 127260 368050 127316 368060
rect 128298 400350 128918 417922
rect 128298 400294 128394 400350
rect 128450 400294 128518 400350
rect 128574 400294 128642 400350
rect 128698 400294 128766 400350
rect 128822 400294 128918 400350
rect 128298 400226 128918 400294
rect 128298 400170 128394 400226
rect 128450 400170 128518 400226
rect 128574 400170 128642 400226
rect 128698 400170 128766 400226
rect 128822 400170 128918 400226
rect 128298 400102 128918 400170
rect 128298 400046 128394 400102
rect 128450 400046 128518 400102
rect 128574 400046 128642 400102
rect 128698 400046 128766 400102
rect 128822 400046 128918 400102
rect 128298 399978 128918 400046
rect 128298 399922 128394 399978
rect 128450 399922 128518 399978
rect 128574 399922 128642 399978
rect 128698 399922 128766 399978
rect 128822 399922 128918 399978
rect 128298 382350 128918 399922
rect 128298 382294 128394 382350
rect 128450 382294 128518 382350
rect 128574 382294 128642 382350
rect 128698 382294 128766 382350
rect 128822 382294 128918 382350
rect 128298 382226 128918 382294
rect 128298 382170 128394 382226
rect 128450 382170 128518 382226
rect 128574 382170 128642 382226
rect 128698 382170 128766 382226
rect 128822 382170 128918 382226
rect 128298 382102 128918 382170
rect 128298 382046 128394 382102
rect 128450 382046 128518 382102
rect 128574 382046 128642 382102
rect 128698 382046 128766 382102
rect 128822 382046 128918 382102
rect 128298 381978 128918 382046
rect 128298 381922 128394 381978
rect 128450 381922 128518 381978
rect 128574 381922 128642 381978
rect 128698 381922 128766 381978
rect 128822 381922 128918 381978
rect 127148 364690 127204 364700
rect 97578 364294 97674 364350
rect 97730 364294 97798 364350
rect 97854 364294 97922 364350
rect 97978 364294 98046 364350
rect 98102 364294 98198 364350
rect 97578 364226 98198 364294
rect 97578 364170 97674 364226
rect 97730 364170 97798 364226
rect 97854 364170 97922 364226
rect 97978 364170 98046 364226
rect 98102 364170 98198 364226
rect 97578 364102 98198 364170
rect 97578 364046 97674 364102
rect 97730 364046 97798 364102
rect 97854 364046 97922 364102
rect 97978 364046 98046 364102
rect 98102 364046 98198 364102
rect 97578 363978 98198 364046
rect 97578 363922 97674 363978
rect 97730 363922 97798 363978
rect 97854 363922 97922 363978
rect 97978 363922 98046 363978
rect 98102 363922 98198 363978
rect 86448 346350 86768 346384
rect 86448 346294 86518 346350
rect 86574 346294 86642 346350
rect 86698 346294 86768 346350
rect 86448 346226 86768 346294
rect 86448 346170 86518 346226
rect 86574 346170 86642 346226
rect 86698 346170 86768 346226
rect 86448 346102 86768 346170
rect 86448 346046 86518 346102
rect 86574 346046 86642 346102
rect 86698 346046 86768 346102
rect 86448 345978 86768 346046
rect 86448 345922 86518 345978
rect 86574 345922 86642 345978
rect 86698 345922 86768 345978
rect 86448 345888 86768 345922
rect 97578 346350 98198 363922
rect 128298 364350 128918 381922
rect 128298 364294 128394 364350
rect 128450 364294 128518 364350
rect 128574 364294 128642 364350
rect 128698 364294 128766 364350
rect 128822 364294 128918 364350
rect 128298 364226 128918 364294
rect 128298 364170 128394 364226
rect 128450 364170 128518 364226
rect 128574 364170 128642 364226
rect 128698 364170 128766 364226
rect 128822 364170 128918 364226
rect 128298 364102 128918 364170
rect 128298 364046 128394 364102
rect 128450 364046 128518 364102
rect 128574 364046 128642 364102
rect 128698 364046 128766 364102
rect 128822 364046 128918 364102
rect 128298 363978 128918 364046
rect 128298 363922 128394 363978
rect 128450 363922 128518 363978
rect 128574 363922 128642 363978
rect 128698 363922 128766 363978
rect 128822 363922 128918 363978
rect 101808 352350 102128 352384
rect 101808 352294 101878 352350
rect 101934 352294 102002 352350
rect 102058 352294 102128 352350
rect 101808 352226 102128 352294
rect 101808 352170 101878 352226
rect 101934 352170 102002 352226
rect 102058 352170 102128 352226
rect 101808 352102 102128 352170
rect 101808 352046 101878 352102
rect 101934 352046 102002 352102
rect 102058 352046 102128 352102
rect 101808 351978 102128 352046
rect 101808 351922 101878 351978
rect 101934 351922 102002 351978
rect 102058 351922 102128 351978
rect 101808 351888 102128 351922
rect 97578 346294 97674 346350
rect 97730 346294 97798 346350
rect 97854 346294 97922 346350
rect 97978 346294 98046 346350
rect 98102 346294 98198 346350
rect 97578 346226 98198 346294
rect 97578 346170 97674 346226
rect 97730 346170 97798 346226
rect 97854 346170 97922 346226
rect 97978 346170 98046 346226
rect 98102 346170 98198 346226
rect 97578 346102 98198 346170
rect 97578 346046 97674 346102
rect 97730 346046 97798 346102
rect 97854 346046 97922 346102
rect 97978 346046 98046 346102
rect 98102 346046 98198 346102
rect 97578 345978 98198 346046
rect 97578 345922 97674 345978
rect 97730 345922 97798 345978
rect 97854 345922 97922 345978
rect 97978 345922 98046 345978
rect 98102 345922 98198 345978
rect 82684 341938 82740 341948
rect 82684 341684 82740 341882
rect 82684 341618 82740 341628
rect 82460 340340 82516 340356
rect 82460 340252 82516 340262
rect 82236 338518 82292 338528
rect 82236 337652 82292 338462
rect 82236 337586 82292 337596
rect 70578 334294 70674 334350
rect 70730 334294 70798 334350
rect 70854 334294 70922 334350
rect 70978 334294 71046 334350
rect 71102 334294 71198 334350
rect 70578 334226 71198 334294
rect 70578 334170 70674 334226
rect 70730 334170 70798 334226
rect 70854 334170 70922 334226
rect 70978 334170 71046 334226
rect 71102 334170 71198 334226
rect 70578 334102 71198 334170
rect 70578 334046 70674 334102
rect 70730 334046 70798 334102
rect 70854 334046 70922 334102
rect 70978 334046 71046 334102
rect 71102 334046 71198 334102
rect 70578 333978 71198 334046
rect 70578 333922 70674 333978
rect 70730 333922 70798 333978
rect 70854 333922 70922 333978
rect 70978 333922 71046 333978
rect 71102 333922 71198 333978
rect 66858 328294 66954 328350
rect 67010 328294 67078 328350
rect 67134 328294 67202 328350
rect 67258 328294 67326 328350
rect 67382 328294 67478 328350
rect 66858 328226 67478 328294
rect 66858 328170 66954 328226
rect 67010 328170 67078 328226
rect 67134 328170 67202 328226
rect 67258 328170 67326 328226
rect 67382 328170 67478 328226
rect 66858 328102 67478 328170
rect 66858 328046 66954 328102
rect 67010 328046 67078 328102
rect 67134 328046 67202 328102
rect 67258 328046 67326 328102
rect 67382 328046 67478 328102
rect 66858 327978 67478 328046
rect 66858 327922 66954 327978
rect 67010 327922 67078 327978
rect 67134 327922 67202 327978
rect 67258 327922 67326 327978
rect 67382 327922 67478 327978
rect 66858 310350 67478 327922
rect 66858 310294 66954 310350
rect 67010 310294 67078 310350
rect 67134 310294 67202 310350
rect 67258 310294 67326 310350
rect 67382 310294 67478 310350
rect 66858 310226 67478 310294
rect 66858 310170 66954 310226
rect 67010 310170 67078 310226
rect 67134 310170 67202 310226
rect 67258 310170 67326 310226
rect 67382 310170 67478 310226
rect 66858 310102 67478 310170
rect 66858 310046 66954 310102
rect 67010 310046 67078 310102
rect 67134 310046 67202 310102
rect 67258 310046 67326 310102
rect 67382 310046 67478 310102
rect 66858 309978 67478 310046
rect 66858 309922 66954 309978
rect 67010 309922 67078 309978
rect 67134 309922 67202 309978
rect 67258 309922 67326 309978
rect 67382 309922 67478 309978
rect 64652 303650 64708 303660
rect 36138 292294 36234 292350
rect 36290 292294 36358 292350
rect 36414 292294 36482 292350
rect 36538 292294 36606 292350
rect 36662 292294 36758 292350
rect 36138 292226 36758 292294
rect 36138 292170 36234 292226
rect 36290 292170 36358 292226
rect 36414 292170 36482 292226
rect 36538 292170 36606 292226
rect 36662 292170 36758 292226
rect 36138 292102 36758 292170
rect 36138 292046 36234 292102
rect 36290 292046 36358 292102
rect 36414 292046 36482 292102
rect 36538 292046 36606 292102
rect 36662 292046 36758 292102
rect 36138 291978 36758 292046
rect 36138 291922 36234 291978
rect 36290 291922 36358 291978
rect 36414 291922 36482 291978
rect 36538 291922 36606 291978
rect 36662 291922 36758 291978
rect 24448 274350 24768 274384
rect 24448 274294 24518 274350
rect 24574 274294 24642 274350
rect 24698 274294 24768 274350
rect 24448 274226 24768 274294
rect 24448 274170 24518 274226
rect 24574 274170 24642 274226
rect 24698 274170 24768 274226
rect 24448 274102 24768 274170
rect 24448 274046 24518 274102
rect 24574 274046 24642 274102
rect 24698 274046 24768 274102
rect 24448 273978 24768 274046
rect 24448 273922 24518 273978
rect 24574 273922 24642 273978
rect 24698 273922 24768 273978
rect 24448 273888 24768 273922
rect 36138 274350 36758 291922
rect 66858 292350 67478 309922
rect 69692 332276 69748 332286
rect 69692 308308 69748 332220
rect 69692 308242 69748 308252
rect 70578 316350 71198 333922
rect 80556 336420 80612 336430
rect 80556 331492 80612 336364
rect 80556 331426 80612 331436
rect 81452 331492 81508 331502
rect 70578 316294 70674 316350
rect 70730 316294 70798 316350
rect 70854 316294 70922 316350
rect 70978 316294 71046 316350
rect 71102 316294 71198 316350
rect 70578 316226 71198 316294
rect 70578 316170 70674 316226
rect 70730 316170 70798 316226
rect 70854 316170 70922 316226
rect 70978 316170 71046 316226
rect 71102 316170 71198 316226
rect 70578 316102 71198 316170
rect 70578 316046 70674 316102
rect 70730 316046 70798 316102
rect 70854 316046 70922 316102
rect 70978 316046 71046 316102
rect 71102 316046 71198 316102
rect 70578 315978 71198 316046
rect 70578 315922 70674 315978
rect 70730 315922 70798 315978
rect 70854 315922 70922 315978
rect 70978 315922 71046 315978
rect 71102 315922 71198 315978
rect 66858 292294 66954 292350
rect 67010 292294 67078 292350
rect 67134 292294 67202 292350
rect 67258 292294 67326 292350
rect 67382 292294 67478 292350
rect 66858 292226 67478 292294
rect 66858 292170 66954 292226
rect 67010 292170 67078 292226
rect 67134 292170 67202 292226
rect 67258 292170 67326 292226
rect 67382 292170 67478 292226
rect 66858 292102 67478 292170
rect 66858 292046 66954 292102
rect 67010 292046 67078 292102
rect 67134 292046 67202 292102
rect 67258 292046 67326 292102
rect 67382 292046 67478 292102
rect 66858 291978 67478 292046
rect 66858 291922 66954 291978
rect 67010 291922 67078 291978
rect 67134 291922 67202 291978
rect 67258 291922 67326 291978
rect 67382 291922 67478 291978
rect 39808 280350 40128 280384
rect 39808 280294 39878 280350
rect 39934 280294 40002 280350
rect 40058 280294 40128 280350
rect 39808 280226 40128 280294
rect 39808 280170 39878 280226
rect 39934 280170 40002 280226
rect 40058 280170 40128 280226
rect 39808 280102 40128 280170
rect 39808 280046 39878 280102
rect 39934 280046 40002 280102
rect 40058 280046 40128 280102
rect 39808 279978 40128 280046
rect 39808 279922 39878 279978
rect 39934 279922 40002 279978
rect 40058 279922 40128 279978
rect 39808 279888 40128 279922
rect 64204 277172 64260 277182
rect 64204 275698 64260 277116
rect 64204 275632 64260 275642
rect 36138 274294 36234 274350
rect 36290 274294 36358 274350
rect 36414 274294 36482 274350
rect 36538 274294 36606 274350
rect 36662 274294 36758 274350
rect 36138 274226 36758 274294
rect 36138 274170 36234 274226
rect 36290 274170 36358 274226
rect 36414 274170 36482 274226
rect 36538 274170 36606 274226
rect 36662 274170 36758 274226
rect 36138 274102 36758 274170
rect 36138 274046 36234 274102
rect 36290 274046 36358 274102
rect 36414 274046 36482 274102
rect 36538 274046 36606 274102
rect 36662 274046 36758 274102
rect 36138 273978 36758 274046
rect 36138 273922 36234 273978
rect 36290 273922 36358 273978
rect 36414 273922 36482 273978
rect 36538 273922 36606 273978
rect 36662 273922 36758 273978
rect 20076 270478 20132 270490
rect 20076 270386 20132 270396
rect 9138 262294 9234 262350
rect 9290 262294 9358 262350
rect 9414 262294 9482 262350
rect 9538 262294 9606 262350
rect 9662 262294 9758 262350
rect 9138 262226 9758 262294
rect 9138 262170 9234 262226
rect 9290 262170 9358 262226
rect 9414 262170 9482 262226
rect 9538 262170 9606 262226
rect 9662 262170 9758 262226
rect 9138 262102 9758 262170
rect 9138 262046 9234 262102
rect 9290 262046 9358 262102
rect 9414 262046 9482 262102
rect 9538 262046 9606 262102
rect 9662 262046 9758 262102
rect 9138 261978 9758 262046
rect 9138 261922 9234 261978
rect 9290 261922 9358 261978
rect 9414 261922 9482 261978
rect 9538 261922 9606 261978
rect 9662 261922 9758 261978
rect 9138 244350 9758 261922
rect 18396 268436 18452 268446
rect 18396 245364 18452 268380
rect 36138 267966 36758 273922
rect 55168 274350 55488 274384
rect 55168 274294 55238 274350
rect 55294 274294 55362 274350
rect 55418 274294 55488 274350
rect 55168 274226 55488 274294
rect 55168 274170 55238 274226
rect 55294 274170 55362 274226
rect 55418 274170 55488 274226
rect 55168 274102 55488 274170
rect 55168 274046 55238 274102
rect 55294 274046 55362 274102
rect 55418 274046 55488 274102
rect 55168 273978 55488 274046
rect 55168 273922 55238 273978
rect 55294 273922 55362 273978
rect 55418 273922 55488 273978
rect 55168 273888 55488 273922
rect 66858 274350 67478 291922
rect 66858 274294 66954 274350
rect 67010 274294 67078 274350
rect 67134 274294 67202 274350
rect 67258 274294 67326 274350
rect 67382 274294 67478 274350
rect 66858 274226 67478 274294
rect 66858 274170 66954 274226
rect 67010 274170 67078 274226
rect 67134 274170 67202 274226
rect 67258 274170 67326 274226
rect 67382 274170 67478 274226
rect 66858 274102 67478 274170
rect 66858 274046 66954 274102
rect 67010 274046 67078 274102
rect 67134 274046 67202 274102
rect 67258 274046 67326 274102
rect 67382 274046 67478 274102
rect 66858 273978 67478 274046
rect 66858 273922 66954 273978
rect 67010 273922 67078 273978
rect 67134 273922 67202 273978
rect 67258 273922 67326 273978
rect 67382 273922 67478 273978
rect 64652 270838 64708 270848
rect 64204 270298 64260 270308
rect 64092 270242 64204 270298
rect 64092 269108 64148 270242
rect 64204 270232 64260 270242
rect 64204 270118 64260 270128
rect 64204 269780 64260 270062
rect 64204 269714 64260 269724
rect 64092 269042 64148 269052
rect 64204 268678 64260 268688
rect 18396 245298 18452 245308
rect 20076 267764 20132 267774
rect 9138 244294 9234 244350
rect 9290 244294 9358 244350
rect 9414 244294 9482 244350
rect 9538 244294 9606 244350
rect 9662 244294 9758 244350
rect 9138 244226 9758 244294
rect 9138 244170 9234 244226
rect 9290 244170 9358 244226
rect 9414 244170 9482 244226
rect 9538 244170 9606 244226
rect 9662 244170 9758 244226
rect 9138 244102 9758 244170
rect 9138 244046 9234 244102
rect 9290 244046 9358 244102
rect 9414 244046 9482 244102
rect 9538 244046 9606 244102
rect 9662 244046 9758 244102
rect 9138 243978 9758 244046
rect 9138 243922 9234 243978
rect 9290 243922 9358 243978
rect 9414 243922 9482 243978
rect 9538 243922 9606 243978
rect 9662 243922 9758 243978
rect 9138 226350 9758 243922
rect 20076 240996 20132 267708
rect 64204 267764 64260 268622
rect 64204 267698 64260 267708
rect 64652 265748 64708 270782
rect 64652 265682 64708 265692
rect 64204 264538 64260 264548
rect 64204 263732 64260 264482
rect 64204 263666 64260 263676
rect 64204 263060 64260 263070
rect 39808 262350 40128 262384
rect 39808 262294 39878 262350
rect 39934 262294 40002 262350
rect 40058 262294 40128 262350
rect 39808 262226 40128 262294
rect 39808 262170 39878 262226
rect 39934 262170 40002 262226
rect 40058 262170 40128 262226
rect 39808 262102 40128 262170
rect 39808 262046 39878 262102
rect 39934 262046 40002 262102
rect 40058 262046 40128 262102
rect 39808 261978 40128 262046
rect 39808 261922 39878 261978
rect 39934 261922 40002 261978
rect 40058 261922 40128 261978
rect 39808 261888 40128 261922
rect 64204 261268 64260 263004
rect 64204 261202 64260 261212
rect 64764 261716 64820 261726
rect 64652 260372 64708 260382
rect 24448 256350 24768 256384
rect 24448 256294 24518 256350
rect 24574 256294 24642 256350
rect 24698 256294 24768 256350
rect 24448 256226 24768 256294
rect 24448 256170 24518 256226
rect 24574 256170 24642 256226
rect 24698 256170 24768 256226
rect 24448 256102 24768 256170
rect 24448 256046 24518 256102
rect 24574 256046 24642 256102
rect 24698 256046 24768 256102
rect 24448 255978 24768 256046
rect 24448 255922 24518 255978
rect 24574 255922 24642 255978
rect 24698 255922 24768 255978
rect 24448 255888 24768 255922
rect 36138 256350 36758 256610
rect 36138 256294 36234 256350
rect 36290 256294 36358 256350
rect 36414 256294 36482 256350
rect 36538 256294 36606 256350
rect 36662 256294 36758 256350
rect 36138 256226 36758 256294
rect 36138 256170 36234 256226
rect 36290 256170 36358 256226
rect 36414 256170 36482 256226
rect 36538 256170 36606 256226
rect 36662 256170 36758 256226
rect 36138 256102 36758 256170
rect 36138 256046 36234 256102
rect 36290 256046 36358 256102
rect 36414 256046 36482 256102
rect 36538 256046 36606 256102
rect 36662 256046 36758 256102
rect 36138 255978 36758 256046
rect 36138 255922 36234 255978
rect 36290 255922 36358 255978
rect 36414 255922 36482 255978
rect 36538 255922 36606 255978
rect 36662 255922 36758 255978
rect 20972 245364 21028 245374
rect 20972 242116 21028 245308
rect 20972 242050 21028 242060
rect 20076 240930 20132 240940
rect 9138 226294 9234 226350
rect 9290 226294 9358 226350
rect 9414 226294 9482 226350
rect 9538 226294 9606 226350
rect 9662 226294 9758 226350
rect 9138 226226 9758 226294
rect 9138 226170 9234 226226
rect 9290 226170 9358 226226
rect 9414 226170 9482 226226
rect 9538 226170 9606 226226
rect 9662 226170 9758 226226
rect 9138 226102 9758 226170
rect 9138 226046 9234 226102
rect 9290 226046 9358 226102
rect 9414 226046 9482 226102
rect 9538 226046 9606 226102
rect 9662 226046 9758 226102
rect 9138 225978 9758 226046
rect 9138 225922 9234 225978
rect 9290 225922 9358 225978
rect 9414 225922 9482 225978
rect 9538 225922 9606 225978
rect 9662 225922 9758 225978
rect 9138 208350 9758 225922
rect 36138 238350 36758 255922
rect 55168 256350 55488 256384
rect 55168 256294 55238 256350
rect 55294 256294 55362 256350
rect 55418 256294 55488 256350
rect 55168 256226 55488 256294
rect 55168 256170 55238 256226
rect 55294 256170 55362 256226
rect 55418 256170 55488 256226
rect 55168 256102 55488 256170
rect 55168 256046 55238 256102
rect 55294 256046 55362 256102
rect 55418 256046 55488 256102
rect 55168 255978 55488 256046
rect 55168 255922 55238 255978
rect 55294 255922 55362 255978
rect 55418 255922 55488 255978
rect 55168 255888 55488 255922
rect 64652 245252 64708 260316
rect 64764 252868 64820 261660
rect 64764 252802 64820 252812
rect 66858 256350 67478 273922
rect 70578 298350 71198 315922
rect 80444 329700 80500 329710
rect 80444 314692 80500 329644
rect 80444 314626 80500 314636
rect 80556 329364 80612 329374
rect 80556 312116 80612 329308
rect 80556 312050 80612 312060
rect 81452 308196 81508 331436
rect 86448 328350 86768 328384
rect 86448 328294 86518 328350
rect 86574 328294 86642 328350
rect 86698 328294 86768 328350
rect 86448 328226 86768 328294
rect 86448 328170 86518 328226
rect 86574 328170 86642 328226
rect 86698 328170 86768 328226
rect 86448 328102 86768 328170
rect 86448 328046 86518 328102
rect 86574 328046 86642 328102
rect 86698 328046 86768 328102
rect 86448 327978 86768 328046
rect 86448 327922 86518 327978
rect 86574 327922 86642 327978
rect 86698 327922 86768 327978
rect 86448 327888 86768 327922
rect 97578 328350 98198 345922
rect 117168 346350 117488 346384
rect 117168 346294 117238 346350
rect 117294 346294 117362 346350
rect 117418 346294 117488 346350
rect 117168 346226 117488 346294
rect 117168 346170 117238 346226
rect 117294 346170 117362 346226
rect 117418 346170 117488 346226
rect 117168 346102 117488 346170
rect 117168 346046 117238 346102
rect 117294 346046 117362 346102
rect 117418 346046 117488 346102
rect 117168 345978 117488 346046
rect 117168 345922 117238 345978
rect 117294 345922 117362 345978
rect 117418 345922 117488 345978
rect 117168 345888 117488 345922
rect 128298 346350 128918 363922
rect 128298 346294 128394 346350
rect 128450 346294 128518 346350
rect 128574 346294 128642 346350
rect 128698 346294 128766 346350
rect 128822 346294 128918 346350
rect 128298 346226 128918 346294
rect 128298 346170 128394 346226
rect 128450 346170 128518 346226
rect 128574 346170 128642 346226
rect 128698 346170 128766 346226
rect 128822 346170 128918 346226
rect 128298 346102 128918 346170
rect 128298 346046 128394 346102
rect 128450 346046 128518 346102
rect 128574 346046 128642 346102
rect 128698 346046 128766 346102
rect 128822 346046 128918 346102
rect 128298 345978 128918 346046
rect 128298 345922 128394 345978
rect 128450 345922 128518 345978
rect 128574 345922 128642 345978
rect 128698 345922 128766 345978
rect 128822 345922 128918 345978
rect 122668 340498 122724 340508
rect 122668 338518 122724 340442
rect 127484 340340 127540 340350
rect 122668 338452 122724 338462
rect 126140 339332 126196 339342
rect 124348 336178 124404 336188
rect 101808 334350 102128 334384
rect 101808 334294 101878 334350
rect 101934 334294 102002 334350
rect 102058 334294 102128 334350
rect 101808 334226 102128 334294
rect 101808 334170 101878 334226
rect 101934 334170 102002 334226
rect 102058 334170 102128 334226
rect 101808 334102 102128 334170
rect 101808 334046 101878 334102
rect 101934 334046 102002 334102
rect 102058 334046 102128 334102
rect 101808 333978 102128 334046
rect 101808 333922 101878 333978
rect 101934 333922 102002 333978
rect 102058 333922 102128 333978
rect 101808 333888 102128 333922
rect 97578 328294 97674 328350
rect 97730 328294 97798 328350
rect 97854 328294 97922 328350
rect 97978 328294 98046 328350
rect 98102 328294 98198 328350
rect 97578 328226 98198 328294
rect 97578 328170 97674 328226
rect 97730 328170 97798 328226
rect 97854 328170 97922 328226
rect 97978 328170 98046 328226
rect 98102 328170 98198 328226
rect 97578 328102 98198 328170
rect 97578 328046 97674 328102
rect 97730 328046 97798 328102
rect 97854 328046 97922 328102
rect 97978 328046 98046 328102
rect 98102 328046 98198 328102
rect 97578 327978 98198 328046
rect 97578 327922 97674 327978
rect 97730 327922 97798 327978
rect 97854 327922 97922 327978
rect 97978 327922 98046 327978
rect 98102 327922 98198 327978
rect 81452 308130 81508 308140
rect 97578 310350 98198 327922
rect 117168 328350 117488 328384
rect 117168 328294 117238 328350
rect 117294 328294 117362 328350
rect 117418 328294 117488 328350
rect 117168 328226 117488 328294
rect 117168 328170 117238 328226
rect 117294 328170 117362 328226
rect 117418 328170 117488 328226
rect 117168 328102 117488 328170
rect 117168 328046 117238 328102
rect 117294 328046 117362 328102
rect 117418 328046 117488 328102
rect 117168 327978 117488 328046
rect 117168 327922 117238 327978
rect 117294 327922 117362 327978
rect 117418 327922 117488 327978
rect 117168 327888 117488 327922
rect 124348 327358 124404 336122
rect 126140 333620 126196 339276
rect 127484 338548 127540 340284
rect 127484 338482 127540 338492
rect 127596 339238 127652 339248
rect 127596 338324 127652 339182
rect 127596 338258 127652 338268
rect 127596 336980 127652 336990
rect 127596 336178 127652 336924
rect 127596 336112 127652 336122
rect 126140 333554 126196 333564
rect 127596 332948 127652 332958
rect 127596 332758 127652 332892
rect 127596 332692 127652 332702
rect 127596 330778 127652 330788
rect 124348 327292 124404 327302
rect 126812 330260 126868 330270
rect 126812 313348 126868 330204
rect 127596 329588 127652 330722
rect 127596 329522 127652 329532
rect 126812 313282 126868 313292
rect 128298 328350 128918 345922
rect 132018 442350 132638 459922
rect 133532 480004 133588 480014
rect 133532 457044 133588 479948
rect 133532 456978 133588 456988
rect 135212 476644 135268 476654
rect 135212 456036 135268 476588
rect 135212 455970 135268 455980
rect 136892 455476 136948 482076
rect 140924 480452 140980 492716
rect 141036 483812 141092 483822
rect 141036 483058 141092 483756
rect 141036 482992 141092 483002
rect 142044 481348 142100 481358
rect 140924 480386 140980 480396
rect 141036 480676 141092 480686
rect 140924 477316 140980 477326
rect 140812 476644 140868 476654
rect 136892 455410 136948 455420
rect 138572 476308 138628 476318
rect 138572 454356 138628 476252
rect 138572 454290 138628 454300
rect 140812 444500 140868 476588
rect 140924 466138 140980 477260
rect 141036 475524 141092 480620
rect 141036 475458 141092 475468
rect 141932 475524 141988 475534
rect 140924 466072 140980 466082
rect 140812 444434 140868 444444
rect 132018 442294 132114 442350
rect 132170 442294 132238 442350
rect 132294 442294 132362 442350
rect 132418 442294 132486 442350
rect 132542 442294 132638 442350
rect 132018 442226 132638 442294
rect 132018 442170 132114 442226
rect 132170 442170 132238 442226
rect 132294 442170 132362 442226
rect 132418 442170 132486 442226
rect 132542 442170 132638 442226
rect 132018 442102 132638 442170
rect 132018 442046 132114 442102
rect 132170 442046 132238 442102
rect 132294 442046 132362 442102
rect 132418 442046 132486 442102
rect 132542 442046 132638 442102
rect 132018 441978 132638 442046
rect 132018 441922 132114 441978
rect 132170 441922 132238 441978
rect 132294 441922 132362 441978
rect 132418 441922 132486 441978
rect 132542 441922 132638 441978
rect 132018 424350 132638 441922
rect 141932 433076 141988 475468
rect 142044 457940 142100 481292
rect 142044 457874 142100 457884
rect 142156 461188 142212 461198
rect 142156 450996 142212 461132
rect 142156 450930 142212 450940
rect 143612 450436 143668 493388
rect 148448 490350 148768 490384
rect 148448 490294 148518 490350
rect 148574 490294 148642 490350
rect 148698 490294 148768 490350
rect 148448 490226 148768 490294
rect 148448 490170 148518 490226
rect 148574 490170 148642 490226
rect 148698 490170 148768 490226
rect 148448 490102 148768 490170
rect 148448 490046 148518 490102
rect 148574 490046 148642 490102
rect 148698 490046 148768 490102
rect 148448 489978 148768 490046
rect 148448 489922 148518 489978
rect 148574 489922 148642 489978
rect 148698 489922 148768 489978
rect 148448 489888 148768 489922
rect 159018 490350 159638 507922
rect 159018 490294 159114 490350
rect 159170 490294 159238 490350
rect 159294 490294 159362 490350
rect 159418 490294 159486 490350
rect 159542 490294 159638 490350
rect 159018 490226 159638 490294
rect 159018 490170 159114 490226
rect 159170 490170 159238 490226
rect 159294 490170 159362 490226
rect 159418 490170 159486 490226
rect 159542 490170 159638 490226
rect 159018 490102 159638 490170
rect 159018 490046 159114 490102
rect 159170 490046 159238 490102
rect 159294 490046 159362 490102
rect 159418 490046 159486 490102
rect 159542 490046 159638 490102
rect 159018 489978 159638 490046
rect 159018 489922 159114 489978
rect 159170 489922 159238 489978
rect 159294 489922 159362 489978
rect 159418 489922 159486 489978
rect 159542 489922 159638 489978
rect 143724 480452 143780 480462
rect 143724 459172 143780 480396
rect 148448 472350 148768 472384
rect 148448 472294 148518 472350
rect 148574 472294 148642 472350
rect 148698 472294 148768 472350
rect 148448 472226 148768 472294
rect 148448 472170 148518 472226
rect 148574 472170 148642 472226
rect 148698 472170 148768 472226
rect 148448 472102 148768 472170
rect 148448 472046 148518 472102
rect 148574 472046 148642 472102
rect 148698 472046 148768 472102
rect 148448 471978 148768 472046
rect 148448 471922 148518 471978
rect 148574 471922 148642 471978
rect 148698 471922 148768 471978
rect 148448 471888 148768 471922
rect 159018 472350 159638 489922
rect 159018 472294 159114 472350
rect 159170 472294 159238 472350
rect 159294 472294 159362 472350
rect 159418 472294 159486 472350
rect 159542 472294 159638 472350
rect 159018 472226 159638 472294
rect 159018 472170 159114 472226
rect 159170 472170 159238 472226
rect 159294 472170 159362 472226
rect 159418 472170 159486 472226
rect 159542 472170 159638 472226
rect 159018 472102 159638 472170
rect 159018 472046 159114 472102
rect 159170 472046 159238 472102
rect 159294 472046 159362 472102
rect 159418 472046 159486 472102
rect 159542 472046 159638 472102
rect 159018 471978 159638 472046
rect 159018 471922 159114 471978
rect 159170 471922 159238 471978
rect 159294 471922 159362 471978
rect 159418 471922 159486 471978
rect 159542 471922 159638 471978
rect 144396 471268 144452 471278
rect 144396 469558 144452 471212
rect 144396 469492 144452 469502
rect 143724 459106 143780 459116
rect 143612 450370 143668 450380
rect 159018 454350 159638 471922
rect 162738 532350 163358 542754
rect 162738 532294 162834 532350
rect 162890 532294 162958 532350
rect 163014 532294 163082 532350
rect 163138 532294 163206 532350
rect 163262 532294 163358 532350
rect 162738 532226 163358 532294
rect 162738 532170 162834 532226
rect 162890 532170 162958 532226
rect 163014 532170 163082 532226
rect 163138 532170 163206 532226
rect 163262 532170 163358 532226
rect 162738 532102 163358 532170
rect 162738 532046 162834 532102
rect 162890 532046 162958 532102
rect 163014 532046 163082 532102
rect 163138 532046 163206 532102
rect 163262 532046 163358 532102
rect 162738 531978 163358 532046
rect 162738 531922 162834 531978
rect 162890 531922 162958 531978
rect 163014 531922 163082 531978
rect 163138 531922 163206 531978
rect 163262 531922 163358 531978
rect 162738 514350 163358 531922
rect 163808 532350 164128 532384
rect 163808 532294 163878 532350
rect 163934 532294 164002 532350
rect 164058 532294 164128 532350
rect 163808 532226 164128 532294
rect 163808 532170 163878 532226
rect 163934 532170 164002 532226
rect 164058 532170 164128 532226
rect 163808 532102 164128 532170
rect 163808 532046 163878 532102
rect 163934 532046 164002 532102
rect 164058 532046 164128 532102
rect 163808 531978 164128 532046
rect 163808 531922 163878 531978
rect 163934 531922 164002 531978
rect 164058 531922 164128 531978
rect 163808 531888 164128 531922
rect 162738 514294 162834 514350
rect 162890 514294 162958 514350
rect 163014 514294 163082 514350
rect 163138 514294 163206 514350
rect 163262 514294 163358 514350
rect 162738 514226 163358 514294
rect 162738 514170 162834 514226
rect 162890 514170 162958 514226
rect 163014 514170 163082 514226
rect 163138 514170 163206 514226
rect 163262 514170 163358 514226
rect 162738 514102 163358 514170
rect 162738 514046 162834 514102
rect 162890 514046 162958 514102
rect 163014 514046 163082 514102
rect 163138 514046 163206 514102
rect 163262 514046 163358 514102
rect 162738 513978 163358 514046
rect 162738 513922 162834 513978
rect 162890 513922 162958 513978
rect 163014 513922 163082 513978
rect 163138 513922 163206 513978
rect 163262 513922 163358 513978
rect 162738 496350 163358 513922
rect 188972 503300 189028 549836
rect 189084 506772 189140 551180
rect 189196 548548 189252 548558
rect 189196 522116 189252 548492
rect 189196 522050 189252 522060
rect 189420 545188 189476 545198
rect 189420 521556 189476 545132
rect 189420 521490 189476 521500
rect 189738 544350 190358 561922
rect 189738 544294 189834 544350
rect 189890 544294 189958 544350
rect 190014 544294 190082 544350
rect 190138 544294 190206 544350
rect 190262 544294 190358 544350
rect 189738 544226 190358 544294
rect 189738 544170 189834 544226
rect 189890 544170 189958 544226
rect 190014 544170 190082 544226
rect 190138 544170 190206 544226
rect 190262 544170 190358 544226
rect 189738 544102 190358 544170
rect 189738 544046 189834 544102
rect 189890 544046 189958 544102
rect 190014 544046 190082 544102
rect 190138 544046 190206 544102
rect 190262 544046 190358 544102
rect 189738 543978 190358 544046
rect 189738 543922 189834 543978
rect 189890 543922 189958 543978
rect 190014 543922 190082 543978
rect 190138 543922 190206 543978
rect 190262 543922 190358 543978
rect 189738 526350 190358 543922
rect 189738 526294 189834 526350
rect 189890 526294 189958 526350
rect 190014 526294 190082 526350
rect 190138 526294 190206 526350
rect 190262 526294 190358 526350
rect 189738 526226 190358 526294
rect 189738 526170 189834 526226
rect 189890 526170 189958 526226
rect 190014 526170 190082 526226
rect 190138 526170 190206 526226
rect 190262 526170 190358 526226
rect 189738 526102 190358 526170
rect 189738 526046 189834 526102
rect 189890 526046 189958 526102
rect 190014 526046 190082 526102
rect 190138 526046 190206 526102
rect 190262 526046 190358 526102
rect 189738 525978 190358 526046
rect 189738 525922 189834 525978
rect 189890 525922 189958 525978
rect 190014 525922 190082 525978
rect 190138 525922 190206 525978
rect 190262 525922 190358 525978
rect 189084 506706 189140 506716
rect 189738 508350 190358 525922
rect 189738 508294 189834 508350
rect 189890 508294 189958 508350
rect 190014 508294 190082 508350
rect 190138 508294 190206 508350
rect 190262 508294 190358 508350
rect 189738 508226 190358 508294
rect 189738 508170 189834 508226
rect 189890 508170 189958 508226
rect 190014 508170 190082 508226
rect 190138 508170 190206 508226
rect 190262 508170 190358 508226
rect 189738 508102 190358 508170
rect 189738 508046 189834 508102
rect 189890 508046 189958 508102
rect 190014 508046 190082 508102
rect 190138 508046 190206 508102
rect 190262 508046 190358 508102
rect 189738 507978 190358 508046
rect 189738 507922 189834 507978
rect 189890 507922 189958 507978
rect 190014 507922 190082 507978
rect 190138 507922 190206 507978
rect 190262 507922 190358 507978
rect 188972 503234 189028 503244
rect 162738 496294 162834 496350
rect 162890 496294 162958 496350
rect 163014 496294 163082 496350
rect 163138 496294 163206 496350
rect 163262 496294 163358 496350
rect 162738 496226 163358 496294
rect 162738 496170 162834 496226
rect 162890 496170 162958 496226
rect 163014 496170 163082 496226
rect 163138 496170 163206 496226
rect 163262 496170 163358 496226
rect 162738 496102 163358 496170
rect 162738 496046 162834 496102
rect 162890 496046 162958 496102
rect 163014 496046 163082 496102
rect 163138 496046 163206 496102
rect 163262 496046 163358 496102
rect 162738 495978 163358 496046
rect 162738 495922 162834 495978
rect 162890 495922 162958 495978
rect 163014 495922 163082 495978
rect 163138 495922 163206 495978
rect 163262 495922 163358 495978
rect 162738 478350 163358 495922
rect 179168 490350 179488 490384
rect 179168 490294 179238 490350
rect 179294 490294 179362 490350
rect 179418 490294 179488 490350
rect 179168 490226 179488 490294
rect 179168 490170 179238 490226
rect 179294 490170 179362 490226
rect 179418 490170 179488 490226
rect 179168 490102 179488 490170
rect 179168 490046 179238 490102
rect 179294 490046 179362 490102
rect 179418 490046 179488 490102
rect 179168 489978 179488 490046
rect 179168 489922 179238 489978
rect 179294 489922 179362 489978
rect 179418 489922 179488 489978
rect 179168 489888 179488 489922
rect 189738 490350 190358 507922
rect 189738 490294 189834 490350
rect 189890 490294 189958 490350
rect 190014 490294 190082 490350
rect 190138 490294 190206 490350
rect 190262 490294 190358 490350
rect 189738 490226 190358 490294
rect 189738 490170 189834 490226
rect 189890 490170 189958 490226
rect 190014 490170 190082 490226
rect 190138 490170 190206 490226
rect 190262 490170 190358 490226
rect 189738 490102 190358 490170
rect 189738 490046 189834 490102
rect 189890 490046 189958 490102
rect 190014 490046 190082 490102
rect 190138 490046 190206 490102
rect 190262 490046 190358 490102
rect 189738 489978 190358 490046
rect 189738 489922 189834 489978
rect 189890 489922 189958 489978
rect 190014 489922 190082 489978
rect 190138 489922 190206 489978
rect 190262 489922 190358 489978
rect 189084 482692 189140 482702
rect 188972 478660 189028 478670
rect 162738 478294 162834 478350
rect 162890 478294 162958 478350
rect 163014 478294 163082 478350
rect 163138 478294 163206 478350
rect 163262 478294 163358 478350
rect 162738 478226 163358 478294
rect 162738 478170 162834 478226
rect 162890 478170 162958 478226
rect 163014 478170 163082 478226
rect 163138 478170 163206 478226
rect 163262 478170 163358 478226
rect 162738 478102 163358 478170
rect 162738 478046 162834 478102
rect 162890 478046 162958 478102
rect 163014 478046 163082 478102
rect 163138 478046 163206 478102
rect 163262 478046 163358 478102
rect 162738 477978 163358 478046
rect 162738 477922 162834 477978
rect 162890 477922 162958 477978
rect 163014 477922 163082 477978
rect 163138 477922 163206 477978
rect 163262 477922 163358 477978
rect 162738 460350 163358 477922
rect 163808 478350 164128 478384
rect 163808 478294 163878 478350
rect 163934 478294 164002 478350
rect 164058 478294 164128 478350
rect 163808 478226 164128 478294
rect 163808 478170 163878 478226
rect 163934 478170 164002 478226
rect 164058 478170 164128 478226
rect 163808 478102 164128 478170
rect 163808 478046 163878 478102
rect 163934 478046 164002 478102
rect 164058 478046 164128 478102
rect 163808 477978 164128 478046
rect 163808 477922 163878 477978
rect 163934 477922 164002 477978
rect 164058 477922 164128 477978
rect 163808 477888 164128 477922
rect 179168 472350 179488 472384
rect 179168 472294 179238 472350
rect 179294 472294 179362 472350
rect 179418 472294 179488 472350
rect 179168 472226 179488 472294
rect 179168 472170 179238 472226
rect 179294 472170 179362 472226
rect 179418 472170 179488 472226
rect 179168 472102 179488 472170
rect 179168 472046 179238 472102
rect 179294 472046 179362 472102
rect 179418 472046 179488 472102
rect 179168 471978 179488 472046
rect 179168 471922 179238 471978
rect 179294 471922 179362 471978
rect 179418 471922 179488 471978
rect 179168 471888 179488 471922
rect 188972 461188 189028 478604
rect 189084 467908 189140 482636
rect 189532 475972 189588 475982
rect 189532 475498 189588 475916
rect 189532 475432 189588 475442
rect 189532 473956 189588 473966
rect 189532 473878 189588 473900
rect 189532 473812 189588 473822
rect 189084 467842 189140 467852
rect 189738 472350 190358 489922
rect 189738 472294 189834 472350
rect 189890 472294 189958 472350
rect 190014 472294 190082 472350
rect 190138 472294 190206 472350
rect 190262 472294 190358 472350
rect 189738 472226 190358 472294
rect 189738 472170 189834 472226
rect 189890 472170 189958 472226
rect 190014 472170 190082 472226
rect 190138 472170 190206 472226
rect 190262 472170 190358 472226
rect 189738 472102 190358 472170
rect 189738 472046 189834 472102
rect 189890 472046 189958 472102
rect 190014 472046 190082 472102
rect 190138 472046 190206 472102
rect 190262 472046 190358 472102
rect 189738 471978 190358 472046
rect 189738 471922 189834 471978
rect 189890 471922 189958 471978
rect 190014 471922 190082 471978
rect 190138 471922 190206 471978
rect 190262 471922 190358 471978
rect 188972 461122 189028 461132
rect 162738 460294 162834 460350
rect 162890 460294 162958 460350
rect 163014 460294 163082 460350
rect 163138 460294 163206 460350
rect 163262 460294 163358 460350
rect 162738 460226 163358 460294
rect 162738 460170 162834 460226
rect 162890 460170 162958 460226
rect 163014 460170 163082 460226
rect 163138 460170 163206 460226
rect 163262 460170 163358 460226
rect 162738 460102 163358 460170
rect 162738 460046 162834 460102
rect 162890 460046 162958 460102
rect 163014 460046 163082 460102
rect 163138 460046 163206 460102
rect 163262 460046 163358 460102
rect 162738 459978 163358 460046
rect 162738 459922 162834 459978
rect 162890 459922 162958 459978
rect 163014 459922 163082 459978
rect 163138 459922 163206 459978
rect 163262 459922 163358 459978
rect 160860 458052 160916 458062
rect 160860 456932 160916 457996
rect 160860 456866 160916 456876
rect 159018 454294 159114 454350
rect 159170 454294 159238 454350
rect 159294 454294 159362 454350
rect 159418 454294 159486 454350
rect 159542 454294 159638 454350
rect 159018 454226 159638 454294
rect 159018 454170 159114 454226
rect 159170 454170 159238 454226
rect 159294 454170 159362 454226
rect 159418 454170 159486 454226
rect 159542 454170 159638 454226
rect 159018 454102 159638 454170
rect 159018 454046 159114 454102
rect 159170 454046 159238 454102
rect 159294 454046 159362 454102
rect 159418 454046 159486 454102
rect 159542 454046 159638 454102
rect 159018 453978 159638 454046
rect 159018 453922 159114 453978
rect 159170 453922 159238 453978
rect 159294 453922 159362 453978
rect 159418 453922 159486 453978
rect 159542 453922 159638 453978
rect 141932 433010 141988 433020
rect 159018 436350 159638 453922
rect 159018 436294 159114 436350
rect 159170 436294 159238 436350
rect 159294 436294 159362 436350
rect 159418 436294 159486 436350
rect 159542 436294 159638 436350
rect 159018 436226 159638 436294
rect 159018 436170 159114 436226
rect 159170 436170 159238 436226
rect 159294 436170 159362 436226
rect 159418 436170 159486 436226
rect 159542 436170 159638 436226
rect 159018 436102 159638 436170
rect 159018 436046 159114 436102
rect 159170 436046 159238 436102
rect 159294 436046 159362 436102
rect 159418 436046 159486 436102
rect 159542 436046 159638 436102
rect 159018 435978 159638 436046
rect 159018 435922 159114 435978
rect 159170 435922 159238 435978
rect 159294 435922 159362 435978
rect 159418 435922 159486 435978
rect 159542 435922 159638 435978
rect 132018 424294 132114 424350
rect 132170 424294 132238 424350
rect 132294 424294 132362 424350
rect 132418 424294 132486 424350
rect 132542 424294 132638 424350
rect 132018 424226 132638 424294
rect 132018 424170 132114 424226
rect 132170 424170 132238 424226
rect 132294 424170 132362 424226
rect 132418 424170 132486 424226
rect 132542 424170 132638 424226
rect 132018 424102 132638 424170
rect 132018 424046 132114 424102
rect 132170 424046 132238 424102
rect 132294 424046 132362 424102
rect 132418 424046 132486 424102
rect 132542 424046 132638 424102
rect 132018 423978 132638 424046
rect 132018 423922 132114 423978
rect 132170 423922 132238 423978
rect 132294 423922 132362 423978
rect 132418 423922 132486 423978
rect 132542 423922 132638 423978
rect 132018 406350 132638 423922
rect 148448 418350 148768 418384
rect 148448 418294 148518 418350
rect 148574 418294 148642 418350
rect 148698 418294 148768 418350
rect 148448 418226 148768 418294
rect 148448 418170 148518 418226
rect 148574 418170 148642 418226
rect 148698 418170 148768 418226
rect 148448 418102 148768 418170
rect 148448 418046 148518 418102
rect 148574 418046 148642 418102
rect 148698 418046 148768 418102
rect 148448 417978 148768 418046
rect 148448 417922 148518 417978
rect 148574 417922 148642 417978
rect 148698 417922 148768 417978
rect 148448 417888 148768 417922
rect 159018 418350 159638 435922
rect 159018 418294 159114 418350
rect 159170 418294 159238 418350
rect 159294 418294 159362 418350
rect 159418 418294 159486 418350
rect 159542 418294 159638 418350
rect 159018 418226 159638 418294
rect 159018 418170 159114 418226
rect 159170 418170 159238 418226
rect 159294 418170 159362 418226
rect 159418 418170 159486 418226
rect 159542 418170 159638 418226
rect 159018 418102 159638 418170
rect 159018 418046 159114 418102
rect 159170 418046 159238 418102
rect 159294 418046 159362 418102
rect 159418 418046 159486 418102
rect 159542 418046 159638 418102
rect 159018 417978 159638 418046
rect 159018 417922 159114 417978
rect 159170 417922 159238 417978
rect 159294 417922 159362 417978
rect 159418 417922 159486 417978
rect 159542 417922 159638 417978
rect 141036 412804 141092 412814
rect 141036 412498 141092 412748
rect 144060 412804 144116 412814
rect 144060 412678 144116 412748
rect 144060 412612 144116 412622
rect 141036 412432 141092 412442
rect 132018 406294 132114 406350
rect 132170 406294 132238 406350
rect 132294 406294 132362 406350
rect 132418 406294 132486 406350
rect 132542 406294 132638 406350
rect 132018 406226 132638 406294
rect 132018 406170 132114 406226
rect 132170 406170 132238 406226
rect 132294 406170 132362 406226
rect 132418 406170 132486 406226
rect 132542 406170 132638 406226
rect 132018 406102 132638 406170
rect 132018 406046 132114 406102
rect 132170 406046 132238 406102
rect 132294 406046 132362 406102
rect 132418 406046 132486 406102
rect 132542 406046 132638 406102
rect 132018 405978 132638 406046
rect 132018 405922 132114 405978
rect 132170 405922 132238 405978
rect 132294 405922 132362 405978
rect 132418 405922 132486 405978
rect 132542 405922 132638 405978
rect 132018 388350 132638 405922
rect 135212 411460 135268 411470
rect 132018 388294 132114 388350
rect 132170 388294 132238 388350
rect 132294 388294 132362 388350
rect 132418 388294 132486 388350
rect 132542 388294 132638 388350
rect 132018 388226 132638 388294
rect 132018 388170 132114 388226
rect 132170 388170 132238 388226
rect 132294 388170 132362 388226
rect 132418 388170 132486 388226
rect 132542 388170 132638 388226
rect 132018 388102 132638 388170
rect 132018 388046 132114 388102
rect 132170 388046 132238 388102
rect 132294 388046 132362 388102
rect 132418 388046 132486 388102
rect 132542 388046 132638 388102
rect 132018 387978 132638 388046
rect 132018 387922 132114 387978
rect 132170 387922 132238 387978
rect 132294 387922 132362 387978
rect 132418 387922 132486 387978
rect 132542 387922 132638 387978
rect 132018 370350 132638 387922
rect 133532 401380 133588 401390
rect 133532 380772 133588 401324
rect 135212 393058 135268 411404
rect 142716 410116 142772 410126
rect 136108 406756 136164 406766
rect 136108 399718 136164 406700
rect 136108 399652 136164 399662
rect 141036 403396 141092 403406
rect 135212 392992 135268 393002
rect 133532 380706 133588 380716
rect 141036 377076 141092 403340
rect 141036 377010 141092 377020
rect 142716 374276 142772 410060
rect 144284 409978 144340 409988
rect 144284 409892 144340 409922
rect 144284 409826 144340 409836
rect 144284 408436 144340 408446
rect 144284 408358 144340 408380
rect 144284 408292 144340 408302
rect 144396 407316 144452 407326
rect 144396 406738 144452 407260
rect 144396 406672 144452 406682
rect 144284 406644 144340 406654
rect 144284 404218 144340 406588
rect 144284 404152 144340 404162
rect 142716 374210 142772 374220
rect 143612 402724 143668 402734
rect 132018 370294 132114 370350
rect 132170 370294 132238 370350
rect 132294 370294 132362 370350
rect 132418 370294 132486 370350
rect 132542 370294 132638 370350
rect 132018 370226 132638 370294
rect 132018 370170 132114 370226
rect 132170 370170 132238 370226
rect 132294 370170 132362 370226
rect 132418 370170 132486 370226
rect 132542 370170 132638 370226
rect 132018 370102 132638 370170
rect 132018 370046 132114 370102
rect 132170 370046 132238 370102
rect 132294 370046 132362 370102
rect 132418 370046 132486 370102
rect 132542 370046 132638 370102
rect 132018 369978 132638 370046
rect 132018 369922 132114 369978
rect 132170 369922 132238 369978
rect 132294 369922 132362 369978
rect 132418 369922 132486 369978
rect 132542 369922 132638 369978
rect 132018 352350 132638 369922
rect 143612 364196 143668 402668
rect 148448 400350 148768 400384
rect 148448 400294 148518 400350
rect 148574 400294 148642 400350
rect 148698 400294 148768 400350
rect 148448 400226 148768 400294
rect 148448 400170 148518 400226
rect 148574 400170 148642 400226
rect 148698 400170 148768 400226
rect 148448 400102 148768 400170
rect 148448 400046 148518 400102
rect 148574 400046 148642 400102
rect 148698 400046 148768 400102
rect 148448 399978 148768 400046
rect 148448 399922 148518 399978
rect 148574 399922 148642 399978
rect 148698 399922 148768 399978
rect 148448 399888 148768 399922
rect 159018 400350 159638 417922
rect 159018 400294 159114 400350
rect 159170 400294 159238 400350
rect 159294 400294 159362 400350
rect 159418 400294 159486 400350
rect 159542 400294 159638 400350
rect 159018 400226 159638 400294
rect 159018 400170 159114 400226
rect 159170 400170 159238 400226
rect 159294 400170 159362 400226
rect 159418 400170 159486 400226
rect 159542 400170 159638 400226
rect 159018 400102 159638 400170
rect 159018 400046 159114 400102
rect 159170 400046 159238 400102
rect 159294 400046 159362 400102
rect 159418 400046 159486 400102
rect 159542 400046 159638 400102
rect 159018 399978 159638 400046
rect 159018 399922 159114 399978
rect 159170 399922 159238 399978
rect 159294 399922 159362 399978
rect 159418 399922 159486 399978
rect 159542 399922 159638 399978
rect 143612 364130 143668 364140
rect 159018 382350 159638 399922
rect 159018 382294 159114 382350
rect 159170 382294 159238 382350
rect 159294 382294 159362 382350
rect 159418 382294 159486 382350
rect 159542 382294 159638 382350
rect 159018 382226 159638 382294
rect 159018 382170 159114 382226
rect 159170 382170 159238 382226
rect 159294 382170 159362 382226
rect 159418 382170 159486 382226
rect 159542 382170 159638 382226
rect 159018 382102 159638 382170
rect 159018 382046 159114 382102
rect 159170 382046 159238 382102
rect 159294 382046 159362 382102
rect 159418 382046 159486 382102
rect 159542 382046 159638 382102
rect 159018 381978 159638 382046
rect 159018 381922 159114 381978
rect 159170 381922 159238 381978
rect 159294 381922 159362 381978
rect 159418 381922 159486 381978
rect 159542 381922 159638 381978
rect 159018 364350 159638 381922
rect 159018 364294 159114 364350
rect 159170 364294 159238 364350
rect 159294 364294 159362 364350
rect 159418 364294 159486 364350
rect 159542 364294 159638 364350
rect 159018 364226 159638 364294
rect 159018 364170 159114 364226
rect 159170 364170 159238 364226
rect 159294 364170 159362 364226
rect 159418 364170 159486 364226
rect 159542 364170 159638 364226
rect 132018 352294 132114 352350
rect 132170 352294 132238 352350
rect 132294 352294 132362 352350
rect 132418 352294 132486 352350
rect 132542 352294 132638 352350
rect 132018 352226 132638 352294
rect 132018 352170 132114 352226
rect 132170 352170 132238 352226
rect 132294 352170 132362 352226
rect 132418 352170 132486 352226
rect 132542 352170 132638 352226
rect 132018 352102 132638 352170
rect 132018 352046 132114 352102
rect 132170 352046 132238 352102
rect 132294 352046 132362 352102
rect 132418 352046 132486 352102
rect 132542 352046 132638 352102
rect 132018 351978 132638 352046
rect 132018 351922 132114 351978
rect 132170 351922 132238 351978
rect 132294 351922 132362 351978
rect 132418 351922 132486 351978
rect 132542 351922 132638 351978
rect 130060 341758 130116 341768
rect 130060 339332 130116 341702
rect 130060 339266 130116 339276
rect 128298 328294 128394 328350
rect 128450 328294 128518 328350
rect 128574 328294 128642 328350
rect 128698 328294 128766 328350
rect 128822 328294 128918 328350
rect 128298 328226 128918 328294
rect 128298 328170 128394 328226
rect 128450 328170 128518 328226
rect 128574 328170 128642 328226
rect 128698 328170 128766 328226
rect 128822 328170 128918 328226
rect 128298 328102 128918 328170
rect 128298 328046 128394 328102
rect 128450 328046 128518 328102
rect 128574 328046 128642 328102
rect 128698 328046 128766 328102
rect 128822 328046 128918 328102
rect 128298 327978 128918 328046
rect 128298 327922 128394 327978
rect 128450 327922 128518 327978
rect 128574 327922 128642 327978
rect 128698 327922 128766 327978
rect 128822 327922 128918 327978
rect 97578 310294 97674 310350
rect 97730 310294 97798 310350
rect 97854 310294 97922 310350
rect 97978 310294 98046 310350
rect 98102 310294 98198 310350
rect 97578 310226 98198 310294
rect 97578 310170 97674 310226
rect 97730 310170 97798 310226
rect 97854 310170 97922 310226
rect 97978 310170 98046 310226
rect 98102 310170 98198 310226
rect 97578 310102 98198 310170
rect 97578 310046 97674 310102
rect 97730 310046 97798 310102
rect 97854 310046 97922 310102
rect 97978 310046 98046 310102
rect 98102 310046 98198 310102
rect 97578 309978 98198 310046
rect 97578 309922 97674 309978
rect 97730 309922 97798 309978
rect 97854 309922 97922 309978
rect 97978 309922 98046 309978
rect 98102 309922 98198 309978
rect 70578 298294 70674 298350
rect 70730 298294 70798 298350
rect 70854 298294 70922 298350
rect 70978 298294 71046 298350
rect 71102 298294 71198 298350
rect 70578 298226 71198 298294
rect 70578 298170 70674 298226
rect 70730 298170 70798 298226
rect 70854 298170 70922 298226
rect 70978 298170 71046 298226
rect 71102 298170 71198 298226
rect 70578 298102 71198 298170
rect 70578 298046 70674 298102
rect 70730 298046 70798 298102
rect 70854 298046 70922 298102
rect 70978 298046 71046 298102
rect 71102 298046 71198 298102
rect 70578 297978 71198 298046
rect 70578 297922 70674 297978
rect 70730 297922 70798 297978
rect 70854 297922 70922 297978
rect 70978 297922 71046 297978
rect 71102 297922 71198 297978
rect 70578 280350 71198 297922
rect 97578 292350 98198 309922
rect 97578 292294 97674 292350
rect 97730 292294 97798 292350
rect 97854 292294 97922 292350
rect 97978 292294 98046 292350
rect 98102 292294 98198 292350
rect 97578 292226 98198 292294
rect 97578 292170 97674 292226
rect 97730 292170 97798 292226
rect 97854 292170 97922 292226
rect 97978 292170 98046 292226
rect 98102 292170 98198 292226
rect 97578 292102 98198 292170
rect 97578 292046 97674 292102
rect 97730 292046 97798 292102
rect 97854 292046 97922 292102
rect 97978 292046 98046 292102
rect 98102 292046 98198 292102
rect 97578 291978 98198 292046
rect 97578 291922 97674 291978
rect 97730 291922 97798 291978
rect 97854 291922 97922 291978
rect 97978 291922 98046 291978
rect 98102 291922 98198 291978
rect 70578 280294 70674 280350
rect 70730 280294 70798 280350
rect 70854 280294 70922 280350
rect 70978 280294 71046 280350
rect 71102 280294 71198 280350
rect 70578 280226 71198 280294
rect 70578 280170 70674 280226
rect 70730 280170 70798 280226
rect 70854 280170 70922 280226
rect 70978 280170 71046 280226
rect 71102 280170 71198 280226
rect 70578 280102 71198 280170
rect 70578 280046 70674 280102
rect 70730 280046 70798 280102
rect 70854 280046 70922 280102
rect 70978 280046 71046 280102
rect 71102 280046 71198 280102
rect 70578 279978 71198 280046
rect 70578 279922 70674 279978
rect 70730 279922 70798 279978
rect 70854 279922 70922 279978
rect 70978 279922 71046 279978
rect 71102 279922 71198 279978
rect 66858 256294 66954 256350
rect 67010 256294 67078 256350
rect 67134 256294 67202 256350
rect 67258 256294 67326 256350
rect 67382 256294 67478 256350
rect 66858 256226 67478 256294
rect 66858 256170 66954 256226
rect 67010 256170 67078 256226
rect 67134 256170 67202 256226
rect 67258 256170 67326 256226
rect 67382 256170 67478 256226
rect 66858 256102 67478 256170
rect 66858 256046 66954 256102
rect 67010 256046 67078 256102
rect 67134 256046 67202 256102
rect 67258 256046 67326 256102
rect 67382 256046 67478 256102
rect 66858 255978 67478 256046
rect 66858 255922 66954 255978
rect 67010 255922 67078 255978
rect 67134 255922 67202 255978
rect 67258 255922 67326 255978
rect 67382 255922 67478 255978
rect 64652 245186 64708 245196
rect 36138 238294 36234 238350
rect 36290 238294 36358 238350
rect 36414 238294 36482 238350
rect 36538 238294 36606 238350
rect 36662 238294 36758 238350
rect 36138 238226 36758 238294
rect 36138 238170 36234 238226
rect 36290 238170 36358 238226
rect 36414 238170 36482 238226
rect 36538 238170 36606 238226
rect 36662 238170 36758 238226
rect 36138 238102 36758 238170
rect 36138 238046 36234 238102
rect 36290 238046 36358 238102
rect 36414 238046 36482 238102
rect 36538 238046 36606 238102
rect 36662 238046 36758 238102
rect 36138 237978 36758 238046
rect 36138 237922 36234 237978
rect 36290 237922 36358 237978
rect 36414 237922 36482 237978
rect 36538 237922 36606 237978
rect 36662 237922 36758 237978
rect 36138 220350 36758 237922
rect 36138 220294 36234 220350
rect 36290 220294 36358 220350
rect 36414 220294 36482 220350
rect 36538 220294 36606 220350
rect 36662 220294 36758 220350
rect 36138 220226 36758 220294
rect 36138 220170 36234 220226
rect 36290 220170 36358 220226
rect 36414 220170 36482 220226
rect 36538 220170 36606 220226
rect 36662 220170 36758 220226
rect 36138 220102 36758 220170
rect 36138 220046 36234 220102
rect 36290 220046 36358 220102
rect 36414 220046 36482 220102
rect 36538 220046 36606 220102
rect 36662 220046 36758 220102
rect 36138 219978 36758 220046
rect 36138 219922 36234 219978
rect 36290 219922 36358 219978
rect 36414 219922 36482 219978
rect 36538 219922 36606 219978
rect 36662 219922 36758 219978
rect 9138 208294 9234 208350
rect 9290 208294 9358 208350
rect 9414 208294 9482 208350
rect 9538 208294 9606 208350
rect 9662 208294 9758 208350
rect 9138 208226 9758 208294
rect 9138 208170 9234 208226
rect 9290 208170 9358 208226
rect 9414 208170 9482 208226
rect 9538 208170 9606 208226
rect 9662 208170 9758 208226
rect 9138 208102 9758 208170
rect 9138 208046 9234 208102
rect 9290 208046 9358 208102
rect 9414 208046 9482 208102
rect 9538 208046 9606 208102
rect 9662 208046 9758 208102
rect 9138 207978 9758 208046
rect 9138 207922 9234 207978
rect 9290 207922 9358 207978
rect 9414 207922 9482 207978
rect 9538 207922 9606 207978
rect 9662 207922 9758 207978
rect 9138 190350 9758 207922
rect 20076 210420 20132 210430
rect 18396 199018 18452 199034
rect 18396 198930 18452 198940
rect 20076 194516 20132 210364
rect 24448 202350 24768 202384
rect 24448 202294 24518 202350
rect 24574 202294 24642 202350
rect 24698 202294 24768 202350
rect 24448 202226 24768 202294
rect 24448 202170 24518 202226
rect 24574 202170 24642 202226
rect 24698 202170 24768 202226
rect 24448 202102 24768 202170
rect 24448 202046 24518 202102
rect 24574 202046 24642 202102
rect 24698 202046 24768 202102
rect 24448 201978 24768 202046
rect 24448 201922 24518 201978
rect 24574 201922 24642 201978
rect 24698 201922 24768 201978
rect 24448 201888 24768 201922
rect 36138 202350 36758 219922
rect 66858 238350 67478 255922
rect 69692 265076 69748 265086
rect 69692 243236 69748 265020
rect 69692 243170 69748 243180
rect 70578 262350 71198 279922
rect 80332 282436 80388 282446
rect 80332 263060 80388 282380
rect 82012 281540 82068 281550
rect 80332 262994 80388 263004
rect 80444 265748 80500 265758
rect 70578 262294 70674 262350
rect 70730 262294 70798 262350
rect 70854 262294 70922 262350
rect 70978 262294 71046 262350
rect 71102 262294 71198 262350
rect 70578 262226 71198 262294
rect 70578 262170 70674 262226
rect 70730 262170 70798 262226
rect 70854 262170 70922 262226
rect 70978 262170 71046 262226
rect 71102 262170 71198 262226
rect 70578 262102 71198 262170
rect 70578 262046 70674 262102
rect 70730 262046 70798 262102
rect 70854 262046 70922 262102
rect 70978 262046 71046 262102
rect 71102 262046 71198 262102
rect 70578 261978 71198 262046
rect 70578 261922 70674 261978
rect 70730 261922 70798 261978
rect 70854 261922 70922 261978
rect 70978 261922 71046 261978
rect 71102 261922 71198 261978
rect 70578 244350 71198 261922
rect 80444 253558 80500 265692
rect 80444 253492 80500 253502
rect 81452 261268 81508 261278
rect 80556 252868 80612 252878
rect 80556 244916 80612 252812
rect 80556 244850 80612 244860
rect 70578 244294 70674 244350
rect 70730 244294 70798 244350
rect 70854 244294 70922 244350
rect 70978 244294 71046 244350
rect 71102 244294 71198 244350
rect 70578 244226 71198 244294
rect 70578 244170 70674 244226
rect 70730 244170 70798 244226
rect 70854 244170 70922 244226
rect 70978 244170 71046 244226
rect 71102 244170 71198 244226
rect 70578 244102 71198 244170
rect 70578 244046 70674 244102
rect 70730 244046 70798 244102
rect 70854 244046 70922 244102
rect 70978 244046 71046 244102
rect 71102 244046 71198 244102
rect 70578 243978 71198 244046
rect 70578 243922 70674 243978
rect 70730 243922 70798 243978
rect 70854 243922 70922 243978
rect 70978 243922 71046 243978
rect 71102 243922 71198 243978
rect 66858 238294 66954 238350
rect 67010 238294 67078 238350
rect 67134 238294 67202 238350
rect 67258 238294 67326 238350
rect 67382 238294 67478 238350
rect 66858 238226 67478 238294
rect 66858 238170 66954 238226
rect 67010 238170 67078 238226
rect 67134 238170 67202 238226
rect 67258 238170 67326 238226
rect 67382 238170 67478 238226
rect 66858 238102 67478 238170
rect 66858 238046 66954 238102
rect 67010 238046 67078 238102
rect 67134 238046 67202 238102
rect 67258 238046 67326 238102
rect 67382 238046 67478 238102
rect 66858 237978 67478 238046
rect 66858 237922 66954 237978
rect 67010 237922 67078 237978
rect 67134 237922 67202 237978
rect 67258 237922 67326 237978
rect 67382 237922 67478 237978
rect 66858 220350 67478 237922
rect 66858 220294 66954 220350
rect 67010 220294 67078 220350
rect 67134 220294 67202 220350
rect 67258 220294 67326 220350
rect 67382 220294 67478 220350
rect 66858 220226 67478 220294
rect 66858 220170 66954 220226
rect 67010 220170 67078 220226
rect 67134 220170 67202 220226
rect 67258 220170 67326 220226
rect 67382 220170 67478 220226
rect 66858 220102 67478 220170
rect 66858 220046 66954 220102
rect 67010 220046 67078 220102
rect 67134 220046 67202 220102
rect 67258 220046 67326 220102
rect 67382 220046 67478 220102
rect 66858 219978 67478 220046
rect 66858 219922 66954 219978
rect 67010 219922 67078 219978
rect 67134 219922 67202 219978
rect 67258 219922 67326 219978
rect 67382 219922 67478 219978
rect 64652 211092 64708 211102
rect 39808 208350 40128 208384
rect 39808 208294 39878 208350
rect 39934 208294 40002 208350
rect 40058 208294 40128 208350
rect 39808 208226 40128 208294
rect 39808 208170 39878 208226
rect 39934 208170 40002 208226
rect 40058 208170 40128 208226
rect 39808 208102 40128 208170
rect 39808 208046 39878 208102
rect 39934 208046 40002 208102
rect 40058 208046 40128 208102
rect 39808 207978 40128 208046
rect 39808 207922 39878 207978
rect 39934 207922 40002 207978
rect 40058 207922 40128 207978
rect 39808 207888 40128 207922
rect 36138 202294 36234 202350
rect 36290 202294 36358 202350
rect 36414 202294 36482 202350
rect 36538 202294 36606 202350
rect 36662 202294 36758 202350
rect 36138 202226 36758 202294
rect 36138 202170 36234 202226
rect 36290 202170 36358 202226
rect 36414 202170 36482 202226
rect 36538 202170 36606 202226
rect 36662 202170 36758 202226
rect 36138 202102 36758 202170
rect 36138 202046 36234 202102
rect 36290 202046 36358 202102
rect 36414 202046 36482 202102
rect 36538 202046 36606 202102
rect 36662 202046 36758 202102
rect 36138 201978 36758 202046
rect 36138 201922 36234 201978
rect 36290 201922 36358 201978
rect 36414 201922 36482 201978
rect 36538 201922 36606 201978
rect 36662 201922 36758 201978
rect 20636 196084 20692 196094
rect 20636 195058 20692 196028
rect 20636 194992 20692 195002
rect 20076 194450 20132 194460
rect 20300 194964 20356 194974
rect 20300 194158 20356 194908
rect 20300 194092 20356 194102
rect 9138 190294 9234 190350
rect 9290 190294 9358 190350
rect 9414 190294 9482 190350
rect 9538 190294 9606 190350
rect 9662 190294 9758 190350
rect 9138 190226 9758 190294
rect 9138 190170 9234 190226
rect 9290 190170 9358 190226
rect 9414 190170 9482 190226
rect 9538 190170 9606 190226
rect 9662 190170 9758 190226
rect 9138 190102 9758 190170
rect 9138 190046 9234 190102
rect 9290 190046 9358 190102
rect 9414 190046 9482 190102
rect 9538 190046 9606 190102
rect 9662 190046 9758 190102
rect 9138 189978 9758 190046
rect 9138 189922 9234 189978
rect 9290 189922 9358 189978
rect 9414 189922 9482 189978
rect 9538 189922 9606 189978
rect 9662 189922 9758 189978
rect 9138 172350 9758 189922
rect 20076 188244 20132 188254
rect 20076 186418 20132 188188
rect 20076 186352 20132 186362
rect 24448 184350 24768 184384
rect 24448 184294 24518 184350
rect 24574 184294 24642 184350
rect 24698 184294 24768 184350
rect 24448 184226 24768 184294
rect 24448 184170 24518 184226
rect 24574 184170 24642 184226
rect 24698 184170 24768 184226
rect 24448 184102 24768 184170
rect 24448 184046 24518 184102
rect 24574 184046 24642 184102
rect 24698 184046 24768 184102
rect 24448 183978 24768 184046
rect 24448 183922 24518 183978
rect 24574 183922 24642 183978
rect 24698 183922 24768 183978
rect 24448 183888 24768 183922
rect 36138 184350 36758 201922
rect 55168 202350 55488 202384
rect 55168 202294 55238 202350
rect 55294 202294 55362 202350
rect 55418 202294 55488 202350
rect 55168 202226 55488 202294
rect 55168 202170 55238 202226
rect 55294 202170 55362 202226
rect 55418 202170 55488 202226
rect 55168 202102 55488 202170
rect 55168 202046 55238 202102
rect 55294 202046 55362 202102
rect 55418 202046 55488 202102
rect 55168 201978 55488 202046
rect 55168 201922 55238 201978
rect 55294 201922 55362 201978
rect 55418 201922 55488 201978
rect 55168 201888 55488 201922
rect 64204 197204 64260 197214
rect 64204 196678 64260 197148
rect 64204 196612 64260 196622
rect 64204 195238 64260 195248
rect 64204 195122 64260 195132
rect 39808 190350 40128 190384
rect 39808 190294 39878 190350
rect 39934 190294 40002 190350
rect 40058 190294 40128 190350
rect 39808 190226 40128 190294
rect 39808 190170 39878 190226
rect 39934 190170 40002 190226
rect 40058 190170 40128 190226
rect 39808 190102 40128 190170
rect 39808 190046 39878 190102
rect 39934 190046 40002 190102
rect 40058 190046 40128 190102
rect 39808 189978 40128 190046
rect 39808 189922 39878 189978
rect 39934 189922 40002 189978
rect 40058 189922 40128 189978
rect 39808 189888 40128 189922
rect 64652 187124 64708 211036
rect 64652 187058 64708 187068
rect 66858 202350 67478 219922
rect 66858 202294 66954 202350
rect 67010 202294 67078 202350
rect 67134 202294 67202 202350
rect 67258 202294 67326 202350
rect 67382 202294 67478 202350
rect 66858 202226 67478 202294
rect 66858 202170 66954 202226
rect 67010 202170 67078 202226
rect 67134 202170 67202 202226
rect 67258 202170 67326 202226
rect 67382 202170 67478 202226
rect 66858 202102 67478 202170
rect 66858 202046 66954 202102
rect 67010 202046 67078 202102
rect 67134 202046 67202 202102
rect 67258 202046 67326 202102
rect 67382 202046 67478 202102
rect 66858 201978 67478 202046
rect 66858 201922 66954 201978
rect 67010 201922 67078 201978
rect 67134 201922 67202 201978
rect 67258 201922 67326 201978
rect 67382 201922 67478 201978
rect 36138 184294 36234 184350
rect 36290 184294 36358 184350
rect 36414 184294 36482 184350
rect 36538 184294 36606 184350
rect 36662 184294 36758 184350
rect 36138 184226 36758 184294
rect 36138 184170 36234 184226
rect 36290 184170 36358 184226
rect 36414 184170 36482 184226
rect 36538 184170 36606 184226
rect 36662 184170 36758 184226
rect 36138 184102 36758 184170
rect 36138 184046 36234 184102
rect 36290 184046 36358 184102
rect 36414 184046 36482 184102
rect 36538 184046 36606 184102
rect 36662 184046 36758 184102
rect 36138 183978 36758 184046
rect 36138 183922 36234 183978
rect 36290 183922 36358 183978
rect 36414 183922 36482 183978
rect 36538 183922 36606 183978
rect 36662 183922 36758 183978
rect 9138 172294 9234 172350
rect 9290 172294 9358 172350
rect 9414 172294 9482 172350
rect 9538 172294 9606 172350
rect 9662 172294 9758 172350
rect 9138 172226 9758 172294
rect 9138 172170 9234 172226
rect 9290 172170 9358 172226
rect 9414 172170 9482 172226
rect 9538 172170 9606 172226
rect 9662 172170 9758 172226
rect 9138 172102 9758 172170
rect 9138 172046 9234 172102
rect 9290 172046 9358 172102
rect 9414 172046 9482 172102
rect 9538 172046 9606 172102
rect 9662 172046 9758 172102
rect 9138 171978 9758 172046
rect 9138 171922 9234 171978
rect 9290 171922 9358 171978
rect 9414 171922 9482 171978
rect 9538 171922 9606 171978
rect 9662 171922 9758 171978
rect 9138 154350 9758 171922
rect 36138 166350 36758 183922
rect 55168 184350 55488 184384
rect 55168 184294 55238 184350
rect 55294 184294 55362 184350
rect 55418 184294 55488 184350
rect 55168 184226 55488 184294
rect 55168 184170 55238 184226
rect 55294 184170 55362 184226
rect 55418 184170 55488 184226
rect 55168 184102 55488 184170
rect 55168 184046 55238 184102
rect 55294 184046 55362 184102
rect 55418 184046 55488 184102
rect 55168 183978 55488 184046
rect 55168 183922 55238 183978
rect 55294 183922 55362 183978
rect 55418 183922 55488 183978
rect 55168 183888 55488 183922
rect 66858 184350 67478 201922
rect 66858 184294 66954 184350
rect 67010 184294 67078 184350
rect 67134 184294 67202 184350
rect 67258 184294 67326 184350
rect 67382 184294 67478 184350
rect 66858 184226 67478 184294
rect 66858 184170 66954 184226
rect 67010 184170 67078 184226
rect 67134 184170 67202 184226
rect 67258 184170 67326 184226
rect 67382 184170 67478 184226
rect 66858 184102 67478 184170
rect 66858 184046 66954 184102
rect 67010 184046 67078 184102
rect 67134 184046 67202 184102
rect 67258 184046 67326 184102
rect 67382 184046 67478 184102
rect 66858 183978 67478 184046
rect 66858 183922 66954 183978
rect 67010 183922 67078 183978
rect 67134 183922 67202 183978
rect 67258 183922 67326 183978
rect 67382 183922 67478 183978
rect 36138 166294 36234 166350
rect 36290 166294 36358 166350
rect 36414 166294 36482 166350
rect 36538 166294 36606 166350
rect 36662 166294 36758 166350
rect 36138 166226 36758 166294
rect 36138 166170 36234 166226
rect 36290 166170 36358 166226
rect 36414 166170 36482 166226
rect 36538 166170 36606 166226
rect 36662 166170 36758 166226
rect 36138 166102 36758 166170
rect 36138 166046 36234 166102
rect 36290 166046 36358 166102
rect 36414 166046 36482 166102
rect 36538 166046 36606 166102
rect 36662 166046 36758 166102
rect 36138 165978 36758 166046
rect 36138 165922 36234 165978
rect 36290 165922 36358 165978
rect 36414 165922 36482 165978
rect 36538 165922 36606 165978
rect 36662 165922 36758 165978
rect 9138 154294 9234 154350
rect 9290 154294 9358 154350
rect 9414 154294 9482 154350
rect 9538 154294 9606 154350
rect 9662 154294 9758 154350
rect 9138 154226 9758 154294
rect 9138 154170 9234 154226
rect 9290 154170 9358 154226
rect 9414 154170 9482 154226
rect 9538 154170 9606 154226
rect 9662 154170 9758 154226
rect 9138 154102 9758 154170
rect 9138 154046 9234 154102
rect 9290 154046 9358 154102
rect 9414 154046 9482 154102
rect 9538 154046 9606 154102
rect 9662 154046 9758 154102
rect 9138 153978 9758 154046
rect 9138 153922 9234 153978
rect 9290 153922 9358 153978
rect 9414 153922 9482 153978
rect 9538 153922 9606 153978
rect 9662 153922 9758 153978
rect 9138 136350 9758 153922
rect 9138 136294 9234 136350
rect 9290 136294 9358 136350
rect 9414 136294 9482 136350
rect 9538 136294 9606 136350
rect 9662 136294 9758 136350
rect 9138 136226 9758 136294
rect 9138 136170 9234 136226
rect 9290 136170 9358 136226
rect 9414 136170 9482 136226
rect 9538 136170 9606 136226
rect 9662 136170 9758 136226
rect 9138 136102 9758 136170
rect 9138 136046 9234 136102
rect 9290 136046 9358 136102
rect 9414 136046 9482 136102
rect 9538 136046 9606 136102
rect 9662 136046 9758 136102
rect 9138 135978 9758 136046
rect 9138 135922 9234 135978
rect 9290 135922 9358 135978
rect 9414 135922 9482 135978
rect 9538 135922 9606 135978
rect 9662 135922 9758 135978
rect 9138 118350 9758 135922
rect 18172 156436 18228 156446
rect 18172 121268 18228 156380
rect 36138 148350 36758 165922
rect 36138 148294 36234 148350
rect 36290 148294 36358 148350
rect 36414 148294 36482 148350
rect 36538 148294 36606 148350
rect 36662 148294 36758 148350
rect 36138 148226 36758 148294
rect 36138 148170 36234 148226
rect 36290 148170 36358 148226
rect 36414 148170 36482 148226
rect 36538 148170 36606 148226
rect 36662 148170 36758 148226
rect 36138 148102 36758 148170
rect 36138 148046 36234 148102
rect 36290 148046 36358 148102
rect 36414 148046 36482 148102
rect 36538 148046 36606 148102
rect 36662 148046 36758 148102
rect 36138 147978 36758 148046
rect 36138 147922 36234 147978
rect 36290 147922 36358 147978
rect 36414 147922 36482 147978
rect 36538 147922 36606 147978
rect 36662 147922 36758 147978
rect 20076 131338 20132 131348
rect 19964 131282 20076 131338
rect 18396 131158 18452 131168
rect 18284 128638 18340 128648
rect 18284 126028 18340 128582
rect 18396 127316 18452 131102
rect 18396 127250 18452 127260
rect 19964 126028 20020 131282
rect 20076 131272 20132 131282
rect 24448 130350 24768 130384
rect 24448 130294 24518 130350
rect 24574 130294 24642 130350
rect 24698 130294 24768 130350
rect 24448 130226 24768 130294
rect 24448 130170 24518 130226
rect 24574 130170 24642 130226
rect 24698 130170 24768 130226
rect 24448 130102 24768 130170
rect 24448 130046 24518 130102
rect 24574 130046 24642 130102
rect 24698 130046 24768 130102
rect 24448 129978 24768 130046
rect 24448 129922 24518 129978
rect 24574 129922 24642 129978
rect 24698 129922 24768 129978
rect 24448 129888 24768 129922
rect 36138 130350 36758 147922
rect 39858 172350 40478 172564
rect 39858 172294 39954 172350
rect 40010 172294 40078 172350
rect 40134 172294 40202 172350
rect 40258 172294 40326 172350
rect 40382 172294 40478 172350
rect 39858 172226 40478 172294
rect 39858 172170 39954 172226
rect 40010 172170 40078 172226
rect 40134 172170 40202 172226
rect 40258 172170 40326 172226
rect 40382 172170 40478 172226
rect 39858 172102 40478 172170
rect 39858 172046 39954 172102
rect 40010 172046 40078 172102
rect 40134 172046 40202 172102
rect 40258 172046 40326 172102
rect 40382 172046 40478 172102
rect 39858 171978 40478 172046
rect 39858 171922 39954 171978
rect 40010 171922 40078 171978
rect 40134 171922 40202 171978
rect 40258 171922 40326 171978
rect 40382 171922 40478 171978
rect 39858 154350 40478 171922
rect 66858 166350 67478 183922
rect 66858 166294 66954 166350
rect 67010 166294 67078 166350
rect 67134 166294 67202 166350
rect 67258 166294 67326 166350
rect 67382 166294 67478 166350
rect 66858 166226 67478 166294
rect 66858 166170 66954 166226
rect 67010 166170 67078 166226
rect 67134 166170 67202 166226
rect 67258 166170 67326 166226
rect 67382 166170 67478 166226
rect 66858 166102 67478 166170
rect 66858 166046 66954 166102
rect 67010 166046 67078 166102
rect 67134 166046 67202 166102
rect 67258 166046 67326 166102
rect 67382 166046 67478 166102
rect 66858 165978 67478 166046
rect 66858 165922 66954 165978
rect 67010 165922 67078 165978
rect 67134 165922 67202 165978
rect 67258 165922 67326 165978
rect 67382 165922 67478 165978
rect 64876 158676 64932 158686
rect 64764 156996 64820 157006
rect 39858 154294 39954 154350
rect 40010 154294 40078 154350
rect 40134 154294 40202 154350
rect 40258 154294 40326 154350
rect 40382 154294 40478 154350
rect 39858 154226 40478 154294
rect 39858 154170 39954 154226
rect 40010 154170 40078 154226
rect 40134 154170 40202 154226
rect 40258 154170 40326 154226
rect 40382 154170 40478 154226
rect 39858 154102 40478 154170
rect 39858 154046 39954 154102
rect 40010 154046 40078 154102
rect 40134 154046 40202 154102
rect 40258 154046 40326 154102
rect 40382 154046 40478 154102
rect 39858 153978 40478 154046
rect 39858 153922 39954 153978
rect 40010 153922 40078 153978
rect 40134 153922 40202 153978
rect 40258 153922 40326 153978
rect 40382 153922 40478 153978
rect 39858 140988 40478 153922
rect 64652 154756 64708 154766
rect 39808 136350 40128 136384
rect 39808 136294 39878 136350
rect 39934 136294 40002 136350
rect 40058 136294 40128 136350
rect 39808 136226 40128 136294
rect 39808 136170 39878 136226
rect 39934 136170 40002 136226
rect 40058 136170 40128 136226
rect 39808 136102 40128 136170
rect 39808 136046 39878 136102
rect 39934 136046 40002 136102
rect 40058 136046 40128 136102
rect 39808 135978 40128 136046
rect 39808 135922 39878 135978
rect 39934 135922 40002 135978
rect 40058 135922 40128 135978
rect 39808 135888 40128 135922
rect 36138 130294 36234 130350
rect 36290 130294 36358 130350
rect 36414 130294 36482 130350
rect 36538 130294 36606 130350
rect 36662 130294 36758 130350
rect 36138 130226 36758 130294
rect 36138 130170 36234 130226
rect 36290 130170 36358 130226
rect 36414 130170 36482 130226
rect 36538 130170 36606 130226
rect 36662 130170 36758 130226
rect 36138 130102 36758 130170
rect 36138 130046 36234 130102
rect 36290 130046 36358 130102
rect 36414 130046 36482 130102
rect 36538 130046 36606 130102
rect 36662 130046 36758 130102
rect 36138 129978 36758 130046
rect 36138 129922 36234 129978
rect 36290 129922 36358 129978
rect 36414 129922 36482 129978
rect 36538 129922 36606 129978
rect 36662 129922 36758 129978
rect 36138 129486 36758 129922
rect 55168 130350 55488 130384
rect 55168 130294 55238 130350
rect 55294 130294 55362 130350
rect 55418 130294 55488 130350
rect 55168 130226 55488 130294
rect 55168 130170 55238 130226
rect 55294 130170 55362 130226
rect 55418 130170 55488 130226
rect 55168 130102 55488 130170
rect 55168 130046 55238 130102
rect 55294 130046 55362 130102
rect 55418 130046 55488 130102
rect 55168 129978 55488 130046
rect 55168 129922 55238 129978
rect 55294 129922 55362 129978
rect 55418 129922 55488 129978
rect 55168 129888 55488 129922
rect 20076 127988 20132 127998
rect 20076 127918 20132 127932
rect 20076 127852 20132 127862
rect 37772 127918 37828 127928
rect 20636 127558 20692 127568
rect 20636 127204 20692 127502
rect 37772 127558 37828 127862
rect 37772 127492 37828 127502
rect 20636 127138 20692 127148
rect 18284 125972 18452 126028
rect 19964 125972 20132 126028
rect 18172 121202 18228 121212
rect 18396 119252 18452 125972
rect 18396 119186 18452 119196
rect 20076 118580 20132 125972
rect 64204 124318 64260 124328
rect 64204 123284 64260 124262
rect 64204 123218 64260 123228
rect 64204 120898 64260 120908
rect 64204 119924 64260 120842
rect 64204 119858 64260 119868
rect 20076 118514 20132 118524
rect 9138 118294 9234 118350
rect 9290 118294 9358 118350
rect 9414 118294 9482 118350
rect 9538 118294 9606 118350
rect 9662 118294 9758 118350
rect 9138 118226 9758 118294
rect 9138 118170 9234 118226
rect 9290 118170 9358 118226
rect 9414 118170 9482 118226
rect 9538 118170 9606 118226
rect 9662 118170 9758 118226
rect 9138 118102 9758 118170
rect 9138 118046 9234 118102
rect 9290 118046 9358 118102
rect 9414 118046 9482 118102
rect 9538 118046 9606 118102
rect 9662 118046 9758 118102
rect 9138 117978 9758 118046
rect 9138 117922 9234 117978
rect 9290 117922 9358 117978
rect 9414 117922 9482 117978
rect 9538 117922 9606 117978
rect 9662 117922 9758 117978
rect 9138 100350 9758 117922
rect 39808 118350 40128 118384
rect 39808 118294 39878 118350
rect 39934 118294 40002 118350
rect 40058 118294 40128 118350
rect 39808 118226 40128 118294
rect 39808 118170 39878 118226
rect 39934 118170 40002 118226
rect 40058 118170 40128 118226
rect 39808 118102 40128 118170
rect 39808 118046 39878 118102
rect 39934 118046 40002 118102
rect 40058 118046 40128 118102
rect 39808 117978 40128 118046
rect 39808 117922 39878 117978
rect 39934 117922 40002 117978
rect 40058 117922 40128 117978
rect 39808 117888 40128 117922
rect 64652 117908 64708 154700
rect 64764 121940 64820 156940
rect 64876 126644 64932 158620
rect 64876 126578 64932 126588
rect 64988 157556 65044 157566
rect 64764 121874 64820 121884
rect 64988 121268 65044 157500
rect 64988 121202 65044 121212
rect 66858 148350 67478 165922
rect 66858 148294 66954 148350
rect 67010 148294 67078 148350
rect 67134 148294 67202 148350
rect 67258 148294 67326 148350
rect 67382 148294 67478 148350
rect 66858 148226 67478 148294
rect 66858 148170 66954 148226
rect 67010 148170 67078 148226
rect 67134 148170 67202 148226
rect 67258 148170 67326 148226
rect 67382 148170 67478 148226
rect 66858 148102 67478 148170
rect 66858 148046 66954 148102
rect 67010 148046 67078 148102
rect 67134 148046 67202 148102
rect 67258 148046 67326 148102
rect 67382 148046 67478 148102
rect 66858 147978 67478 148046
rect 66858 147922 66954 147978
rect 67010 147922 67078 147978
rect 67134 147922 67202 147978
rect 67258 147922 67326 147978
rect 67382 147922 67478 147978
rect 66858 130350 67478 147922
rect 70578 226350 71198 243922
rect 81452 242676 81508 261212
rect 82012 260372 82068 281484
rect 86448 274350 86768 274384
rect 86448 274294 86518 274350
rect 86574 274294 86642 274350
rect 86698 274294 86768 274350
rect 86448 274226 86768 274294
rect 86448 274170 86518 274226
rect 86574 274170 86642 274226
rect 86698 274170 86768 274226
rect 86448 274102 86768 274170
rect 86448 274046 86518 274102
rect 86574 274046 86642 274102
rect 86698 274046 86768 274102
rect 86448 273978 86768 274046
rect 86448 273922 86518 273978
rect 86574 273922 86642 273978
rect 86698 273922 86768 273978
rect 86448 273888 86768 273922
rect 97578 274350 98198 291922
rect 128298 310350 128918 327922
rect 128298 310294 128394 310350
rect 128450 310294 128518 310350
rect 128574 310294 128642 310350
rect 128698 310294 128766 310350
rect 128822 310294 128918 310350
rect 128298 310226 128918 310294
rect 128298 310170 128394 310226
rect 128450 310170 128518 310226
rect 128574 310170 128642 310226
rect 128698 310170 128766 310226
rect 128822 310170 128918 310226
rect 128298 310102 128918 310170
rect 128298 310046 128394 310102
rect 128450 310046 128518 310102
rect 128574 310046 128642 310102
rect 128698 310046 128766 310102
rect 128822 310046 128918 310102
rect 128298 309978 128918 310046
rect 128298 309922 128394 309978
rect 128450 309922 128518 309978
rect 128574 309922 128642 309978
rect 128698 309922 128766 309978
rect 128822 309922 128918 309978
rect 128298 292350 128918 309922
rect 128298 292294 128394 292350
rect 128450 292294 128518 292350
rect 128574 292294 128642 292350
rect 128698 292294 128766 292350
rect 128822 292294 128918 292350
rect 128298 292226 128918 292294
rect 128298 292170 128394 292226
rect 128450 292170 128518 292226
rect 128574 292170 128642 292226
rect 128698 292170 128766 292226
rect 128822 292170 128918 292226
rect 128298 292102 128918 292170
rect 128298 292046 128394 292102
rect 128450 292046 128518 292102
rect 128574 292046 128642 292102
rect 128698 292046 128766 292102
rect 128822 292046 128918 292102
rect 128298 291978 128918 292046
rect 128298 291922 128394 291978
rect 128450 291922 128518 291978
rect 128574 291922 128642 291978
rect 128698 291922 128766 291978
rect 128822 291922 128918 291978
rect 101808 280350 102128 280384
rect 101808 280294 101878 280350
rect 101934 280294 102002 280350
rect 102058 280294 102128 280350
rect 101808 280226 102128 280294
rect 101808 280170 101878 280226
rect 101934 280170 102002 280226
rect 102058 280170 102128 280226
rect 101808 280102 102128 280170
rect 101808 280046 101878 280102
rect 101934 280046 102002 280102
rect 102058 280046 102128 280102
rect 101808 279978 102128 280046
rect 101808 279922 101878 279978
rect 101934 279922 102002 279978
rect 102058 279922 102128 279978
rect 101808 279888 102128 279922
rect 126812 278038 126868 278048
rect 124348 275698 124404 275708
rect 97578 274294 97674 274350
rect 97730 274294 97798 274350
rect 97854 274294 97922 274350
rect 97978 274294 98046 274350
rect 98102 274294 98198 274350
rect 97578 274226 98198 274294
rect 97578 274170 97674 274226
rect 97730 274170 97798 274226
rect 97854 274170 97922 274226
rect 97978 274170 98046 274226
rect 98102 274170 98198 274226
rect 97578 274102 98198 274170
rect 97578 274046 97674 274102
rect 97730 274046 97798 274102
rect 97854 274046 97922 274102
rect 97978 274046 98046 274102
rect 98102 274046 98198 274102
rect 97578 273978 98198 274046
rect 97578 273922 97674 273978
rect 97730 273922 97798 273978
rect 97854 273922 97922 273978
rect 97978 273922 98046 273978
rect 98102 273922 98198 273978
rect 82460 270658 82516 270668
rect 82460 270452 82516 270602
rect 82460 270386 82516 270396
rect 82460 267058 82516 267068
rect 82460 266980 82516 267002
rect 82460 266914 82516 266924
rect 82012 260306 82068 260316
rect 82684 262388 82740 262398
rect 82684 259498 82740 262332
rect 82684 259432 82740 259442
rect 81564 258356 81620 258366
rect 81564 244356 81620 258300
rect 86448 256350 86768 256384
rect 86448 256294 86518 256350
rect 86574 256294 86642 256350
rect 86698 256294 86768 256350
rect 86448 256226 86768 256294
rect 86448 256170 86518 256226
rect 86574 256170 86642 256226
rect 86698 256170 86768 256226
rect 86448 256102 86768 256170
rect 86448 256046 86518 256102
rect 86574 256046 86642 256102
rect 86698 256046 86768 256102
rect 86448 255978 86768 256046
rect 86448 255922 86518 255978
rect 86574 255922 86642 255978
rect 86698 255922 86768 255978
rect 86448 255888 86768 255922
rect 97578 256350 98198 273922
rect 117168 274350 117488 274384
rect 117168 274294 117238 274350
rect 117294 274294 117362 274350
rect 117418 274294 117488 274350
rect 117168 274226 117488 274294
rect 117168 274170 117238 274226
rect 117294 274170 117362 274226
rect 117418 274170 117488 274226
rect 117168 274102 117488 274170
rect 117168 274046 117238 274102
rect 117294 274046 117362 274102
rect 117418 274046 117488 274102
rect 117168 273978 117488 274046
rect 117168 273922 117238 273978
rect 117294 273922 117362 273978
rect 117418 273922 117488 273978
rect 117168 273888 117488 273922
rect 124348 268498 124404 275642
rect 124348 268432 124404 268442
rect 126812 265748 126868 277982
rect 127596 276418 127652 276428
rect 127484 276362 127596 276418
rect 127484 269108 127540 276362
rect 127596 276352 127652 276362
rect 128298 274350 128918 291922
rect 132018 334350 132638 351922
rect 159018 364102 159638 364170
rect 159018 364046 159114 364102
rect 159170 364046 159238 364102
rect 159294 364046 159362 364102
rect 159418 364046 159486 364102
rect 159542 364046 159638 364102
rect 159018 363978 159638 364046
rect 159018 363922 159114 363978
rect 159170 363922 159238 363978
rect 159294 363922 159362 363978
rect 159418 363922 159486 363978
rect 159542 363922 159638 363978
rect 148448 346350 148768 346384
rect 148448 346294 148518 346350
rect 148574 346294 148642 346350
rect 148698 346294 148768 346350
rect 148448 346226 148768 346294
rect 148448 346170 148518 346226
rect 148574 346170 148642 346226
rect 148698 346170 148768 346226
rect 148448 346102 148768 346170
rect 148448 346046 148518 346102
rect 148574 346046 148642 346102
rect 148698 346046 148768 346102
rect 148448 345978 148768 346046
rect 148448 345922 148518 345978
rect 148574 345922 148642 345978
rect 148698 345922 148768 345978
rect 148448 345888 148768 345922
rect 159018 346350 159638 363922
rect 159018 346294 159114 346350
rect 159170 346294 159238 346350
rect 159294 346294 159362 346350
rect 159418 346294 159486 346350
rect 159542 346294 159638 346350
rect 159018 346226 159638 346294
rect 159018 346170 159114 346226
rect 159170 346170 159238 346226
rect 159294 346170 159362 346226
rect 159418 346170 159486 346226
rect 159542 346170 159638 346226
rect 159018 346102 159638 346170
rect 159018 346046 159114 346102
rect 159170 346046 159238 346102
rect 159294 346046 159362 346102
rect 159418 346046 159486 346102
rect 159542 346046 159638 346102
rect 159018 345978 159638 346046
rect 159018 345922 159114 345978
rect 159170 345922 159238 345978
rect 159294 345922 159362 345978
rect 159418 345922 159486 345978
rect 159542 345922 159638 345978
rect 141036 341684 141092 341694
rect 141036 341218 141092 341628
rect 144060 341684 144116 341694
rect 144060 341578 144116 341628
rect 144060 341512 144116 341522
rect 141036 341152 141092 341162
rect 141036 340340 141092 340350
rect 132018 334294 132114 334350
rect 132170 334294 132238 334350
rect 132294 334294 132362 334350
rect 132418 334294 132486 334350
rect 132542 334294 132638 334350
rect 132018 334226 132638 334294
rect 132018 334170 132114 334226
rect 132170 334170 132238 334226
rect 132294 334170 132362 334226
rect 132418 334170 132486 334226
rect 132542 334170 132638 334226
rect 132018 334102 132638 334170
rect 132018 334046 132114 334102
rect 132170 334046 132238 334102
rect 132294 334046 132362 334102
rect 132418 334046 132486 334102
rect 132542 334046 132638 334102
rect 132018 333978 132638 334046
rect 132018 333922 132114 333978
rect 132170 333922 132238 333978
rect 132294 333922 132362 333978
rect 132418 333922 132486 333978
rect 132542 333922 132638 333978
rect 132018 316350 132638 333922
rect 140924 337652 140980 337662
rect 140924 319172 140980 337596
rect 140924 319106 140980 319116
rect 132018 316294 132114 316350
rect 132170 316294 132238 316350
rect 132294 316294 132362 316350
rect 132418 316294 132486 316350
rect 132542 316294 132638 316350
rect 132018 316226 132638 316294
rect 132018 316170 132114 316226
rect 132170 316170 132238 316226
rect 132294 316170 132362 316226
rect 132418 316170 132486 316226
rect 132542 316170 132638 316226
rect 132018 316102 132638 316170
rect 132018 316046 132114 316102
rect 132170 316046 132238 316102
rect 132294 316046 132362 316102
rect 132418 316046 132486 316102
rect 132542 316046 132638 316102
rect 132018 315978 132638 316046
rect 132018 315922 132114 315978
rect 132170 315922 132238 315978
rect 132294 315922 132362 315978
rect 132418 315922 132486 315978
rect 132542 315922 132638 315978
rect 132018 298350 132638 315922
rect 141036 314356 141092 340284
rect 143612 338548 143668 338558
rect 141036 314290 141092 314300
rect 141932 337428 141988 337438
rect 141932 307636 141988 337372
rect 142828 319172 142884 319182
rect 142828 316596 142884 319116
rect 142828 316530 142884 316540
rect 143612 310436 143668 338492
rect 148448 328350 148768 328384
rect 148448 328294 148518 328350
rect 148574 328294 148642 328350
rect 148698 328294 148768 328350
rect 148448 328226 148768 328294
rect 148448 328170 148518 328226
rect 148574 328170 148642 328226
rect 148698 328170 148768 328226
rect 148448 328102 148768 328170
rect 148448 328046 148518 328102
rect 148574 328046 148642 328102
rect 148698 328046 148768 328102
rect 148448 327978 148768 328046
rect 148448 327922 148518 327978
rect 148574 327922 148642 327978
rect 148698 327922 148768 327978
rect 148448 327888 148768 327922
rect 159018 328350 159638 345922
rect 162738 442350 163358 459922
rect 163808 460350 164128 460384
rect 163808 460294 163878 460350
rect 163934 460294 164002 460350
rect 164058 460294 164128 460350
rect 163808 460226 164128 460294
rect 163808 460170 163878 460226
rect 163934 460170 164002 460226
rect 164058 460170 164128 460226
rect 163808 460102 164128 460170
rect 163808 460046 163878 460102
rect 163934 460046 164002 460102
rect 164058 460046 164128 460102
rect 163808 459978 164128 460046
rect 163808 459922 163878 459978
rect 163934 459922 164002 459978
rect 164058 459922 164128 459978
rect 163808 459888 164128 459922
rect 162738 442294 162834 442350
rect 162890 442294 162958 442350
rect 163014 442294 163082 442350
rect 163138 442294 163206 442350
rect 163262 442294 163358 442350
rect 162738 442226 163358 442294
rect 162738 442170 162834 442226
rect 162890 442170 162958 442226
rect 163014 442170 163082 442226
rect 163138 442170 163206 442226
rect 163262 442170 163358 442226
rect 162738 442102 163358 442170
rect 162738 442046 162834 442102
rect 162890 442046 162958 442102
rect 163014 442046 163082 442102
rect 163138 442046 163206 442102
rect 163262 442046 163358 442102
rect 162738 441978 163358 442046
rect 162738 441922 162834 441978
rect 162890 441922 162958 441978
rect 163014 441922 163082 441978
rect 163138 441922 163206 441978
rect 163262 441922 163358 441978
rect 162738 424350 163358 441922
rect 189738 454350 190358 471922
rect 193458 598172 194078 598268
rect 193458 598116 193554 598172
rect 193610 598116 193678 598172
rect 193734 598116 193802 598172
rect 193858 598116 193926 598172
rect 193982 598116 194078 598172
rect 193458 598048 194078 598116
rect 193458 597992 193554 598048
rect 193610 597992 193678 598048
rect 193734 597992 193802 598048
rect 193858 597992 193926 598048
rect 193982 597992 194078 598048
rect 193458 597924 194078 597992
rect 193458 597868 193554 597924
rect 193610 597868 193678 597924
rect 193734 597868 193802 597924
rect 193858 597868 193926 597924
rect 193982 597868 194078 597924
rect 193458 597800 194078 597868
rect 193458 597744 193554 597800
rect 193610 597744 193678 597800
rect 193734 597744 193802 597800
rect 193858 597744 193926 597800
rect 193982 597744 194078 597800
rect 193458 586350 194078 597744
rect 193458 586294 193554 586350
rect 193610 586294 193678 586350
rect 193734 586294 193802 586350
rect 193858 586294 193926 586350
rect 193982 586294 194078 586350
rect 193458 586226 194078 586294
rect 193458 586170 193554 586226
rect 193610 586170 193678 586226
rect 193734 586170 193802 586226
rect 193858 586170 193926 586226
rect 193982 586170 194078 586226
rect 193458 586102 194078 586170
rect 193458 586046 193554 586102
rect 193610 586046 193678 586102
rect 193734 586046 193802 586102
rect 193858 586046 193926 586102
rect 193982 586046 194078 586102
rect 193458 585978 194078 586046
rect 193458 585922 193554 585978
rect 193610 585922 193678 585978
rect 193734 585922 193802 585978
rect 193858 585922 193926 585978
rect 193982 585922 194078 585978
rect 193458 568350 194078 585922
rect 220458 597212 221078 598268
rect 220458 597156 220554 597212
rect 220610 597156 220678 597212
rect 220734 597156 220802 597212
rect 220858 597156 220926 597212
rect 220982 597156 221078 597212
rect 220458 597088 221078 597156
rect 220458 597032 220554 597088
rect 220610 597032 220678 597088
rect 220734 597032 220802 597088
rect 220858 597032 220926 597088
rect 220982 597032 221078 597088
rect 220458 596964 221078 597032
rect 220458 596908 220554 596964
rect 220610 596908 220678 596964
rect 220734 596908 220802 596964
rect 220858 596908 220926 596964
rect 220982 596908 221078 596964
rect 220458 596840 221078 596908
rect 220458 596784 220554 596840
rect 220610 596784 220678 596840
rect 220734 596784 220802 596840
rect 220858 596784 220926 596840
rect 220982 596784 221078 596840
rect 220458 580350 221078 596784
rect 220458 580294 220554 580350
rect 220610 580294 220678 580350
rect 220734 580294 220802 580350
rect 220858 580294 220926 580350
rect 220982 580294 221078 580350
rect 220458 580226 221078 580294
rect 220458 580170 220554 580226
rect 220610 580170 220678 580226
rect 220734 580170 220802 580226
rect 220858 580170 220926 580226
rect 220982 580170 221078 580226
rect 220458 580102 221078 580170
rect 220458 580046 220554 580102
rect 220610 580046 220678 580102
rect 220734 580046 220802 580102
rect 220858 580046 220926 580102
rect 220982 580046 221078 580102
rect 220458 579978 221078 580046
rect 220458 579922 220554 579978
rect 220610 579922 220678 579978
rect 220734 579922 220802 579978
rect 220858 579922 220926 579978
rect 220982 579922 221078 579978
rect 193458 568294 193554 568350
rect 193610 568294 193678 568350
rect 193734 568294 193802 568350
rect 193858 568294 193926 568350
rect 193982 568294 194078 568350
rect 193458 568226 194078 568294
rect 193458 568170 193554 568226
rect 193610 568170 193678 568226
rect 193734 568170 193802 568226
rect 193858 568170 193926 568226
rect 193982 568170 194078 568226
rect 193458 568102 194078 568170
rect 193458 568046 193554 568102
rect 193610 568046 193678 568102
rect 193734 568046 193802 568102
rect 193858 568046 193926 568102
rect 193982 568046 194078 568102
rect 193458 567978 194078 568046
rect 193458 567922 193554 567978
rect 193610 567922 193678 567978
rect 193734 567922 193802 567978
rect 193858 567922 193926 567978
rect 193982 567922 194078 567978
rect 193458 550350 194078 567922
rect 193458 550294 193554 550350
rect 193610 550294 193678 550350
rect 193734 550294 193802 550350
rect 193858 550294 193926 550350
rect 193982 550294 194078 550350
rect 193458 550226 194078 550294
rect 193458 550170 193554 550226
rect 193610 550170 193678 550226
rect 193734 550170 193802 550226
rect 193858 550170 193926 550226
rect 193982 550170 194078 550226
rect 193458 550102 194078 550170
rect 193458 550046 193554 550102
rect 193610 550046 193678 550102
rect 193734 550046 193802 550102
rect 193858 550046 193926 550102
rect 193982 550046 194078 550102
rect 193458 549978 194078 550046
rect 193458 549922 193554 549978
rect 193610 549922 193678 549978
rect 193734 549922 193802 549978
rect 193858 549922 193926 549978
rect 193982 549922 194078 549978
rect 193458 532350 194078 549922
rect 200844 571258 200900 571268
rect 193458 532294 193554 532350
rect 193610 532294 193678 532350
rect 193734 532294 193802 532350
rect 193858 532294 193926 532350
rect 193982 532294 194078 532350
rect 193458 532226 194078 532294
rect 193458 532170 193554 532226
rect 193610 532170 193678 532226
rect 193734 532170 193802 532226
rect 193858 532170 193926 532226
rect 193982 532170 194078 532226
rect 193458 532102 194078 532170
rect 193458 532046 193554 532102
rect 193610 532046 193678 532102
rect 193734 532046 193802 532102
rect 193858 532046 193926 532102
rect 193982 532046 194078 532102
rect 193458 531978 194078 532046
rect 193458 531922 193554 531978
rect 193610 531922 193678 531978
rect 193734 531922 193802 531978
rect 193858 531922 193926 531978
rect 193982 531922 194078 531978
rect 193458 514350 194078 531922
rect 197372 545860 197428 545870
rect 197372 522676 197428 545804
rect 197372 522610 197428 522620
rect 193458 514294 193554 514350
rect 193610 514294 193678 514350
rect 193734 514294 193802 514350
rect 193858 514294 193926 514350
rect 193982 514294 194078 514350
rect 193458 514226 194078 514294
rect 193458 514170 193554 514226
rect 193610 514170 193678 514226
rect 193734 514170 193802 514226
rect 193858 514170 193926 514226
rect 193982 514170 194078 514226
rect 193458 514102 194078 514170
rect 193458 514046 193554 514102
rect 193610 514046 193678 514102
rect 193734 514046 193802 514102
rect 193858 514046 193926 514102
rect 193982 514046 194078 514102
rect 193458 513978 194078 514046
rect 193458 513922 193554 513978
rect 193610 513922 193678 513978
rect 193734 513922 193802 513978
rect 193858 513922 193926 513978
rect 193982 513922 194078 513978
rect 193458 496350 194078 513922
rect 193458 496294 193554 496350
rect 193610 496294 193678 496350
rect 193734 496294 193802 496350
rect 193858 496294 193926 496350
rect 193982 496294 194078 496350
rect 193458 496226 194078 496294
rect 193458 496170 193554 496226
rect 193610 496170 193678 496226
rect 193734 496170 193802 496226
rect 193858 496170 193926 496226
rect 193982 496170 194078 496226
rect 193458 496102 194078 496170
rect 193458 496046 193554 496102
rect 193610 496046 193678 496102
rect 193734 496046 193802 496102
rect 193858 496046 193926 496102
rect 193982 496046 194078 496102
rect 193458 495978 194078 496046
rect 193458 495922 193554 495978
rect 193610 495922 193678 495978
rect 193734 495922 193802 495978
rect 193858 495922 193926 495978
rect 193982 495922 194078 495978
rect 193458 478350 194078 495922
rect 193458 478294 193554 478350
rect 193610 478294 193678 478350
rect 193734 478294 193802 478350
rect 193858 478294 193926 478350
rect 193982 478294 194078 478350
rect 193458 478226 194078 478294
rect 193458 478170 193554 478226
rect 193610 478170 193678 478226
rect 193734 478170 193802 478226
rect 193858 478170 193926 478226
rect 193982 478170 194078 478226
rect 193458 478102 194078 478170
rect 193458 478046 193554 478102
rect 193610 478046 193678 478102
rect 193734 478046 193802 478102
rect 193858 478046 193926 478102
rect 193982 478046 194078 478102
rect 193458 477978 194078 478046
rect 197372 480004 197428 480014
rect 193458 477922 193554 477978
rect 193610 477922 193678 477978
rect 193734 477922 193802 477978
rect 193858 477922 193926 477978
rect 193982 477922 194078 477978
rect 193116 469558 193172 469568
rect 193116 465238 193172 469502
rect 193116 465172 193172 465182
rect 189738 454294 189834 454350
rect 189890 454294 189958 454350
rect 190014 454294 190082 454350
rect 190138 454294 190206 454350
rect 190262 454294 190358 454350
rect 189738 454226 190358 454294
rect 189738 454170 189834 454226
rect 189890 454170 189958 454226
rect 190014 454170 190082 454226
rect 190138 454170 190206 454226
rect 190262 454170 190358 454226
rect 189738 454102 190358 454170
rect 189738 454046 189834 454102
rect 189890 454046 189958 454102
rect 190014 454046 190082 454102
rect 190138 454046 190206 454102
rect 190262 454046 190358 454102
rect 189738 453978 190358 454046
rect 189738 453922 189834 453978
rect 189890 453922 189958 453978
rect 190014 453922 190082 453978
rect 190138 453922 190206 453978
rect 190262 453922 190358 453978
rect 189738 436350 190358 453922
rect 189738 436294 189834 436350
rect 189890 436294 189958 436350
rect 190014 436294 190082 436350
rect 190138 436294 190206 436350
rect 190262 436294 190358 436350
rect 189738 436226 190358 436294
rect 189738 436170 189834 436226
rect 189890 436170 189958 436226
rect 190014 436170 190082 436226
rect 190138 436170 190206 436226
rect 190262 436170 190358 436226
rect 189738 436102 190358 436170
rect 189738 436046 189834 436102
rect 189890 436046 189958 436102
rect 190014 436046 190082 436102
rect 190138 436046 190206 436102
rect 190262 436046 190358 436102
rect 189738 435978 190358 436046
rect 189738 435922 189834 435978
rect 189890 435922 189958 435978
rect 190014 435922 190082 435978
rect 190138 435922 190206 435978
rect 190262 435922 190358 435978
rect 173852 426692 173908 426702
rect 170268 426468 170324 426478
rect 170268 426132 170324 426412
rect 170268 426066 170324 426076
rect 173740 426356 173796 426366
rect 173740 425908 173796 426300
rect 173852 426132 173908 426636
rect 173852 426066 173908 426076
rect 173740 425842 173796 425852
rect 162738 424294 162834 424350
rect 162890 424294 162958 424350
rect 163014 424294 163082 424350
rect 163138 424294 163206 424350
rect 163262 424294 163358 424350
rect 162738 424226 163358 424294
rect 162738 424170 162834 424226
rect 162890 424170 162958 424226
rect 163014 424170 163082 424226
rect 163138 424170 163206 424226
rect 163262 424170 163358 424226
rect 162738 424102 163358 424170
rect 162738 424046 162834 424102
rect 162890 424046 162958 424102
rect 163014 424046 163082 424102
rect 163138 424046 163206 424102
rect 163262 424046 163358 424102
rect 162738 423978 163358 424046
rect 162738 423922 162834 423978
rect 162890 423922 162958 423978
rect 163014 423922 163082 423978
rect 163138 423922 163206 423978
rect 163262 423922 163358 423978
rect 162738 406350 163358 423922
rect 179168 418350 179488 418384
rect 179168 418294 179238 418350
rect 179294 418294 179362 418350
rect 179418 418294 179488 418350
rect 179168 418226 179488 418294
rect 179168 418170 179238 418226
rect 179294 418170 179362 418226
rect 179418 418170 179488 418226
rect 179168 418102 179488 418170
rect 179168 418046 179238 418102
rect 179294 418046 179362 418102
rect 179418 418046 179488 418102
rect 179168 417978 179488 418046
rect 179168 417922 179238 417978
rect 179294 417922 179362 417978
rect 179418 417922 179488 417978
rect 179168 417888 179488 417922
rect 189738 418350 190358 435922
rect 189738 418294 189834 418350
rect 189890 418294 189958 418350
rect 190014 418294 190082 418350
rect 190138 418294 190206 418350
rect 190262 418294 190358 418350
rect 189738 418226 190358 418294
rect 189738 418170 189834 418226
rect 189890 418170 189958 418226
rect 190014 418170 190082 418226
rect 190138 418170 190206 418226
rect 190262 418170 190358 418226
rect 189738 418102 190358 418170
rect 189738 418046 189834 418102
rect 189890 418046 189958 418102
rect 190014 418046 190082 418102
rect 190138 418046 190206 418102
rect 190262 418046 190358 418102
rect 189738 417978 190358 418046
rect 189738 417922 189834 417978
rect 189890 417922 189958 417978
rect 190014 417922 190082 417978
rect 190138 417922 190206 417978
rect 190262 417922 190358 417978
rect 188972 408100 189028 408110
rect 162738 406294 162834 406350
rect 162890 406294 162958 406350
rect 163014 406294 163082 406350
rect 163138 406294 163206 406350
rect 163262 406294 163358 406350
rect 162738 406226 163358 406294
rect 162738 406170 162834 406226
rect 162890 406170 162958 406226
rect 163014 406170 163082 406226
rect 163138 406170 163206 406226
rect 163262 406170 163358 406226
rect 162738 406102 163358 406170
rect 162738 406046 162834 406102
rect 162890 406046 162958 406102
rect 163014 406046 163082 406102
rect 163138 406046 163206 406102
rect 163262 406046 163358 406102
rect 162738 405978 163358 406046
rect 162738 405922 162834 405978
rect 162890 405922 162958 405978
rect 163014 405922 163082 405978
rect 163138 405922 163206 405978
rect 163262 405922 163358 405978
rect 162738 388350 163358 405922
rect 163808 406350 164128 406384
rect 163808 406294 163878 406350
rect 163934 406294 164002 406350
rect 164058 406294 164128 406350
rect 163808 406226 164128 406294
rect 163808 406170 163878 406226
rect 163934 406170 164002 406226
rect 164058 406170 164128 406226
rect 163808 406102 164128 406170
rect 163808 406046 163878 406102
rect 163934 406046 164002 406102
rect 164058 406046 164128 406102
rect 163808 405978 164128 406046
rect 163808 405922 163878 405978
rect 163934 405922 164002 405978
rect 164058 405922 164128 405978
rect 163808 405888 164128 405922
rect 179168 400350 179488 400384
rect 179168 400294 179238 400350
rect 179294 400294 179362 400350
rect 179418 400294 179488 400350
rect 179168 400226 179488 400294
rect 179168 400170 179238 400226
rect 179294 400170 179362 400226
rect 179418 400170 179488 400226
rect 179168 400102 179488 400170
rect 179168 400046 179238 400102
rect 179294 400046 179362 400102
rect 179418 400046 179488 400102
rect 179168 399978 179488 400046
rect 179168 399922 179238 399978
rect 179294 399922 179362 399978
rect 179418 399922 179488 399978
rect 179168 399888 179488 399922
rect 188972 395668 189028 408044
rect 189308 404758 189364 404768
rect 189308 403396 189364 404702
rect 189420 404740 189476 404750
rect 189420 404038 189476 404684
rect 189532 404578 189588 404588
rect 189532 404068 189588 404522
rect 189532 404002 189588 404012
rect 189420 403972 189476 403982
rect 189308 403330 189364 403340
rect 189532 402052 189588 402062
rect 189532 399538 189588 401996
rect 189532 399472 189588 399482
rect 189738 400350 190358 417922
rect 193458 460350 194078 477922
rect 194908 477988 194964 477998
rect 194908 467938 194964 477932
rect 197372 469558 197428 479948
rect 197372 469492 197428 469502
rect 199052 473284 199108 473294
rect 194908 467872 194964 467882
rect 199052 463618 199108 473228
rect 199052 463552 199108 463562
rect 193458 460294 193554 460350
rect 193610 460294 193678 460350
rect 193734 460294 193802 460350
rect 193858 460294 193926 460350
rect 193982 460294 194078 460350
rect 193458 460226 194078 460294
rect 193458 460170 193554 460226
rect 193610 460170 193678 460226
rect 193734 460170 193802 460226
rect 193858 460170 193926 460226
rect 193982 460170 194078 460226
rect 193458 460102 194078 460170
rect 193458 460046 193554 460102
rect 193610 460046 193678 460102
rect 193734 460046 193802 460102
rect 193858 460046 193926 460102
rect 193982 460046 194078 460102
rect 193458 459978 194078 460046
rect 193458 459922 193554 459978
rect 193610 459922 193678 459978
rect 193734 459922 193802 459978
rect 193858 459922 193926 459978
rect 193982 459922 194078 459978
rect 193458 442350 194078 459922
rect 193458 442294 193554 442350
rect 193610 442294 193678 442350
rect 193734 442294 193802 442350
rect 193858 442294 193926 442350
rect 193982 442294 194078 442350
rect 193458 442226 194078 442294
rect 193458 442170 193554 442226
rect 193610 442170 193678 442226
rect 193734 442170 193802 442226
rect 193858 442170 193926 442226
rect 193982 442170 194078 442226
rect 193458 442102 194078 442170
rect 193458 442046 193554 442102
rect 193610 442046 193678 442102
rect 193734 442046 193802 442102
rect 193858 442046 193926 442102
rect 193982 442046 194078 442102
rect 193458 441978 194078 442046
rect 193458 441922 193554 441978
rect 193610 441922 193678 441978
rect 193734 441922 193802 441978
rect 193858 441922 193926 441978
rect 193982 441922 194078 441978
rect 193458 424350 194078 441922
rect 193458 424294 193554 424350
rect 193610 424294 193678 424350
rect 193734 424294 193802 424350
rect 193858 424294 193926 424350
rect 193982 424294 194078 424350
rect 193458 424226 194078 424294
rect 193458 424170 193554 424226
rect 193610 424170 193678 424226
rect 193734 424170 193802 424226
rect 193858 424170 193926 424226
rect 193982 424170 194078 424226
rect 193458 424102 194078 424170
rect 193458 424046 193554 424102
rect 193610 424046 193678 424102
rect 193734 424046 193802 424102
rect 193858 424046 193926 424102
rect 193982 424046 194078 424102
rect 193458 423978 194078 424046
rect 193458 423922 193554 423978
rect 193610 423922 193678 423978
rect 193734 423922 193802 423978
rect 193858 423922 193926 423978
rect 193982 423922 194078 423978
rect 191548 406918 191604 406928
rect 191548 406084 191604 406862
rect 191548 406018 191604 406028
rect 193458 406350 194078 423922
rect 193458 406294 193554 406350
rect 193610 406294 193678 406350
rect 193734 406294 193802 406350
rect 193858 406294 193926 406350
rect 193982 406294 194078 406350
rect 193458 406226 194078 406294
rect 193458 406170 193554 406226
rect 193610 406170 193678 406226
rect 193734 406170 193802 406226
rect 193858 406170 193926 406226
rect 193982 406170 194078 406226
rect 193458 406102 194078 406170
rect 193458 406046 193554 406102
rect 193610 406046 193678 406102
rect 193734 406046 193802 406102
rect 193858 406046 193926 406102
rect 193982 406046 194078 406102
rect 193458 405978 194078 406046
rect 193458 405922 193554 405978
rect 193610 405922 193678 405978
rect 193734 405922 193802 405978
rect 193858 405922 193926 405978
rect 193982 405922 194078 405978
rect 189738 400294 189834 400350
rect 189890 400294 189958 400350
rect 190014 400294 190082 400350
rect 190138 400294 190206 400350
rect 190262 400294 190358 400350
rect 189738 400226 190358 400294
rect 189738 400170 189834 400226
rect 189890 400170 189958 400226
rect 190014 400170 190082 400226
rect 190138 400170 190206 400226
rect 190262 400170 190358 400226
rect 189738 400102 190358 400170
rect 189738 400046 189834 400102
rect 189890 400046 189958 400102
rect 190014 400046 190082 400102
rect 190138 400046 190206 400102
rect 190262 400046 190358 400102
rect 189738 399978 190358 400046
rect 189738 399922 189834 399978
rect 189890 399922 189958 399978
rect 190014 399922 190082 399978
rect 190138 399922 190206 399978
rect 190262 399922 190358 399978
rect 188972 395602 189028 395612
rect 162738 388294 162834 388350
rect 162890 388294 162958 388350
rect 163014 388294 163082 388350
rect 163138 388294 163206 388350
rect 163262 388294 163358 388350
rect 162738 388226 163358 388294
rect 163808 388389 164128 388446
rect 163808 388333 163836 388389
rect 163892 388333 163940 388389
rect 163996 388333 164044 388389
rect 164100 388333 164128 388389
rect 163808 388276 164128 388333
rect 162738 388170 162834 388226
rect 162890 388170 162958 388226
rect 163014 388170 163082 388226
rect 163138 388170 163206 388226
rect 163262 388170 163358 388226
rect 162738 388102 163358 388170
rect 162738 388046 162834 388102
rect 162890 388046 162958 388102
rect 163014 388046 163082 388102
rect 163138 388046 163206 388102
rect 163262 388046 163358 388102
rect 162738 387978 163358 388046
rect 162738 387922 162834 387978
rect 162890 387922 162958 387978
rect 163014 387922 163082 387978
rect 163138 387922 163206 387978
rect 163262 387922 163358 387978
rect 162738 370350 163358 387922
rect 162738 370294 162834 370350
rect 162890 370294 162958 370350
rect 163014 370294 163082 370350
rect 163138 370294 163206 370350
rect 163262 370294 163358 370350
rect 162738 370226 163358 370294
rect 162738 370170 162834 370226
rect 162890 370170 162958 370226
rect 163014 370170 163082 370226
rect 163138 370170 163206 370226
rect 163262 370170 163358 370226
rect 162738 370102 163358 370170
rect 162738 370046 162834 370102
rect 162890 370046 162958 370102
rect 163014 370046 163082 370102
rect 163138 370046 163206 370102
rect 163262 370046 163358 370102
rect 162738 369978 163358 370046
rect 162738 369922 162834 369978
rect 162890 369922 162958 369978
rect 163014 369922 163082 369978
rect 163138 369922 163206 369978
rect 163262 369922 163358 369978
rect 162738 352350 163358 369922
rect 189738 382350 190358 399922
rect 189738 382294 189834 382350
rect 189890 382294 189958 382350
rect 190014 382294 190082 382350
rect 190138 382294 190206 382350
rect 190262 382294 190358 382350
rect 189738 382226 190358 382294
rect 189738 382170 189834 382226
rect 189890 382170 189958 382226
rect 190014 382170 190082 382226
rect 190138 382170 190206 382226
rect 190262 382170 190358 382226
rect 189738 382102 190358 382170
rect 189738 382046 189834 382102
rect 189890 382046 189958 382102
rect 190014 382046 190082 382102
rect 190138 382046 190206 382102
rect 190262 382046 190358 382102
rect 189738 381978 190358 382046
rect 189738 381922 189834 381978
rect 189890 381922 189958 381978
rect 190014 381922 190082 381978
rect 190138 381922 190206 381978
rect 190262 381922 190358 381978
rect 189738 364350 190358 381922
rect 192332 401380 192388 401390
rect 192332 372036 192388 401324
rect 192332 371970 192388 371980
rect 193458 388350 194078 405922
rect 199836 407428 199892 407438
rect 199836 403138 199892 407372
rect 199836 403072 199892 403082
rect 199052 402418 199108 402428
rect 199052 396298 199108 402362
rect 199052 396232 199108 396242
rect 193458 388294 193554 388350
rect 193610 388294 193678 388350
rect 193734 388294 193802 388350
rect 193858 388294 193926 388350
rect 193982 388294 194078 388350
rect 193458 388226 194078 388294
rect 193458 388170 193554 388226
rect 193610 388170 193678 388226
rect 193734 388170 193802 388226
rect 193858 388170 193926 388226
rect 193982 388170 194078 388226
rect 193458 388102 194078 388170
rect 193458 388046 193554 388102
rect 193610 388046 193678 388102
rect 193734 388046 193802 388102
rect 193858 388046 193926 388102
rect 193982 388046 194078 388102
rect 193458 387978 194078 388046
rect 193458 387922 193554 387978
rect 193610 387922 193678 387978
rect 193734 387922 193802 387978
rect 193858 387922 193926 387978
rect 193982 387922 194078 387978
rect 189738 364294 189834 364350
rect 189890 364294 189958 364350
rect 190014 364294 190082 364350
rect 190138 364294 190206 364350
rect 190262 364294 190358 364350
rect 189738 364226 190358 364294
rect 189738 364170 189834 364226
rect 189890 364170 189958 364226
rect 190014 364170 190082 364226
rect 190138 364170 190206 364226
rect 190262 364170 190358 364226
rect 189738 364102 190358 364170
rect 189738 364046 189834 364102
rect 189890 364046 189958 364102
rect 190014 364046 190082 364102
rect 190138 364046 190206 364102
rect 190262 364046 190358 364102
rect 189738 363978 190358 364046
rect 189738 363922 189834 363978
rect 189890 363922 189958 363978
rect 190014 363922 190082 363978
rect 190138 363922 190206 363978
rect 190262 363922 190358 363978
rect 162738 352294 162834 352350
rect 162890 352294 162958 352350
rect 163014 352294 163082 352350
rect 163138 352294 163206 352350
rect 163262 352294 163358 352350
rect 162738 352226 163358 352294
rect 162738 352170 162834 352226
rect 162890 352170 162958 352226
rect 163014 352170 163082 352226
rect 163138 352170 163206 352226
rect 163262 352170 163358 352226
rect 162738 352102 163358 352170
rect 162738 352046 162834 352102
rect 162890 352046 162958 352102
rect 163014 352046 163082 352102
rect 163138 352046 163206 352102
rect 163262 352046 163358 352102
rect 162738 351978 163358 352046
rect 162738 351922 162834 351978
rect 162890 351922 162958 351978
rect 163014 351922 163082 351978
rect 163138 351922 163206 351978
rect 163262 351922 163358 351978
rect 160524 342838 160580 342848
rect 159740 341578 159796 341588
rect 159740 339238 159796 341522
rect 159740 339172 159796 339182
rect 160524 337618 160580 342782
rect 162738 342190 163358 351922
rect 163808 352350 164128 352384
rect 163808 352294 163878 352350
rect 163934 352294 164002 352350
rect 164058 352294 164128 352350
rect 163808 352226 164128 352294
rect 163808 352170 163878 352226
rect 163934 352170 164002 352226
rect 164058 352170 164128 352226
rect 163808 352102 164128 352170
rect 163808 352046 163878 352102
rect 163934 352046 164002 352102
rect 164058 352046 164128 352102
rect 163808 351978 164128 352046
rect 163808 351922 163878 351978
rect 163934 351922 164002 351978
rect 164058 351922 164128 351978
rect 163808 351888 164128 351922
rect 179168 346350 179488 346384
rect 179168 346294 179238 346350
rect 179294 346294 179362 346350
rect 179418 346294 179488 346350
rect 179168 346226 179488 346294
rect 179168 346170 179238 346226
rect 179294 346170 179362 346226
rect 179418 346170 179488 346226
rect 179168 346102 179488 346170
rect 179168 346046 179238 346102
rect 179294 346046 179362 346102
rect 179418 346046 179488 346102
rect 179168 345978 179488 346046
rect 179168 345922 179238 345978
rect 179294 345922 179362 345978
rect 179418 345922 179488 345978
rect 179168 345888 179488 345922
rect 189738 346350 190358 363922
rect 189738 346294 189834 346350
rect 189890 346294 189958 346350
rect 190014 346294 190082 346350
rect 190138 346294 190206 346350
rect 190262 346294 190358 346350
rect 189738 346226 190358 346294
rect 189738 346170 189834 346226
rect 189890 346170 189958 346226
rect 190014 346170 190082 346226
rect 190138 346170 190206 346226
rect 190262 346170 190358 346226
rect 189738 346102 190358 346170
rect 189738 346046 189834 346102
rect 189890 346046 189958 346102
rect 190014 346046 190082 346102
rect 190138 346046 190206 346102
rect 190262 346046 190358 346102
rect 189738 345978 190358 346046
rect 189738 345922 189834 345978
rect 189890 345922 189958 345978
rect 190014 345922 190082 345978
rect 190138 345922 190206 345978
rect 190262 345922 190358 345978
rect 189084 343558 189140 343568
rect 160524 337552 160580 337562
rect 188972 336980 189028 336990
rect 159018 328294 159114 328350
rect 159170 328294 159238 328350
rect 159294 328294 159362 328350
rect 159418 328294 159486 328350
rect 159542 328294 159638 328350
rect 159018 328226 159638 328294
rect 159018 328170 159114 328226
rect 159170 328170 159238 328226
rect 159294 328170 159362 328226
rect 159418 328170 159486 328226
rect 159542 328170 159638 328226
rect 159018 328102 159638 328170
rect 159018 328046 159114 328102
rect 159170 328046 159238 328102
rect 159294 328046 159362 328102
rect 159418 328046 159486 328102
rect 159542 328046 159638 328102
rect 159018 327978 159638 328046
rect 159018 327922 159114 327978
rect 159170 327922 159238 327978
rect 159294 327922 159362 327978
rect 159418 327922 159486 327978
rect 159542 327922 159638 327978
rect 143612 310370 143668 310380
rect 141932 307570 141988 307580
rect 159018 310350 159638 327922
rect 160412 336178 160468 336188
rect 160412 325918 160468 336122
rect 163808 334350 164128 334384
rect 163808 334294 163878 334350
rect 163934 334294 164002 334350
rect 164058 334294 164128 334350
rect 163808 334226 164128 334294
rect 163808 334170 163878 334226
rect 163934 334170 164002 334226
rect 164058 334170 164128 334226
rect 163808 334102 164128 334170
rect 163808 334046 163878 334102
rect 163934 334046 164002 334102
rect 164058 334046 164128 334102
rect 163808 333978 164128 334046
rect 163808 333922 163878 333978
rect 163934 333922 164002 333978
rect 164058 333922 164128 333978
rect 163808 333888 164128 333922
rect 160412 325852 160468 325862
rect 160524 332758 160580 332768
rect 160524 325738 160580 332702
rect 162540 331858 162596 331868
rect 162540 330598 162596 331802
rect 162540 330532 162596 330542
rect 166236 331138 166292 331148
rect 166236 330418 166292 331082
rect 166236 330352 166292 330362
rect 160524 325672 160580 325682
rect 162738 316350 163358 329602
rect 179168 328350 179488 328384
rect 179168 328294 179238 328350
rect 179294 328294 179362 328350
rect 179418 328294 179488 328350
rect 179168 328226 179488 328294
rect 179168 328170 179238 328226
rect 179294 328170 179362 328226
rect 179418 328170 179488 328226
rect 179168 328102 179488 328170
rect 179168 328046 179238 328102
rect 179294 328046 179362 328102
rect 179418 328046 179488 328102
rect 179168 327978 179488 328046
rect 179168 327922 179238 327978
rect 179294 327922 179362 327978
rect 179418 327922 179488 327978
rect 179168 327888 179488 327922
rect 188972 318388 189028 336924
rect 189084 333620 189140 343502
rect 189532 340340 189588 340350
rect 189532 338548 189588 340284
rect 189084 333554 189140 333564
rect 189420 338518 189476 338528
rect 189532 338482 189588 338492
rect 189420 331604 189476 338462
rect 189420 331538 189476 331548
rect 188972 318322 189028 318332
rect 189738 328350 190358 345922
rect 193458 370350 194078 387922
rect 193458 370294 193554 370350
rect 193610 370294 193678 370350
rect 193734 370294 193802 370350
rect 193858 370294 193926 370350
rect 193982 370294 194078 370350
rect 193458 370226 194078 370294
rect 193458 370170 193554 370226
rect 193610 370170 193678 370226
rect 193734 370170 193802 370226
rect 193858 370170 193926 370226
rect 193982 370170 194078 370226
rect 193458 370102 194078 370170
rect 193458 370046 193554 370102
rect 193610 370046 193678 370102
rect 193734 370046 193802 370102
rect 193858 370046 193926 370102
rect 193982 370046 194078 370102
rect 193458 369978 194078 370046
rect 193458 369922 193554 369978
rect 193610 369922 193678 369978
rect 193734 369922 193802 369978
rect 193858 369922 193926 369978
rect 193982 369922 194078 369978
rect 193458 352350 194078 369922
rect 193458 352294 193554 352350
rect 193610 352294 193678 352350
rect 193734 352294 193802 352350
rect 193858 352294 193926 352350
rect 193982 352294 194078 352350
rect 193458 352226 194078 352294
rect 193458 352170 193554 352226
rect 193610 352170 193678 352226
rect 193734 352170 193802 352226
rect 193858 352170 193926 352226
rect 193982 352170 194078 352226
rect 193458 352102 194078 352170
rect 193458 352046 193554 352102
rect 193610 352046 193678 352102
rect 193734 352046 193802 352102
rect 193858 352046 193926 352102
rect 193982 352046 194078 352102
rect 193458 351978 194078 352046
rect 193458 351922 193554 351978
rect 193610 351922 193678 351978
rect 193734 351922 193802 351978
rect 193858 351922 193926 351978
rect 193982 351922 194078 351978
rect 192444 344458 192500 344468
rect 192332 341758 192388 341768
rect 192332 332948 192388 341702
rect 192444 337652 192500 344402
rect 192444 337586 192500 337596
rect 192332 332882 192388 332892
rect 193458 334350 194078 351922
rect 197372 347878 197428 347888
rect 195692 344638 195748 344648
rect 195692 335636 195748 344582
rect 195804 343018 195860 343028
rect 195804 336308 195860 342962
rect 195804 336242 195860 336252
rect 195692 335570 195748 335580
rect 193458 334294 193554 334350
rect 193610 334294 193678 334350
rect 193734 334294 193802 334350
rect 193858 334294 193926 334350
rect 193982 334294 194078 334350
rect 193458 334226 194078 334294
rect 193458 334170 193554 334226
rect 193610 334170 193678 334226
rect 193734 334170 193802 334226
rect 193858 334170 193926 334226
rect 193982 334170 194078 334226
rect 193458 334102 194078 334170
rect 193458 334046 193554 334102
rect 193610 334046 193678 334102
rect 193734 334046 193802 334102
rect 193858 334046 193926 334102
rect 193982 334046 194078 334102
rect 193458 333978 194078 334046
rect 193458 333922 193554 333978
rect 193610 333922 193678 333978
rect 193734 333922 193802 333978
rect 193858 333922 193926 333978
rect 193982 333922 194078 333978
rect 189738 328294 189834 328350
rect 189890 328294 189958 328350
rect 190014 328294 190082 328350
rect 190138 328294 190206 328350
rect 190262 328294 190358 328350
rect 189738 328226 190358 328294
rect 189738 328170 189834 328226
rect 189890 328170 189958 328226
rect 190014 328170 190082 328226
rect 190138 328170 190206 328226
rect 190262 328170 190358 328226
rect 189738 328102 190358 328170
rect 189738 328046 189834 328102
rect 189890 328046 189958 328102
rect 190014 328046 190082 328102
rect 190138 328046 190206 328102
rect 190262 328046 190358 328102
rect 189738 327978 190358 328046
rect 189738 327922 189834 327978
rect 189890 327922 189958 327978
rect 190014 327922 190082 327978
rect 190138 327922 190206 327978
rect 190262 327922 190358 327978
rect 162738 316294 162834 316350
rect 162890 316294 162958 316350
rect 163014 316294 163082 316350
rect 163138 316294 163206 316350
rect 163262 316294 163358 316350
rect 162738 316226 163358 316294
rect 162738 316170 162834 316226
rect 162890 316170 162958 316226
rect 163014 316170 163082 316226
rect 163138 316170 163206 316226
rect 163262 316170 163358 316226
rect 162738 316102 163358 316170
rect 162738 316046 162834 316102
rect 162890 316046 162958 316102
rect 163014 316046 163082 316102
rect 163138 316046 163206 316102
rect 163262 316046 163358 316102
rect 162738 315978 163358 316046
rect 162738 315922 162834 315978
rect 162890 315922 162958 315978
rect 163014 315922 163082 315978
rect 163138 315922 163206 315978
rect 163262 315922 163358 315978
rect 161308 314692 161364 314702
rect 161308 311556 161364 314636
rect 161308 311490 161364 311500
rect 159018 310294 159114 310350
rect 159170 310294 159238 310350
rect 159294 310294 159362 310350
rect 159418 310294 159486 310350
rect 159542 310294 159638 310350
rect 159018 310226 159638 310294
rect 159018 310170 159114 310226
rect 159170 310170 159238 310226
rect 159294 310170 159362 310226
rect 159418 310170 159486 310226
rect 159542 310170 159638 310226
rect 159018 310102 159638 310170
rect 159018 310046 159114 310102
rect 159170 310046 159238 310102
rect 159294 310046 159362 310102
rect 159418 310046 159486 310102
rect 159542 310046 159638 310102
rect 159018 309978 159638 310046
rect 159018 309922 159114 309978
rect 159170 309922 159238 309978
rect 159294 309922 159362 309978
rect 159418 309922 159486 309978
rect 159542 309922 159638 309978
rect 132018 298294 132114 298350
rect 132170 298294 132238 298350
rect 132294 298294 132362 298350
rect 132418 298294 132486 298350
rect 132542 298294 132638 298350
rect 132018 298226 132638 298294
rect 132018 298170 132114 298226
rect 132170 298170 132238 298226
rect 132294 298170 132362 298226
rect 132418 298170 132486 298226
rect 132542 298170 132638 298226
rect 132018 298102 132638 298170
rect 132018 298046 132114 298102
rect 132170 298046 132238 298102
rect 132294 298046 132362 298102
rect 132418 298046 132486 298102
rect 132542 298046 132638 298102
rect 132018 297978 132638 298046
rect 132018 297922 132114 297978
rect 132170 297922 132238 297978
rect 132294 297922 132362 297978
rect 132418 297922 132486 297978
rect 132542 297922 132638 297978
rect 128298 274294 128394 274350
rect 128450 274294 128518 274350
rect 128574 274294 128642 274350
rect 128698 274294 128766 274350
rect 128822 274294 128918 274350
rect 128298 274226 128918 274294
rect 128298 274170 128394 274226
rect 128450 274170 128518 274226
rect 128574 274170 128642 274226
rect 128698 274170 128766 274226
rect 128822 274170 128918 274226
rect 128298 274102 128918 274170
rect 128298 274046 128394 274102
rect 128450 274046 128518 274102
rect 128574 274046 128642 274102
rect 128698 274046 128766 274102
rect 128822 274046 128918 274102
rect 128298 273978 128918 274046
rect 128298 273922 128394 273978
rect 128450 273922 128518 273978
rect 128574 273922 128642 273978
rect 128698 273922 128766 273978
rect 128822 273922 128918 273978
rect 127596 272998 127652 273008
rect 127596 270452 127652 272942
rect 127596 270386 127652 270396
rect 127484 269042 127540 269052
rect 126812 265682 126868 265692
rect 127596 265076 127652 265086
rect 126812 263732 126868 263742
rect 101808 262350 102128 262384
rect 101808 262294 101878 262350
rect 101934 262294 102002 262350
rect 102058 262294 102128 262350
rect 101808 262226 102128 262294
rect 101808 262170 101878 262226
rect 101934 262170 102002 262226
rect 102058 262170 102128 262226
rect 101808 262102 102128 262170
rect 101808 262046 101878 262102
rect 101934 262046 102002 262102
rect 102058 262046 102128 262102
rect 101808 261978 102128 262046
rect 101808 261922 101878 261978
rect 101934 261922 102002 261978
rect 102058 261922 102128 261978
rect 101808 261888 102128 261922
rect 125132 259498 125188 259508
rect 97578 256294 97674 256350
rect 97730 256294 97798 256350
rect 97854 256294 97922 256350
rect 97978 256294 98046 256350
rect 98102 256294 98198 256350
rect 97578 256226 98198 256294
rect 97578 256170 97674 256226
rect 97730 256170 97798 256226
rect 97854 256170 97922 256226
rect 97978 256170 98046 256226
rect 98102 256170 98198 256226
rect 97578 256102 98198 256170
rect 97578 256046 97674 256102
rect 97730 256046 97798 256102
rect 97854 256046 97922 256102
rect 97978 256046 98046 256102
rect 98102 256046 98198 256102
rect 97578 255978 98198 256046
rect 97578 255922 97674 255978
rect 97730 255922 97798 255978
rect 97854 255922 97922 255978
rect 97978 255922 98046 255978
rect 98102 255922 98198 255978
rect 81564 244290 81620 244300
rect 81452 242610 81508 242620
rect 70578 226294 70674 226350
rect 70730 226294 70798 226350
rect 70854 226294 70922 226350
rect 70978 226294 71046 226350
rect 71102 226294 71198 226350
rect 70578 226226 71198 226294
rect 70578 226170 70674 226226
rect 70730 226170 70798 226226
rect 70854 226170 70922 226226
rect 70978 226170 71046 226226
rect 71102 226170 71198 226226
rect 70578 226102 71198 226170
rect 70578 226046 70674 226102
rect 70730 226046 70798 226102
rect 70854 226046 70922 226102
rect 70978 226046 71046 226102
rect 71102 226046 71198 226102
rect 70578 225978 71198 226046
rect 70578 225922 70674 225978
rect 70730 225922 70798 225978
rect 70854 225922 70922 225978
rect 70978 225922 71046 225978
rect 71102 225922 71198 225978
rect 70578 208350 71198 225922
rect 97578 238350 98198 255922
rect 117168 256350 117488 256384
rect 117168 256294 117238 256350
rect 117294 256294 117362 256350
rect 117418 256294 117488 256350
rect 117168 256226 117488 256294
rect 117168 256170 117238 256226
rect 117294 256170 117362 256226
rect 117418 256170 117488 256226
rect 117168 256102 117488 256170
rect 117168 256046 117238 256102
rect 117294 256046 117362 256102
rect 117418 256046 117488 256102
rect 117168 255978 117488 256046
rect 117168 255922 117238 255978
rect 117294 255922 117362 255978
rect 117418 255922 117488 255978
rect 117168 255888 117488 255922
rect 125132 253378 125188 259442
rect 126812 254458 126868 263676
rect 127596 263060 127652 265020
rect 127596 262994 127652 263004
rect 126812 254392 126868 254402
rect 128298 256350 128918 273922
rect 130284 281652 130340 281662
rect 128298 256294 128394 256350
rect 128450 256294 128518 256350
rect 128574 256294 128642 256350
rect 128698 256294 128766 256350
rect 128822 256294 128918 256350
rect 128298 256226 128918 256294
rect 128298 256170 128394 256226
rect 128450 256170 128518 256226
rect 128574 256170 128642 256226
rect 128698 256170 128766 256226
rect 128822 256170 128918 256226
rect 128298 256102 128918 256170
rect 128298 256046 128394 256102
rect 128450 256046 128518 256102
rect 128574 256046 128642 256102
rect 128698 256046 128766 256102
rect 128822 256046 128918 256102
rect 128298 255978 128918 256046
rect 128298 255922 128394 255978
rect 128450 255922 128518 255978
rect 128574 255922 128642 255978
rect 128698 255922 128766 255978
rect 128822 255922 128918 255978
rect 125132 253312 125188 253322
rect 97578 238294 97674 238350
rect 97730 238294 97798 238350
rect 97854 238294 97922 238350
rect 97978 238294 98046 238350
rect 98102 238294 98198 238350
rect 97578 238226 98198 238294
rect 97578 238170 97674 238226
rect 97730 238170 97798 238226
rect 97854 238170 97922 238226
rect 97978 238170 98046 238226
rect 98102 238170 98198 238226
rect 97578 238102 98198 238170
rect 97578 238046 97674 238102
rect 97730 238046 97798 238102
rect 97854 238046 97922 238102
rect 97978 238046 98046 238102
rect 98102 238046 98198 238102
rect 97578 237978 98198 238046
rect 97578 237922 97674 237978
rect 97730 237922 97798 237978
rect 97854 237922 97922 237978
rect 97978 237922 98046 237978
rect 98102 237922 98198 237978
rect 80332 224756 80388 224766
rect 80108 223076 80164 223086
rect 74732 214676 74788 214686
rect 70578 208294 70674 208350
rect 70730 208294 70798 208350
rect 70854 208294 70922 208350
rect 70978 208294 71046 208350
rect 71102 208294 71198 208350
rect 70578 208226 71198 208294
rect 70578 208170 70674 208226
rect 70730 208170 70798 208226
rect 70854 208170 70922 208226
rect 70978 208170 71046 208226
rect 71102 208170 71198 208226
rect 70578 208102 71198 208170
rect 70578 208046 70674 208102
rect 70730 208046 70798 208102
rect 70854 208046 70922 208102
rect 70978 208046 71046 208102
rect 71102 208046 71198 208102
rect 70578 207978 71198 208046
rect 70578 207922 70674 207978
rect 70730 207922 70798 207978
rect 70854 207922 70922 207978
rect 70978 207922 71046 207978
rect 71102 207922 71198 207978
rect 70578 190350 71198 207922
rect 70578 190294 70674 190350
rect 70730 190294 70798 190350
rect 70854 190294 70922 190350
rect 70978 190294 71046 190350
rect 71102 190294 71198 190350
rect 70578 190226 71198 190294
rect 70578 190170 70674 190226
rect 70730 190170 70798 190226
rect 70854 190170 70922 190226
rect 70978 190170 71046 190226
rect 71102 190170 71198 190226
rect 70578 190102 71198 190170
rect 70578 190046 70674 190102
rect 70730 190046 70798 190102
rect 70854 190046 70922 190102
rect 70978 190046 71046 190102
rect 71102 190046 71198 190102
rect 70578 189978 71198 190046
rect 70578 189922 70674 189978
rect 70730 189922 70798 189978
rect 70854 189922 70922 189978
rect 70978 189922 71046 189978
rect 71102 189922 71198 189978
rect 70578 172350 71198 189922
rect 73052 213332 73108 213342
rect 73052 189812 73108 213276
rect 73052 189746 73108 189756
rect 74732 188468 74788 214620
rect 74844 212100 74900 212110
rect 74844 192500 74900 212044
rect 79996 211652 80052 211662
rect 79996 194516 80052 211596
rect 79996 194450 80052 194460
rect 74844 192434 74900 192444
rect 80108 190484 80164 223020
rect 80220 211204 80276 211214
rect 80220 193844 80276 211148
rect 80332 197876 80388 224700
rect 80332 197810 80388 197820
rect 80444 222516 80500 222526
rect 80444 195188 80500 222460
rect 83132 221396 83188 221406
rect 82012 219268 82068 219278
rect 80444 195122 80500 195132
rect 81452 214228 81508 214238
rect 81452 193956 81508 214172
rect 81676 210756 81732 210766
rect 81676 194628 81732 210700
rect 82012 208348 82068 219212
rect 82236 217588 82292 217598
rect 82012 208292 82180 208348
rect 81676 194562 81732 194572
rect 81452 193890 81508 193900
rect 80220 193778 80276 193788
rect 80108 190418 80164 190428
rect 74732 188402 74788 188412
rect 82124 187796 82180 208292
rect 82124 187730 82180 187740
rect 82236 187124 82292 217532
rect 83132 211652 83188 221340
rect 83132 211586 83188 211596
rect 97578 220350 98198 237922
rect 128298 238350 128918 255922
rect 130172 269780 130228 269790
rect 130172 250318 130228 269724
rect 130284 266420 130340 281596
rect 130284 266354 130340 266364
rect 132018 280350 132638 297922
rect 159018 292350 159638 309922
rect 159018 292294 159114 292350
rect 159170 292294 159238 292350
rect 159294 292294 159362 292350
rect 159418 292294 159486 292350
rect 159542 292294 159638 292350
rect 159018 292226 159638 292294
rect 159018 292170 159114 292226
rect 159170 292170 159238 292226
rect 159294 292170 159362 292226
rect 159418 292170 159486 292226
rect 159542 292170 159638 292226
rect 159018 292102 159638 292170
rect 159018 292046 159114 292102
rect 159170 292046 159238 292102
rect 159294 292046 159362 292102
rect 159418 292046 159486 292102
rect 159542 292046 159638 292102
rect 159018 291978 159638 292046
rect 159018 291922 159114 291978
rect 159170 291922 159238 291978
rect 159294 291922 159362 291978
rect 159418 291922 159486 291978
rect 159542 291922 159638 291978
rect 140924 289828 140980 289838
rect 138572 282996 138628 283006
rect 132018 280294 132114 280350
rect 132170 280294 132238 280350
rect 132294 280294 132362 280350
rect 132418 280294 132486 280350
rect 132542 280294 132638 280350
rect 132018 280226 132638 280294
rect 132018 280170 132114 280226
rect 132170 280170 132238 280226
rect 132294 280170 132362 280226
rect 132418 280170 132486 280226
rect 132542 280170 132638 280226
rect 132018 280102 132638 280170
rect 132018 280046 132114 280102
rect 132170 280046 132238 280102
rect 132294 280046 132362 280102
rect 132418 280046 132486 280102
rect 132542 280046 132638 280102
rect 132018 279978 132638 280046
rect 132018 279922 132114 279978
rect 132170 279922 132238 279978
rect 132294 279922 132362 279978
rect 132418 279922 132486 279978
rect 132542 279922 132638 279978
rect 130172 250252 130228 250262
rect 132018 262350 132638 279922
rect 136892 281876 136948 281886
rect 133532 275698 133588 275708
rect 133532 265076 133588 275642
rect 133532 265010 133588 265020
rect 136892 264404 136948 281820
rect 136892 264338 136948 264348
rect 132018 262294 132114 262350
rect 132170 262294 132238 262350
rect 132294 262294 132362 262350
rect 132418 262294 132486 262350
rect 132542 262294 132638 262350
rect 132018 262226 132638 262294
rect 132018 262170 132114 262226
rect 132170 262170 132238 262226
rect 132294 262170 132362 262226
rect 132418 262170 132486 262226
rect 132542 262170 132638 262226
rect 132018 262102 132638 262170
rect 132018 262046 132114 262102
rect 132170 262046 132238 262102
rect 132294 262046 132362 262102
rect 132418 262046 132486 262102
rect 132542 262046 132638 262102
rect 132018 261978 132638 262046
rect 132018 261922 132114 261978
rect 132170 261922 132238 261978
rect 132294 261922 132362 261978
rect 132418 261922 132486 261978
rect 132542 261922 132638 261978
rect 128298 238294 128394 238350
rect 128450 238294 128518 238350
rect 128574 238294 128642 238350
rect 128698 238294 128766 238350
rect 128822 238294 128918 238350
rect 128298 238226 128918 238294
rect 128298 238170 128394 238226
rect 128450 238170 128518 238226
rect 128574 238170 128642 238226
rect 128698 238170 128766 238226
rect 128822 238170 128918 238226
rect 128298 238102 128918 238170
rect 128298 238046 128394 238102
rect 128450 238046 128518 238102
rect 128574 238046 128642 238102
rect 128698 238046 128766 238102
rect 128822 238046 128918 238102
rect 128298 237978 128918 238046
rect 128298 237922 128394 237978
rect 128450 237922 128518 237978
rect 128574 237922 128642 237978
rect 128698 237922 128766 237978
rect 128822 237922 128918 237978
rect 97578 220294 97674 220350
rect 97730 220294 97798 220350
rect 97854 220294 97922 220350
rect 97978 220294 98046 220350
rect 98102 220294 98198 220350
rect 97578 220226 98198 220294
rect 97578 220170 97674 220226
rect 97730 220170 97798 220226
rect 97854 220170 97922 220226
rect 97978 220170 98046 220226
rect 98102 220170 98198 220226
rect 97578 220102 98198 220170
rect 97578 220046 97674 220102
rect 97730 220046 97798 220102
rect 97854 220046 97922 220102
rect 97978 220046 98046 220102
rect 98102 220046 98198 220102
rect 97578 219978 98198 220046
rect 97578 219922 97674 219978
rect 97730 219922 97798 219978
rect 97854 219922 97922 219978
rect 97978 219922 98046 219978
rect 98102 219922 98198 219978
rect 86448 202350 86768 202384
rect 86448 202294 86518 202350
rect 86574 202294 86642 202350
rect 86698 202294 86768 202350
rect 86448 202226 86768 202294
rect 86448 202170 86518 202226
rect 86574 202170 86642 202226
rect 86698 202170 86768 202226
rect 86448 202102 86768 202170
rect 86448 202046 86518 202102
rect 86574 202046 86642 202102
rect 86698 202046 86768 202102
rect 86448 201978 86768 202046
rect 86448 201922 86518 201978
rect 86574 201922 86642 201978
rect 86698 201922 86768 201978
rect 86448 201888 86768 201922
rect 97578 202350 98198 219922
rect 126812 223636 126868 223646
rect 101808 208350 102128 208384
rect 101808 208294 101878 208350
rect 101934 208294 102002 208350
rect 102058 208294 102128 208350
rect 101808 208226 102128 208294
rect 101808 208170 101878 208226
rect 101934 208170 102002 208226
rect 102058 208170 102128 208226
rect 101808 208102 102128 208170
rect 101808 208046 101878 208102
rect 101934 208046 102002 208102
rect 102058 208046 102128 208102
rect 101808 207978 102128 208046
rect 101808 207922 101878 207978
rect 101934 207922 102002 207978
rect 102058 207922 102128 207978
rect 101808 207888 102128 207922
rect 97578 202294 97674 202350
rect 97730 202294 97798 202350
rect 97854 202294 97922 202350
rect 97978 202294 98046 202350
rect 98102 202294 98198 202350
rect 97578 202226 98198 202294
rect 97578 202170 97674 202226
rect 97730 202170 97798 202226
rect 97854 202170 97922 202226
rect 97978 202170 98046 202226
rect 98102 202170 98198 202226
rect 97578 202102 98198 202170
rect 97578 202046 97674 202102
rect 97730 202046 97798 202102
rect 97854 202046 97922 202102
rect 97978 202046 98046 202102
rect 98102 202046 98198 202102
rect 97578 201978 98198 202046
rect 97578 201922 97674 201978
rect 97730 201922 97798 201978
rect 97854 201922 97922 201978
rect 97978 201922 98046 201978
rect 98102 201922 98198 201978
rect 82684 199018 82740 199028
rect 82684 198548 82740 198962
rect 82684 198482 82740 198492
rect 82236 187058 82292 187068
rect 82684 186452 82740 186462
rect 82684 186058 82740 186396
rect 82684 185992 82740 186002
rect 86448 184350 86768 184384
rect 86448 184294 86518 184350
rect 86574 184294 86642 184350
rect 86698 184294 86768 184350
rect 86448 184226 86768 184294
rect 86448 184170 86518 184226
rect 86574 184170 86642 184226
rect 86698 184170 86768 184226
rect 86448 184102 86768 184170
rect 86448 184046 86518 184102
rect 86574 184046 86642 184102
rect 86698 184046 86768 184102
rect 86448 183978 86768 184046
rect 86448 183922 86518 183978
rect 86574 183922 86642 183978
rect 86698 183922 86768 183978
rect 86448 183888 86768 183922
rect 97578 184350 98198 201922
rect 117168 202350 117488 202384
rect 117168 202294 117238 202350
rect 117294 202294 117362 202350
rect 117418 202294 117488 202350
rect 117168 202226 117488 202294
rect 117168 202170 117238 202226
rect 117294 202170 117362 202226
rect 117418 202170 117488 202226
rect 117168 202102 117488 202170
rect 117168 202046 117238 202102
rect 117294 202046 117362 202102
rect 117418 202046 117488 202102
rect 117168 201978 117488 202046
rect 117168 201922 117238 201978
rect 117294 201922 117362 201978
rect 117418 201922 117488 201978
rect 117168 201888 117488 201922
rect 101808 190350 102128 190384
rect 101808 190294 101878 190350
rect 101934 190294 102002 190350
rect 102058 190294 102128 190350
rect 101808 190226 102128 190294
rect 101808 190170 101878 190226
rect 101934 190170 102002 190226
rect 102058 190170 102128 190226
rect 101808 190102 102128 190170
rect 101808 190046 101878 190102
rect 101934 190046 102002 190102
rect 102058 190046 102128 190102
rect 101808 189978 102128 190046
rect 101808 189922 101878 189978
rect 101934 189922 102002 189978
rect 102058 189922 102128 189978
rect 101808 189888 102128 189922
rect 126812 189140 126868 223580
rect 126924 221956 126980 221966
rect 126924 192500 126980 221900
rect 128298 220350 128918 237922
rect 132018 244350 132638 261922
rect 135212 261044 135268 261054
rect 133532 259700 133588 259710
rect 133532 251938 133588 259644
rect 135212 255358 135268 260988
rect 138572 260372 138628 282940
rect 140924 265076 140980 289772
rect 144060 284900 144116 284910
rect 142716 283220 142772 283230
rect 141036 271124 141092 271134
rect 141036 270658 141092 271068
rect 141036 270592 141092 270602
rect 140924 265010 140980 265020
rect 141036 268436 141092 268446
rect 141036 264718 141092 268380
rect 141036 264652 141092 264662
rect 142604 266420 142660 266430
rect 138572 260306 138628 260316
rect 142604 258598 142660 266364
rect 142716 261044 142772 283164
rect 144060 278908 144116 284844
rect 143948 278852 144116 278908
rect 143948 267148 144004 278852
rect 148448 274350 148768 274384
rect 148448 274294 148518 274350
rect 148574 274294 148642 274350
rect 148698 274294 148768 274350
rect 148448 274226 148768 274294
rect 148448 274170 148518 274226
rect 148574 274170 148642 274226
rect 148698 274170 148768 274226
rect 148448 274102 148768 274170
rect 148448 274046 148518 274102
rect 148574 274046 148642 274102
rect 148698 274046 148768 274102
rect 148448 273978 148768 274046
rect 148448 273922 148518 273978
rect 148574 273922 148642 273978
rect 148698 273922 148768 273978
rect 148448 273888 148768 273922
rect 159018 274350 159638 291922
rect 159018 274294 159114 274350
rect 159170 274294 159238 274350
rect 159294 274294 159362 274350
rect 159418 274294 159486 274350
rect 159542 274294 159638 274350
rect 159018 274226 159638 274294
rect 159018 274170 159114 274226
rect 159170 274170 159238 274226
rect 159294 274170 159362 274226
rect 159418 274170 159486 274226
rect 159542 274170 159638 274226
rect 159018 274102 159638 274170
rect 159018 274046 159114 274102
rect 159170 274046 159238 274102
rect 159294 274046 159362 274102
rect 159418 274046 159486 274102
rect 159542 274046 159638 274102
rect 159018 273978 159638 274046
rect 159018 273922 159114 273978
rect 159170 273922 159238 273978
rect 159294 273922 159362 273978
rect 159418 273922 159486 273978
rect 159542 273922 159638 273978
rect 144060 271198 144116 271208
rect 144060 271124 144116 271142
rect 144060 271058 144116 271068
rect 143948 267092 144116 267148
rect 142716 260978 142772 260988
rect 144060 260372 144116 267092
rect 144284 262836 144340 262846
rect 144284 260398 144340 262780
rect 144284 260332 144340 260342
rect 144060 260306 144116 260316
rect 142716 258598 142772 258608
rect 142604 258542 142716 258598
rect 142716 258532 142772 258542
rect 148448 256350 148768 256384
rect 148448 256294 148518 256350
rect 148574 256294 148642 256350
rect 148698 256294 148768 256350
rect 148448 256226 148768 256294
rect 148448 256170 148518 256226
rect 148574 256170 148642 256226
rect 148698 256170 148768 256226
rect 148448 256102 148768 256170
rect 148448 256046 148518 256102
rect 148574 256046 148642 256102
rect 148698 256046 148768 256102
rect 148448 255978 148768 256046
rect 148448 255922 148518 255978
rect 148574 255922 148642 255978
rect 148698 255922 148768 255978
rect 148448 255888 148768 255922
rect 159018 256350 159638 273922
rect 162738 298350 163358 315922
rect 162738 298294 162834 298350
rect 162890 298294 162958 298350
rect 163014 298294 163082 298350
rect 163138 298294 163206 298350
rect 163262 298294 163358 298350
rect 162738 298226 163358 298294
rect 162738 298170 162834 298226
rect 162890 298170 162958 298226
rect 163014 298170 163082 298226
rect 163138 298170 163206 298226
rect 163262 298170 163358 298226
rect 162738 298102 163358 298170
rect 162738 298046 162834 298102
rect 162890 298046 162958 298102
rect 163014 298046 163082 298102
rect 163138 298046 163206 298102
rect 163262 298046 163358 298102
rect 162738 297978 163358 298046
rect 162738 297922 162834 297978
rect 162890 297922 162958 297978
rect 163014 297922 163082 297978
rect 163138 297922 163206 297978
rect 163262 297922 163358 297978
rect 162738 280350 163358 297922
rect 189738 310350 190358 327922
rect 189738 310294 189834 310350
rect 189890 310294 189958 310350
rect 190014 310294 190082 310350
rect 190138 310294 190206 310350
rect 190262 310294 190358 310350
rect 189738 310226 190358 310294
rect 189738 310170 189834 310226
rect 189890 310170 189958 310226
rect 190014 310170 190082 310226
rect 190138 310170 190206 310226
rect 190262 310170 190358 310226
rect 189738 310102 190358 310170
rect 189738 310046 189834 310102
rect 189890 310046 189958 310102
rect 190014 310046 190082 310102
rect 190138 310046 190206 310102
rect 190262 310046 190358 310102
rect 189738 309978 190358 310046
rect 189738 309922 189834 309978
rect 189890 309922 189958 309978
rect 190014 309922 190082 309978
rect 190138 309922 190206 309978
rect 190262 309922 190358 309978
rect 189738 292350 190358 309922
rect 189738 292294 189834 292350
rect 189890 292294 189958 292350
rect 190014 292294 190082 292350
rect 190138 292294 190206 292350
rect 190262 292294 190358 292350
rect 189738 292226 190358 292294
rect 189738 292170 189834 292226
rect 189890 292170 189958 292226
rect 190014 292170 190082 292226
rect 190138 292170 190206 292226
rect 190262 292170 190358 292226
rect 189738 292102 190358 292170
rect 189738 292046 189834 292102
rect 189890 292046 189958 292102
rect 190014 292046 190082 292102
rect 190138 292046 190206 292102
rect 190262 292046 190358 292102
rect 189738 291978 190358 292046
rect 189738 291922 189834 291978
rect 189890 291922 189958 291978
rect 190014 291922 190082 291978
rect 190138 291922 190206 291978
rect 190262 291922 190358 291978
rect 189196 290276 189252 290286
rect 188972 289156 189028 289166
rect 162738 280294 162834 280350
rect 162890 280294 162958 280350
rect 163014 280294 163082 280350
rect 163138 280294 163206 280350
rect 163262 280294 163358 280350
rect 162738 280226 163358 280294
rect 162738 280170 162834 280226
rect 162890 280170 162958 280226
rect 163014 280170 163082 280226
rect 163138 280170 163206 280226
rect 163262 280170 163358 280226
rect 162738 280102 163358 280170
rect 162738 280046 162834 280102
rect 162890 280046 162958 280102
rect 163014 280046 163082 280102
rect 163138 280046 163206 280102
rect 163262 280046 163358 280102
rect 162738 279978 163358 280046
rect 162738 279922 162834 279978
rect 162890 279922 162958 279978
rect 163014 279922 163082 279978
rect 163138 279922 163206 279978
rect 163262 279922 163358 279978
rect 162738 266958 163358 279922
rect 163808 280350 164128 280384
rect 163808 280294 163878 280350
rect 163934 280294 164002 280350
rect 164058 280294 164128 280350
rect 163808 280226 164128 280294
rect 163808 280170 163878 280226
rect 163934 280170 164002 280226
rect 164058 280170 164128 280226
rect 163808 280102 164128 280170
rect 163808 280046 163878 280102
rect 163934 280046 164002 280102
rect 164058 280046 164128 280102
rect 163808 279978 164128 280046
rect 163808 279922 163878 279978
rect 163934 279922 164002 279978
rect 164058 279922 164128 279978
rect 163808 279888 164128 279922
rect 179168 274350 179488 274384
rect 179168 274294 179238 274350
rect 179294 274294 179362 274350
rect 179418 274294 179488 274350
rect 179168 274226 179488 274294
rect 179168 274170 179238 274226
rect 179294 274170 179362 274226
rect 179418 274170 179488 274226
rect 179168 274102 179488 274170
rect 179168 274046 179238 274102
rect 179294 274046 179362 274102
rect 179418 274046 179488 274102
rect 179168 273978 179488 274046
rect 179168 273922 179238 273978
rect 179294 273922 179362 273978
rect 179418 273922 179488 273978
rect 179168 273888 179488 273922
rect 163808 262350 164128 262384
rect 163808 262294 163878 262350
rect 163934 262294 164002 262350
rect 164058 262294 164128 262350
rect 163808 262226 164128 262294
rect 163808 262170 163878 262226
rect 163934 262170 164002 262226
rect 164058 262170 164128 262226
rect 163808 262102 164128 262170
rect 159018 256294 159114 256350
rect 159170 256294 159238 256350
rect 159294 256294 159362 256350
rect 159418 256294 159486 256350
rect 159542 256294 159638 256350
rect 159018 256226 159638 256294
rect 159018 256170 159114 256226
rect 159170 256170 159238 256226
rect 159294 256170 159362 256226
rect 159418 256170 159486 256226
rect 159542 256170 159638 256226
rect 159018 256102 159638 256170
rect 159018 256046 159114 256102
rect 159170 256046 159238 256102
rect 159294 256046 159362 256102
rect 159418 256046 159486 256102
rect 159542 256046 159638 256102
rect 159018 255978 159638 256046
rect 159018 255922 159114 255978
rect 159170 255922 159238 255978
rect 159294 255922 159362 255978
rect 159418 255922 159486 255978
rect 159542 255922 159638 255978
rect 135212 255292 135268 255302
rect 133532 251872 133588 251882
rect 132018 244294 132114 244350
rect 132170 244294 132238 244350
rect 132294 244294 132362 244350
rect 132418 244294 132486 244350
rect 132542 244294 132638 244350
rect 132018 244226 132638 244294
rect 132018 244170 132114 244226
rect 132170 244170 132238 244226
rect 132294 244170 132362 244226
rect 132418 244170 132486 244226
rect 132542 244170 132638 244226
rect 132018 244102 132638 244170
rect 132018 244046 132114 244102
rect 132170 244046 132238 244102
rect 132294 244046 132362 244102
rect 132418 244046 132486 244102
rect 132542 244046 132638 244102
rect 132018 243978 132638 244046
rect 132018 243922 132114 243978
rect 132170 243922 132238 243978
rect 132294 243922 132362 243978
rect 132418 243922 132486 243978
rect 132542 243922 132638 243978
rect 132018 226350 132638 243922
rect 159018 238350 159638 255922
rect 159018 238294 159114 238350
rect 159170 238294 159238 238350
rect 159294 238294 159362 238350
rect 159418 238294 159486 238350
rect 159542 238294 159638 238350
rect 159018 238226 159638 238294
rect 159018 238170 159114 238226
rect 159170 238170 159238 238226
rect 159294 238170 159362 238226
rect 159418 238170 159486 238226
rect 159542 238170 159638 238226
rect 159018 238102 159638 238170
rect 159018 238046 159114 238102
rect 159170 238046 159238 238102
rect 159294 238046 159362 238102
rect 159418 238046 159486 238102
rect 159542 238046 159638 238102
rect 159018 237978 159638 238046
rect 159018 237922 159114 237978
rect 159170 237922 159238 237978
rect 159294 237922 159362 237978
rect 159418 237922 159486 237978
rect 159542 237922 159638 237978
rect 132018 226294 132114 226350
rect 132170 226294 132238 226350
rect 132294 226294 132362 226350
rect 132418 226294 132486 226350
rect 132542 226294 132638 226350
rect 132018 226226 132638 226294
rect 132018 226170 132114 226226
rect 132170 226170 132238 226226
rect 132294 226170 132362 226226
rect 132418 226170 132486 226226
rect 132542 226170 132638 226226
rect 132018 226102 132638 226170
rect 132018 226046 132114 226102
rect 132170 226046 132238 226102
rect 132294 226046 132362 226102
rect 132418 226046 132486 226102
rect 132542 226046 132638 226102
rect 132018 225978 132638 226046
rect 132018 225922 132114 225978
rect 132170 225922 132238 225978
rect 132294 225922 132362 225978
rect 132418 225922 132486 225978
rect 132542 225922 132638 225978
rect 128298 220294 128394 220350
rect 128450 220294 128518 220350
rect 128574 220294 128642 220350
rect 128698 220294 128766 220350
rect 128822 220294 128918 220350
rect 128298 220226 128918 220294
rect 128298 220170 128394 220226
rect 128450 220170 128518 220226
rect 128574 220170 128642 220226
rect 128698 220170 128766 220226
rect 128822 220170 128918 220226
rect 128298 220102 128918 220170
rect 128298 220046 128394 220102
rect 128450 220046 128518 220102
rect 128574 220046 128642 220102
rect 128698 220046 128766 220102
rect 128822 220046 128918 220102
rect 128298 219978 128918 220046
rect 128298 219922 128394 219978
rect 128450 219922 128518 219978
rect 128574 219922 128642 219978
rect 128698 219922 128766 219978
rect 128822 219922 128918 219978
rect 128298 202350 128918 219922
rect 130172 220836 130228 220846
rect 130172 211204 130228 220780
rect 130172 211138 130228 211148
rect 128298 202294 128394 202350
rect 128450 202294 128518 202350
rect 128574 202294 128642 202350
rect 128698 202294 128766 202350
rect 128822 202294 128918 202350
rect 128298 202226 128918 202294
rect 128298 202170 128394 202226
rect 128450 202170 128518 202226
rect 128574 202170 128642 202226
rect 128698 202170 128766 202226
rect 128822 202170 128918 202226
rect 128298 202102 128918 202170
rect 128298 202046 128394 202102
rect 128450 202046 128518 202102
rect 128574 202046 128642 202102
rect 128698 202046 128766 202102
rect 128822 202046 128918 202102
rect 128298 201978 128918 202046
rect 128298 201922 128394 201978
rect 128450 201922 128518 201978
rect 128574 201922 128642 201978
rect 128698 201922 128766 201978
rect 128822 201922 128918 201978
rect 127484 195188 127540 195198
rect 127484 193978 127540 195132
rect 127484 193912 127540 193922
rect 127596 194516 127652 194526
rect 127596 193258 127652 194460
rect 127596 193192 127652 193202
rect 126924 192434 126980 192444
rect 126812 189074 126868 189084
rect 127596 191156 127652 191166
rect 127596 186238 127652 191100
rect 127596 186172 127652 186182
rect 97578 184294 97674 184350
rect 97730 184294 97798 184350
rect 97854 184294 97922 184350
rect 97978 184294 98046 184350
rect 98102 184294 98198 184350
rect 97578 184226 98198 184294
rect 97578 184170 97674 184226
rect 97730 184170 97798 184226
rect 97854 184170 97922 184226
rect 97978 184170 98046 184226
rect 98102 184170 98198 184226
rect 97578 184102 98198 184170
rect 97578 184046 97674 184102
rect 97730 184046 97798 184102
rect 97854 184046 97922 184102
rect 97978 184046 98046 184102
rect 98102 184046 98198 184102
rect 97578 183978 98198 184046
rect 97578 183922 97674 183978
rect 97730 183922 97798 183978
rect 97854 183922 97922 183978
rect 97978 183922 98046 183978
rect 98102 183922 98198 183978
rect 70578 172294 70674 172350
rect 70730 172294 70798 172350
rect 70854 172294 70922 172350
rect 70978 172294 71046 172350
rect 71102 172294 71198 172350
rect 70578 172226 71198 172294
rect 70578 172170 70674 172226
rect 70730 172170 70798 172226
rect 70854 172170 70922 172226
rect 70978 172170 71046 172226
rect 71102 172170 71198 172226
rect 70578 172102 71198 172170
rect 70578 172046 70674 172102
rect 70730 172046 70798 172102
rect 70854 172046 70922 172102
rect 70978 172046 71046 172102
rect 71102 172046 71198 172102
rect 70578 171978 71198 172046
rect 70578 171922 70674 171978
rect 70730 171922 70798 171978
rect 70854 171922 70922 171978
rect 70978 171922 71046 171978
rect 71102 171922 71198 171978
rect 70578 154350 71198 171922
rect 70578 154294 70674 154350
rect 70730 154294 70798 154350
rect 70854 154294 70922 154350
rect 70978 154294 71046 154350
rect 71102 154294 71198 154350
rect 70578 154226 71198 154294
rect 70578 154170 70674 154226
rect 70730 154170 70798 154226
rect 70854 154170 70922 154226
rect 70978 154170 71046 154226
rect 71102 154170 71198 154226
rect 70578 154102 71198 154170
rect 70578 154046 70674 154102
rect 70730 154046 70798 154102
rect 70854 154046 70922 154102
rect 70978 154046 71046 154102
rect 71102 154046 71198 154102
rect 70578 153978 71198 154046
rect 70578 153922 70674 153978
rect 70730 153922 70798 153978
rect 70854 153922 70922 153978
rect 70978 153922 71046 153978
rect 71102 153922 71198 153978
rect 66858 130294 66954 130350
rect 67010 130294 67078 130350
rect 67134 130294 67202 130350
rect 67258 130294 67326 130350
rect 67382 130294 67478 130350
rect 66858 130226 67478 130294
rect 66858 130170 66954 130226
rect 67010 130170 67078 130226
rect 67134 130170 67202 130226
rect 67258 130170 67326 130226
rect 67382 130170 67478 130226
rect 66858 130102 67478 130170
rect 66858 130046 66954 130102
rect 67010 130046 67078 130102
rect 67134 130046 67202 130102
rect 67258 130046 67326 130102
rect 67382 130046 67478 130102
rect 66858 129978 67478 130046
rect 66858 129922 66954 129978
rect 67010 129922 67078 129978
rect 67134 129922 67202 129978
rect 67258 129922 67326 129978
rect 67382 129922 67478 129978
rect 64652 117842 64708 117852
rect 64204 117478 64260 117488
rect 64204 116564 64260 117422
rect 64204 116498 64260 116508
rect 24448 112350 24768 112384
rect 24448 112294 24518 112350
rect 24574 112294 24642 112350
rect 24698 112294 24768 112350
rect 24448 112226 24768 112294
rect 24448 112170 24518 112226
rect 24574 112170 24642 112226
rect 24698 112170 24768 112226
rect 24448 112102 24768 112170
rect 24448 112046 24518 112102
rect 24574 112046 24642 112102
rect 24698 112046 24768 112102
rect 24448 111978 24768 112046
rect 24448 111922 24518 111978
rect 24574 111922 24642 111978
rect 24698 111922 24768 111978
rect 24448 111888 24768 111922
rect 36138 112350 36758 114770
rect 36138 112294 36234 112350
rect 36290 112294 36358 112350
rect 36414 112294 36482 112350
rect 36538 112294 36606 112350
rect 36662 112294 36758 112350
rect 36138 112226 36758 112294
rect 36138 112170 36234 112226
rect 36290 112170 36358 112226
rect 36414 112170 36482 112226
rect 36538 112170 36606 112226
rect 36662 112170 36758 112226
rect 36138 112102 36758 112170
rect 36138 112046 36234 112102
rect 36290 112046 36358 112102
rect 36414 112046 36482 112102
rect 36538 112046 36606 112102
rect 36662 112046 36758 112102
rect 36138 111978 36758 112046
rect 36138 111922 36234 111978
rect 36290 111922 36358 111978
rect 36414 111922 36482 111978
rect 36538 111922 36606 111978
rect 36662 111922 36758 111978
rect 9138 100294 9234 100350
rect 9290 100294 9358 100350
rect 9414 100294 9482 100350
rect 9538 100294 9606 100350
rect 9662 100294 9758 100350
rect 9138 100226 9758 100294
rect 9138 100170 9234 100226
rect 9290 100170 9358 100226
rect 9414 100170 9482 100226
rect 9538 100170 9606 100226
rect 9662 100170 9758 100226
rect 9138 100102 9758 100170
rect 9138 100046 9234 100102
rect 9290 100046 9358 100102
rect 9414 100046 9482 100102
rect 9538 100046 9606 100102
rect 9662 100046 9758 100102
rect 9138 99978 9758 100046
rect 9138 99922 9234 99978
rect 9290 99922 9358 99978
rect 9414 99922 9482 99978
rect 9538 99922 9606 99978
rect 9662 99922 9758 99978
rect 9138 82350 9758 99922
rect 9138 82294 9234 82350
rect 9290 82294 9358 82350
rect 9414 82294 9482 82350
rect 9538 82294 9606 82350
rect 9662 82294 9758 82350
rect 9138 82226 9758 82294
rect 9138 82170 9234 82226
rect 9290 82170 9358 82226
rect 9414 82170 9482 82226
rect 9538 82170 9606 82226
rect 9662 82170 9758 82226
rect 9138 82102 9758 82170
rect 9138 82046 9234 82102
rect 9290 82046 9358 82102
rect 9414 82046 9482 82102
rect 9538 82046 9606 82102
rect 9662 82046 9758 82102
rect 9138 81978 9758 82046
rect 9138 81922 9234 81978
rect 9290 81922 9358 81978
rect 9414 81922 9482 81978
rect 9538 81922 9606 81978
rect 9662 81922 9758 81978
rect 9138 64350 9758 81922
rect 36138 94350 36758 111922
rect 55168 112350 55488 112384
rect 55168 112294 55238 112350
rect 55294 112294 55362 112350
rect 55418 112294 55488 112350
rect 55168 112226 55488 112294
rect 55168 112170 55238 112226
rect 55294 112170 55362 112226
rect 55418 112170 55488 112226
rect 55168 112102 55488 112170
rect 55168 112046 55238 112102
rect 55294 112046 55362 112102
rect 55418 112046 55488 112102
rect 55168 111978 55488 112046
rect 55168 111922 55238 111978
rect 55294 111922 55362 111978
rect 55418 111922 55488 111978
rect 55168 111888 55488 111922
rect 66858 112350 67478 129922
rect 69692 147028 69748 147038
rect 69692 124628 69748 146972
rect 69692 124562 69748 124572
rect 70578 136350 71198 153922
rect 97578 166350 98198 183922
rect 117168 184350 117488 184384
rect 117168 184294 117238 184350
rect 117294 184294 117362 184350
rect 117418 184294 117488 184350
rect 117168 184226 117488 184294
rect 117168 184170 117238 184226
rect 117294 184170 117362 184226
rect 117418 184170 117488 184226
rect 117168 184102 117488 184170
rect 117168 184046 117238 184102
rect 117294 184046 117362 184102
rect 117418 184046 117488 184102
rect 117168 183978 117488 184046
rect 117168 183922 117238 183978
rect 117294 183922 117362 183978
rect 117418 183922 117488 183978
rect 117168 183888 117488 183922
rect 128298 184350 128918 201922
rect 128298 184294 128394 184350
rect 128450 184294 128518 184350
rect 128574 184294 128642 184350
rect 128698 184294 128766 184350
rect 128822 184294 128918 184350
rect 128298 184226 128918 184294
rect 128298 184170 128394 184226
rect 128450 184170 128518 184226
rect 128574 184170 128642 184226
rect 128698 184170 128766 184226
rect 128822 184170 128918 184226
rect 128298 184102 128918 184170
rect 128298 184046 128394 184102
rect 128450 184046 128518 184102
rect 128574 184046 128642 184102
rect 128698 184046 128766 184102
rect 128822 184046 128918 184102
rect 128298 183978 128918 184046
rect 128298 183922 128394 183978
rect 128450 183922 128518 183978
rect 128574 183922 128642 183978
rect 128698 183922 128766 183978
rect 128822 183922 128918 183978
rect 97578 166294 97674 166350
rect 97730 166294 97798 166350
rect 97854 166294 97922 166350
rect 97978 166294 98046 166350
rect 98102 166294 98198 166350
rect 97578 166226 98198 166294
rect 97578 166170 97674 166226
rect 97730 166170 97798 166226
rect 97854 166170 97922 166226
rect 97978 166170 98046 166226
rect 98102 166170 98198 166226
rect 97578 166102 98198 166170
rect 97578 166046 97674 166102
rect 97730 166046 97798 166102
rect 97854 166046 97922 166102
rect 97978 166046 98046 166102
rect 98102 166046 98198 166102
rect 97578 165978 98198 166046
rect 97578 165922 97674 165978
rect 97730 165922 97798 165978
rect 97854 165922 97922 165978
rect 97978 165922 98046 165978
rect 98102 165922 98198 165978
rect 81452 150500 81508 150510
rect 70578 136294 70674 136350
rect 70730 136294 70798 136350
rect 70854 136294 70922 136350
rect 70978 136294 71046 136350
rect 71102 136294 71198 136350
rect 70578 136226 71198 136294
rect 70578 136170 70674 136226
rect 70730 136170 70798 136226
rect 70854 136170 70922 136226
rect 70978 136170 71046 136226
rect 71102 136170 71198 136226
rect 70578 136102 71198 136170
rect 70578 136046 70674 136102
rect 70730 136046 70798 136102
rect 70854 136046 70922 136102
rect 70978 136046 71046 136102
rect 71102 136046 71198 136102
rect 70578 135978 71198 136046
rect 70578 135922 70674 135978
rect 70730 135922 70798 135978
rect 70854 135922 70922 135978
rect 70978 135922 71046 135978
rect 71102 135922 71198 135978
rect 66858 112294 66954 112350
rect 67010 112294 67078 112350
rect 67134 112294 67202 112350
rect 67258 112294 67326 112350
rect 67382 112294 67478 112350
rect 66858 112226 67478 112294
rect 66858 112170 66954 112226
rect 67010 112170 67078 112226
rect 67134 112170 67202 112226
rect 67258 112170 67326 112226
rect 67382 112170 67478 112226
rect 66858 112102 67478 112170
rect 66858 112046 66954 112102
rect 67010 112046 67078 112102
rect 67134 112046 67202 112102
rect 67258 112046 67326 112102
rect 67382 112046 67478 112102
rect 66858 111978 67478 112046
rect 66858 111922 66954 111978
rect 67010 111922 67078 111978
rect 67134 111922 67202 111978
rect 67258 111922 67326 111978
rect 67382 111922 67478 111978
rect 36138 94294 36234 94350
rect 36290 94294 36358 94350
rect 36414 94294 36482 94350
rect 36538 94294 36606 94350
rect 36662 94294 36758 94350
rect 36138 94226 36758 94294
rect 36138 94170 36234 94226
rect 36290 94170 36358 94226
rect 36414 94170 36482 94226
rect 36538 94170 36606 94226
rect 36662 94170 36758 94226
rect 36138 94102 36758 94170
rect 36138 94046 36234 94102
rect 36290 94046 36358 94102
rect 36414 94046 36482 94102
rect 36538 94046 36606 94102
rect 36662 94046 36758 94102
rect 36138 93978 36758 94046
rect 36138 93922 36234 93978
rect 36290 93922 36358 93978
rect 36414 93922 36482 93978
rect 36538 93922 36606 93978
rect 36662 93922 36758 93978
rect 36138 76350 36758 93922
rect 36138 76294 36234 76350
rect 36290 76294 36358 76350
rect 36414 76294 36482 76350
rect 36538 76294 36606 76350
rect 36662 76294 36758 76350
rect 36138 76226 36758 76294
rect 36138 76170 36234 76226
rect 36290 76170 36358 76226
rect 36414 76170 36482 76226
rect 36538 76170 36606 76226
rect 36662 76170 36758 76226
rect 36138 76102 36758 76170
rect 36138 76046 36234 76102
rect 36290 76046 36358 76102
rect 36414 76046 36482 76102
rect 36538 76046 36606 76102
rect 36662 76046 36758 76102
rect 36138 75978 36758 76046
rect 36138 75922 36234 75978
rect 36290 75922 36358 75978
rect 36414 75922 36482 75978
rect 36538 75922 36606 75978
rect 36662 75922 36758 75978
rect 20636 70196 20692 70206
rect 19964 68516 20020 68526
rect 9138 64294 9234 64350
rect 9290 64294 9358 64350
rect 9414 64294 9482 64350
rect 9538 64294 9606 64350
rect 9662 64294 9758 64350
rect 9138 64226 9758 64294
rect 9138 64170 9234 64226
rect 9290 64170 9358 64226
rect 9414 64170 9482 64226
rect 9538 64170 9606 64226
rect 9662 64170 9758 64226
rect 9138 64102 9758 64170
rect 9138 64046 9234 64102
rect 9290 64046 9358 64102
rect 9414 64046 9482 64102
rect 9538 64046 9606 64102
rect 9662 64046 9758 64102
rect 9138 63978 9758 64046
rect 9138 63922 9234 63978
rect 9290 63922 9358 63978
rect 9414 63922 9482 63978
rect 9538 63922 9606 63978
rect 9662 63922 9758 63978
rect 9138 46350 9758 63922
rect 9138 46294 9234 46350
rect 9290 46294 9358 46350
rect 9414 46294 9482 46350
rect 9538 46294 9606 46350
rect 9662 46294 9758 46350
rect 9138 46226 9758 46294
rect 9138 46170 9234 46226
rect 9290 46170 9358 46226
rect 9414 46170 9482 46226
rect 9538 46170 9606 46226
rect 9662 46170 9758 46226
rect 9138 46102 9758 46170
rect 9138 46046 9234 46102
rect 9290 46046 9358 46102
rect 9414 46046 9482 46102
rect 9538 46046 9606 46102
rect 9662 46046 9758 46102
rect 9138 45978 9758 46046
rect 9138 45922 9234 45978
rect 9290 45922 9358 45978
rect 9414 45922 9482 45978
rect 9538 45922 9606 45978
rect 9662 45922 9758 45978
rect 9138 28350 9758 45922
rect 18284 67284 18340 67294
rect 18284 45444 18340 67228
rect 18284 45378 18340 45388
rect 18396 56868 18452 56878
rect 18396 55558 18452 56812
rect 9138 28294 9234 28350
rect 9290 28294 9358 28350
rect 9414 28294 9482 28350
rect 9538 28294 9606 28350
rect 9662 28294 9758 28350
rect 9138 28226 9758 28294
rect 9138 28170 9234 28226
rect 9290 28170 9358 28226
rect 9414 28170 9482 28226
rect 9538 28170 9606 28226
rect 9662 28170 9758 28226
rect 9138 28102 9758 28170
rect 9138 28046 9234 28102
rect 9290 28046 9358 28102
rect 9414 28046 9482 28102
rect 9538 28046 9606 28102
rect 9662 28046 9758 28102
rect 9138 27978 9758 28046
rect 9138 27922 9234 27978
rect 9290 27922 9358 27978
rect 9414 27922 9482 27978
rect 9538 27922 9606 27978
rect 9662 27922 9758 27978
rect 9138 10350 9758 27922
rect 9138 10294 9234 10350
rect 9290 10294 9358 10350
rect 9414 10294 9482 10350
rect 9538 10294 9606 10350
rect 9662 10294 9758 10350
rect 9138 10226 9758 10294
rect 9138 10170 9234 10226
rect 9290 10170 9358 10226
rect 9414 10170 9482 10226
rect 9538 10170 9606 10226
rect 9662 10170 9758 10226
rect 9138 10102 9758 10170
rect 9138 10046 9234 10102
rect 9290 10046 9358 10102
rect 9414 10046 9482 10102
rect 9538 10046 9606 10102
rect 9662 10046 9758 10102
rect 9138 9978 9758 10046
rect 9138 9922 9234 9978
rect 9290 9922 9358 9978
rect 9414 9922 9482 9978
rect 9538 9922 9606 9978
rect 9662 9922 9758 9978
rect 9138 -1120 9758 9922
rect 18396 5124 18452 55502
rect 19964 48244 20020 68460
rect 20076 67956 20132 67966
rect 20076 55524 20132 67900
rect 20636 67284 20692 70140
rect 20636 67218 20692 67228
rect 24448 58350 24768 58384
rect 24448 58294 24518 58350
rect 24574 58294 24642 58350
rect 24698 58294 24768 58350
rect 24448 58226 24768 58294
rect 24448 58170 24518 58226
rect 24574 58170 24642 58226
rect 24698 58170 24768 58226
rect 24448 58102 24768 58170
rect 24448 58046 24518 58102
rect 24574 58046 24642 58102
rect 24698 58046 24768 58102
rect 24448 57978 24768 58046
rect 24448 57922 24518 57978
rect 24574 57922 24642 57978
rect 24698 57922 24768 57978
rect 24448 57888 24768 57922
rect 36138 58350 36758 75922
rect 39858 100350 40478 101364
rect 39858 100294 39954 100350
rect 40010 100294 40078 100350
rect 40134 100294 40202 100350
rect 40258 100294 40326 100350
rect 40382 100294 40478 100350
rect 39858 100226 40478 100294
rect 39858 100170 39954 100226
rect 40010 100170 40078 100226
rect 40134 100170 40202 100226
rect 40258 100170 40326 100226
rect 40382 100170 40478 100226
rect 39858 100102 40478 100170
rect 39858 100046 39954 100102
rect 40010 100046 40078 100102
rect 40134 100046 40202 100102
rect 40258 100046 40326 100102
rect 40382 100046 40478 100102
rect 39858 99978 40478 100046
rect 39858 99922 39954 99978
rect 40010 99922 40078 99978
rect 40134 99922 40202 99978
rect 40258 99922 40326 99978
rect 40382 99922 40478 99978
rect 39858 82350 40478 99922
rect 39858 82294 39954 82350
rect 40010 82294 40078 82350
rect 40134 82294 40202 82350
rect 40258 82294 40326 82350
rect 40382 82294 40478 82350
rect 39858 82226 40478 82294
rect 39858 82170 39954 82226
rect 40010 82170 40078 82226
rect 40134 82170 40202 82226
rect 40258 82170 40326 82226
rect 40382 82170 40478 82226
rect 39858 82102 40478 82170
rect 39858 82046 39954 82102
rect 40010 82046 40078 82102
rect 40134 82046 40202 82102
rect 40258 82046 40326 82102
rect 40382 82046 40478 82102
rect 39858 81978 40478 82046
rect 39858 81922 39954 81978
rect 40010 81922 40078 81978
rect 40134 81922 40202 81978
rect 40258 81922 40326 81978
rect 40382 81922 40478 81978
rect 39858 69788 40478 81922
rect 66858 94350 67478 111922
rect 70578 118350 71198 135922
rect 80332 139524 80388 139534
rect 73836 126118 73892 126128
rect 73836 120596 73892 126062
rect 80332 123956 80388 139468
rect 80332 123890 80388 123900
rect 80444 132778 80500 132788
rect 80444 122500 80500 132722
rect 81452 124068 81508 150444
rect 97578 148350 98198 165922
rect 97578 148294 97674 148350
rect 97730 148294 97798 148350
rect 97854 148294 97922 148350
rect 97978 148294 98046 148350
rect 98102 148294 98198 148350
rect 97578 148226 98198 148294
rect 97578 148170 97674 148226
rect 97730 148170 97798 148226
rect 97854 148170 97922 148226
rect 97978 148170 98046 148226
rect 98102 148170 98198 148226
rect 97578 148102 98198 148170
rect 97578 148046 97674 148102
rect 97730 148046 97798 148102
rect 97854 148046 97922 148102
rect 97978 148046 98046 148102
rect 98102 148046 98198 148102
rect 97578 147978 98198 148046
rect 97578 147922 97674 147978
rect 97730 147922 97798 147978
rect 97854 147922 97922 147978
rect 97978 147922 98046 147978
rect 98102 147922 98198 147978
rect 86448 130350 86768 130384
rect 86448 130294 86518 130350
rect 86574 130294 86642 130350
rect 86698 130294 86768 130350
rect 86448 130226 86768 130294
rect 86448 130170 86518 130226
rect 86574 130170 86642 130226
rect 86698 130170 86768 130226
rect 86448 130102 86768 130170
rect 86448 130046 86518 130102
rect 86574 130046 86642 130102
rect 86698 130046 86768 130102
rect 86448 129978 86768 130046
rect 86448 129922 86518 129978
rect 86574 129922 86642 129978
rect 86698 129922 86768 129978
rect 86448 129888 86768 129922
rect 97578 130350 98198 147922
rect 101298 172350 101918 172564
rect 101298 172294 101394 172350
rect 101450 172294 101518 172350
rect 101574 172294 101642 172350
rect 101698 172294 101766 172350
rect 101822 172294 101918 172350
rect 101298 172226 101918 172294
rect 101298 172170 101394 172226
rect 101450 172170 101518 172226
rect 101574 172170 101642 172226
rect 101698 172170 101766 172226
rect 101822 172170 101918 172226
rect 101298 172102 101918 172170
rect 101298 172046 101394 172102
rect 101450 172046 101518 172102
rect 101574 172046 101642 172102
rect 101698 172046 101766 172102
rect 101822 172046 101918 172102
rect 101298 171978 101918 172046
rect 101298 171922 101394 171978
rect 101450 171922 101518 171978
rect 101574 171922 101642 171978
rect 101698 171922 101766 171978
rect 101822 171922 101918 171978
rect 101298 154350 101918 171922
rect 128298 166350 128918 183922
rect 128298 166294 128394 166350
rect 128450 166294 128518 166350
rect 128574 166294 128642 166350
rect 128698 166294 128766 166350
rect 128822 166294 128918 166350
rect 128298 166226 128918 166294
rect 128298 166170 128394 166226
rect 128450 166170 128518 166226
rect 128574 166170 128642 166226
rect 128698 166170 128766 166226
rect 128822 166170 128918 166226
rect 128298 166102 128918 166170
rect 128298 166046 128394 166102
rect 128450 166046 128518 166102
rect 128574 166046 128642 166102
rect 128698 166046 128766 166102
rect 128822 166046 128918 166102
rect 128298 165978 128918 166046
rect 128298 165922 128394 165978
rect 128450 165922 128518 165978
rect 128574 165922 128642 165978
rect 128698 165922 128766 165978
rect 128822 165922 128918 165978
rect 127148 164276 127204 164286
rect 126924 163716 126980 163726
rect 101298 154294 101394 154350
rect 101450 154294 101518 154350
rect 101574 154294 101642 154350
rect 101698 154294 101766 154350
rect 101822 154294 101918 154350
rect 101298 154226 101918 154294
rect 101298 154170 101394 154226
rect 101450 154170 101518 154226
rect 101574 154170 101642 154226
rect 101698 154170 101766 154226
rect 101822 154170 101918 154226
rect 101298 154102 101918 154170
rect 101298 154046 101394 154102
rect 101450 154046 101518 154102
rect 101574 154046 101642 154102
rect 101698 154046 101766 154102
rect 101822 154046 101918 154102
rect 101298 153978 101918 154046
rect 101298 153922 101394 153978
rect 101450 153922 101518 153978
rect 101574 153922 101642 153978
rect 101698 153922 101766 153978
rect 101822 153922 101918 153978
rect 101298 140988 101918 153922
rect 126812 161476 126868 161486
rect 101808 136350 102128 136384
rect 101808 136294 101878 136350
rect 101934 136294 102002 136350
rect 102058 136294 102128 136350
rect 101808 136226 102128 136294
rect 101808 136170 101878 136226
rect 101934 136170 102002 136226
rect 102058 136170 102128 136226
rect 101808 136102 102128 136170
rect 101808 136046 101878 136102
rect 101934 136046 102002 136102
rect 102058 136046 102128 136102
rect 101808 135978 102128 136046
rect 101808 135922 101878 135978
rect 101934 135922 102002 135978
rect 102058 135922 102128 135978
rect 101808 135888 102128 135922
rect 97578 130294 97674 130350
rect 97730 130294 97798 130350
rect 97854 130294 97922 130350
rect 97978 130294 98046 130350
rect 98102 130294 98198 130350
rect 97578 130226 98198 130294
rect 97578 130170 97674 130226
rect 97730 130170 97798 130226
rect 97854 130170 97922 130226
rect 97978 130170 98046 130226
rect 98102 130170 98198 130226
rect 97578 130102 98198 130170
rect 97578 130046 97674 130102
rect 97730 130046 97798 130102
rect 97854 130046 97922 130102
rect 97978 130046 98046 130102
rect 98102 130046 98198 130102
rect 97578 129978 98198 130046
rect 97578 129922 97674 129978
rect 97730 129922 97798 129978
rect 97854 129922 97922 129978
rect 97978 129922 98046 129978
rect 98102 129922 98198 129978
rect 82684 127738 82740 127748
rect 82684 127316 82740 127682
rect 82684 127250 82740 127260
rect 82460 125938 82516 125948
rect 82460 125524 82516 125882
rect 82460 125458 82516 125468
rect 81452 124002 81508 124012
rect 80444 122434 80500 122444
rect 73836 120530 73892 120540
rect 70578 118294 70674 118350
rect 70730 118294 70798 118350
rect 70854 118294 70922 118350
rect 70978 118294 71046 118350
rect 71102 118294 71198 118350
rect 70578 118226 71198 118294
rect 70578 118170 70674 118226
rect 70730 118170 70798 118226
rect 70854 118170 70922 118226
rect 70978 118170 71046 118226
rect 71102 118170 71198 118226
rect 70578 118102 71198 118170
rect 70578 118046 70674 118102
rect 70730 118046 70798 118102
rect 70854 118046 70922 118102
rect 70978 118046 71046 118102
rect 71102 118046 71198 118102
rect 70578 117978 71198 118046
rect 70578 117922 70674 117978
rect 70730 117922 70798 117978
rect 70854 117922 70922 117978
rect 70978 117922 71046 117978
rect 71102 117922 71198 117978
rect 70578 100350 71198 117922
rect 86448 112350 86768 112384
rect 86448 112294 86518 112350
rect 86574 112294 86642 112350
rect 86698 112294 86768 112350
rect 86448 112226 86768 112294
rect 86448 112170 86518 112226
rect 86574 112170 86642 112226
rect 86698 112170 86768 112226
rect 86448 112102 86768 112170
rect 86448 112046 86518 112102
rect 86574 112046 86642 112102
rect 86698 112046 86768 112102
rect 86448 111978 86768 112046
rect 86448 111922 86518 111978
rect 86574 111922 86642 111978
rect 86698 111922 86768 111978
rect 86448 111888 86768 111922
rect 97578 112350 98198 129922
rect 117168 130350 117488 130384
rect 117168 130294 117238 130350
rect 117294 130294 117362 130350
rect 117418 130294 117488 130350
rect 117168 130226 117488 130294
rect 117168 130170 117238 130226
rect 117294 130170 117362 130226
rect 117418 130170 117488 130226
rect 117168 130102 117488 130170
rect 117168 130046 117238 130102
rect 117294 130046 117362 130102
rect 117418 130046 117488 130102
rect 117168 129978 117488 130046
rect 117168 129922 117238 129978
rect 117294 129922 117362 129978
rect 117418 129922 117488 129978
rect 117168 129888 117488 129922
rect 126812 119252 126868 161420
rect 126924 122612 126980 163660
rect 126924 122546 126980 122556
rect 127036 159796 127092 159806
rect 127036 119924 127092 159740
rect 127148 121940 127204 164220
rect 127372 163156 127428 163166
rect 127260 162596 127316 162606
rect 127260 126644 127316 162540
rect 127260 126578 127316 126588
rect 127372 125972 127428 163100
rect 127484 160916 127540 160926
rect 127484 136724 127540 160860
rect 127484 136658 127540 136668
rect 128298 148350 128918 165922
rect 128298 148294 128394 148350
rect 128450 148294 128518 148350
rect 128574 148294 128642 148350
rect 128698 148294 128766 148350
rect 128822 148294 128918 148350
rect 128298 148226 128918 148294
rect 128298 148170 128394 148226
rect 128450 148170 128518 148226
rect 128574 148170 128642 148226
rect 128698 148170 128766 148226
rect 128822 148170 128918 148226
rect 128298 148102 128918 148170
rect 128298 148046 128394 148102
rect 128450 148046 128518 148102
rect 128574 148046 128642 148102
rect 128698 148046 128766 148102
rect 128822 148046 128918 148102
rect 128298 147978 128918 148046
rect 128298 147922 128394 147978
rect 128450 147922 128518 147978
rect 128574 147922 128642 147978
rect 128698 147922 128766 147978
rect 128822 147922 128918 147978
rect 127372 125906 127428 125916
rect 128298 130350 128918 147922
rect 128298 130294 128394 130350
rect 128450 130294 128518 130350
rect 128574 130294 128642 130350
rect 128698 130294 128766 130350
rect 128822 130294 128918 130350
rect 128298 130226 128918 130294
rect 128298 130170 128394 130226
rect 128450 130170 128518 130226
rect 128574 130170 128642 130226
rect 128698 130170 128766 130226
rect 128822 130170 128918 130226
rect 128298 130102 128918 130170
rect 128298 130046 128394 130102
rect 128450 130046 128518 130102
rect 128574 130046 128642 130102
rect 128698 130046 128766 130102
rect 128822 130046 128918 130102
rect 128298 129978 128918 130046
rect 128298 129922 128394 129978
rect 128450 129922 128518 129978
rect 128574 129922 128642 129978
rect 128698 129922 128766 129978
rect 128822 129922 128918 129978
rect 127148 121874 127204 121884
rect 127036 119858 127092 119868
rect 126812 119186 126868 119196
rect 101808 118350 102128 118384
rect 101808 118294 101878 118350
rect 101934 118294 102002 118350
rect 102058 118294 102128 118350
rect 101808 118226 102128 118294
rect 101808 118170 101878 118226
rect 101934 118170 102002 118226
rect 102058 118170 102128 118226
rect 101808 118102 102128 118170
rect 101808 118046 101878 118102
rect 101934 118046 102002 118102
rect 102058 118046 102128 118102
rect 101808 117978 102128 118046
rect 101808 117922 101878 117978
rect 101934 117922 102002 117978
rect 102058 117922 102128 117978
rect 101808 117888 102128 117922
rect 97578 112294 97674 112350
rect 97730 112294 97798 112350
rect 97854 112294 97922 112350
rect 97978 112294 98046 112350
rect 98102 112294 98198 112350
rect 97578 112226 98198 112294
rect 97578 112170 97674 112226
rect 97730 112170 97798 112226
rect 97854 112170 97922 112226
rect 97978 112170 98046 112226
rect 98102 112170 98198 112226
rect 97578 112102 98198 112170
rect 97578 112046 97674 112102
rect 97730 112046 97798 112102
rect 97854 112046 97922 112102
rect 97978 112046 98046 112102
rect 98102 112046 98198 112102
rect 97578 111978 98198 112046
rect 97578 111922 97674 111978
rect 97730 111922 97798 111978
rect 97854 111922 97922 111978
rect 97978 111922 98046 111978
rect 98102 111922 98198 111978
rect 70578 100294 70674 100350
rect 70730 100294 70798 100350
rect 70854 100294 70922 100350
rect 70978 100294 71046 100350
rect 71102 100294 71198 100350
rect 70578 100226 71198 100294
rect 70578 100170 70674 100226
rect 70730 100170 70798 100226
rect 70854 100170 70922 100226
rect 70978 100170 71046 100226
rect 71102 100170 71198 100226
rect 70578 100102 71198 100170
rect 70578 100046 70674 100102
rect 70730 100046 70798 100102
rect 70854 100046 70922 100102
rect 70978 100046 71046 100102
rect 71102 100046 71198 100102
rect 70578 99978 71198 100046
rect 70578 99922 70674 99978
rect 70730 99922 70798 99978
rect 70854 99922 70922 99978
rect 70978 99922 71046 99978
rect 71102 99922 71198 99978
rect 66858 94294 66954 94350
rect 67010 94294 67078 94350
rect 67134 94294 67202 94350
rect 67258 94294 67326 94350
rect 67382 94294 67478 94350
rect 66858 94226 67478 94294
rect 66858 94170 66954 94226
rect 67010 94170 67078 94226
rect 67134 94170 67202 94226
rect 67258 94170 67326 94226
rect 67382 94170 67478 94226
rect 66858 94102 67478 94170
rect 66858 94046 66954 94102
rect 67010 94046 67078 94102
rect 67134 94046 67202 94102
rect 67258 94046 67326 94102
rect 67382 94046 67478 94102
rect 66858 93978 67478 94046
rect 66858 93922 66954 93978
rect 67010 93922 67078 93978
rect 67134 93922 67202 93978
rect 67258 93922 67326 93978
rect 67382 93922 67478 93978
rect 66858 76350 67478 93922
rect 66858 76294 66954 76350
rect 67010 76294 67078 76350
rect 67134 76294 67202 76350
rect 67258 76294 67326 76350
rect 67382 76294 67478 76350
rect 66858 76226 67478 76294
rect 66858 76170 66954 76226
rect 67010 76170 67078 76226
rect 67134 76170 67202 76226
rect 67258 76170 67326 76226
rect 67382 76170 67478 76226
rect 66858 76102 67478 76170
rect 66858 76046 66954 76102
rect 67010 76046 67078 76102
rect 67134 76046 67202 76102
rect 67258 76046 67326 76102
rect 67382 76046 67478 76102
rect 66858 75978 67478 76046
rect 66858 75922 66954 75978
rect 67010 75922 67078 75978
rect 67134 75922 67202 75978
rect 67258 75922 67326 75978
rect 67382 75922 67478 75978
rect 64652 70756 64708 70766
rect 39808 64350 40128 64384
rect 39808 64294 39878 64350
rect 39934 64294 40002 64350
rect 40058 64294 40128 64350
rect 39808 64226 40128 64294
rect 39808 64170 39878 64226
rect 39934 64170 40002 64226
rect 40058 64170 40128 64226
rect 39808 64102 40128 64170
rect 39808 64046 39878 64102
rect 39934 64046 40002 64102
rect 40058 64046 40128 64102
rect 39808 63978 40128 64046
rect 39808 63922 39878 63978
rect 39934 63922 40002 63978
rect 40058 63922 40128 63978
rect 39808 63888 40128 63922
rect 36138 58294 36234 58350
rect 36290 58294 36358 58350
rect 36414 58294 36482 58350
rect 36538 58294 36606 58350
rect 36662 58294 36758 58350
rect 36138 58226 36758 58294
rect 36138 58170 36234 58226
rect 36290 58170 36358 58226
rect 36414 58170 36482 58226
rect 36538 58170 36606 58226
rect 36662 58170 36758 58226
rect 36138 58102 36758 58170
rect 36138 58046 36234 58102
rect 36290 58046 36358 58102
rect 36414 58046 36482 58102
rect 36538 58046 36606 58102
rect 36662 58046 36758 58102
rect 36138 57978 36758 58046
rect 36138 57922 36234 57978
rect 36290 57922 36358 57978
rect 36414 57922 36482 57978
rect 36538 57922 36606 57978
rect 36662 57922 36758 57978
rect 20076 55458 20132 55468
rect 19964 48178 20020 48188
rect 24448 40350 24768 40384
rect 24448 40294 24518 40350
rect 24574 40294 24642 40350
rect 24698 40294 24768 40350
rect 24448 40226 24768 40294
rect 24448 40170 24518 40226
rect 24574 40170 24642 40226
rect 24698 40170 24768 40226
rect 24448 40102 24768 40170
rect 24448 40046 24518 40102
rect 24574 40046 24642 40102
rect 24698 40046 24768 40102
rect 24448 39978 24768 40046
rect 24448 39922 24518 39978
rect 24574 39922 24642 39978
rect 24698 39922 24768 39978
rect 24448 39888 24768 39922
rect 36138 40350 36758 57922
rect 55168 58350 55488 58384
rect 55168 58294 55238 58350
rect 55294 58294 55362 58350
rect 55418 58294 55488 58350
rect 55168 58226 55488 58294
rect 55168 58170 55238 58226
rect 55294 58170 55362 58226
rect 55418 58170 55488 58226
rect 55168 58102 55488 58170
rect 55168 58046 55238 58102
rect 55294 58046 55362 58102
rect 55418 58046 55488 58102
rect 55168 57978 55488 58046
rect 55168 57922 55238 57978
rect 55294 57922 55362 57978
rect 55418 57922 55488 57978
rect 55168 57888 55488 57922
rect 64652 51492 64708 70700
rect 64764 66388 64820 66398
rect 64764 52164 64820 66332
rect 64764 52098 64820 52108
rect 66858 58350 67478 75922
rect 66858 58294 66954 58350
rect 67010 58294 67078 58350
rect 67134 58294 67202 58350
rect 67258 58294 67326 58350
rect 67382 58294 67478 58350
rect 66858 58226 67478 58294
rect 66858 58170 66954 58226
rect 67010 58170 67078 58226
rect 67134 58170 67202 58226
rect 67258 58170 67326 58226
rect 67382 58170 67478 58226
rect 66858 58102 67478 58170
rect 66858 58046 66954 58102
rect 67010 58046 67078 58102
rect 67134 58046 67202 58102
rect 67258 58046 67326 58102
rect 67382 58046 67478 58102
rect 66858 57978 67478 58046
rect 66858 57922 66954 57978
rect 67010 57922 67078 57978
rect 67134 57922 67202 57978
rect 67258 57922 67326 57978
rect 67382 57922 67478 57978
rect 64652 51426 64708 51436
rect 64316 51380 64372 51390
rect 64092 51268 64148 51278
rect 64092 48132 64148 51212
rect 64316 48804 64372 51324
rect 64316 48738 64372 48748
rect 64092 48066 64148 48076
rect 64204 48692 64260 48702
rect 39808 46350 40128 46384
rect 39808 46294 39878 46350
rect 39934 46294 40002 46350
rect 40058 46294 40128 46350
rect 39808 46226 40128 46294
rect 39808 46170 39878 46226
rect 39934 46170 40002 46226
rect 40058 46170 40128 46226
rect 39808 46102 40128 46170
rect 39808 46046 39878 46102
rect 39934 46046 40002 46102
rect 40058 46046 40128 46102
rect 39808 45978 40128 46046
rect 39808 45922 39878 45978
rect 39934 45922 40002 45978
rect 40058 45922 40128 45978
rect 39808 45888 40128 45922
rect 64204 45444 64260 48636
rect 64204 45378 64260 45388
rect 36138 40294 36234 40350
rect 36290 40294 36358 40350
rect 36414 40294 36482 40350
rect 36538 40294 36606 40350
rect 36662 40294 36758 40350
rect 36138 40226 36758 40294
rect 36138 40170 36234 40226
rect 36290 40170 36358 40226
rect 36414 40170 36482 40226
rect 36538 40170 36606 40226
rect 36662 40170 36758 40226
rect 36138 40102 36758 40170
rect 36138 40046 36234 40102
rect 36290 40046 36358 40102
rect 36414 40046 36482 40102
rect 36538 40046 36606 40102
rect 36662 40046 36758 40102
rect 36138 39978 36758 40046
rect 36138 39922 36234 39978
rect 36290 39922 36358 39978
rect 36414 39922 36482 39978
rect 36538 39922 36606 39978
rect 36662 39922 36758 39978
rect 18396 5058 18452 5068
rect 36138 22350 36758 39922
rect 55168 40350 55488 40384
rect 55168 40294 55238 40350
rect 55294 40294 55362 40350
rect 55418 40294 55488 40350
rect 55168 40226 55488 40294
rect 55168 40170 55238 40226
rect 55294 40170 55362 40226
rect 55418 40170 55488 40226
rect 55168 40102 55488 40170
rect 55168 40046 55238 40102
rect 55294 40046 55362 40102
rect 55418 40046 55488 40102
rect 55168 39978 55488 40046
rect 55168 39922 55238 39978
rect 55294 39922 55362 39978
rect 55418 39922 55488 39978
rect 55168 39888 55488 39922
rect 66858 40350 67478 57922
rect 69692 96516 69748 96526
rect 69692 48692 69748 96460
rect 69692 48626 69748 48636
rect 69804 89908 69860 89918
rect 69804 44772 69860 89852
rect 69804 44706 69860 44716
rect 70578 82350 71198 99922
rect 82012 101108 82068 101118
rect 78092 98196 78148 98206
rect 70578 82294 70674 82350
rect 70730 82294 70798 82350
rect 70854 82294 70922 82350
rect 70978 82294 71046 82350
rect 71102 82294 71198 82350
rect 70578 82226 71198 82294
rect 70578 82170 70674 82226
rect 70730 82170 70798 82226
rect 70854 82170 70922 82226
rect 70978 82170 71046 82226
rect 71102 82170 71198 82226
rect 70578 82102 71198 82170
rect 70578 82046 70674 82102
rect 70730 82046 70798 82102
rect 70854 82046 70922 82102
rect 70978 82046 71046 82102
rect 71102 82046 71198 82102
rect 70578 81978 71198 82046
rect 70578 81922 70674 81978
rect 70730 81922 70798 81978
rect 70854 81922 70922 81978
rect 70978 81922 71046 81978
rect 71102 81922 71198 81978
rect 70578 64350 71198 81922
rect 70578 64294 70674 64350
rect 70730 64294 70798 64350
rect 70854 64294 70922 64350
rect 70978 64294 71046 64350
rect 71102 64294 71198 64350
rect 70578 64226 71198 64294
rect 70578 64170 70674 64226
rect 70730 64170 70798 64226
rect 70854 64170 70922 64226
rect 70978 64170 71046 64226
rect 71102 64170 71198 64226
rect 70578 64102 71198 64170
rect 70578 64046 70674 64102
rect 70730 64046 70798 64102
rect 70854 64046 70922 64102
rect 70978 64046 71046 64102
rect 71102 64046 71198 64102
rect 70578 63978 71198 64046
rect 70578 63922 70674 63978
rect 70730 63922 70798 63978
rect 70854 63922 70922 63978
rect 70978 63922 71046 63978
rect 71102 63922 71198 63978
rect 70578 46350 71198 63922
rect 73052 97076 73108 97086
rect 73052 51380 73108 97020
rect 74732 86548 74788 86558
rect 74732 52836 74788 86492
rect 76412 69076 76468 69086
rect 76412 66388 76468 69020
rect 76412 66322 76468 66332
rect 76524 68068 76580 68078
rect 76524 55468 76580 68012
rect 76412 55412 76580 55468
rect 76412 53508 76468 55412
rect 76412 53442 76468 53452
rect 74732 52770 74788 52780
rect 73052 51314 73108 51324
rect 78092 51268 78148 98140
rect 81452 91700 81508 91710
rect 78092 51202 78148 51212
rect 80220 77476 80276 77486
rect 70578 46294 70674 46350
rect 70730 46294 70798 46350
rect 70854 46294 70922 46350
rect 70978 46294 71046 46350
rect 71102 46294 71198 46350
rect 70578 46226 71198 46294
rect 70578 46170 70674 46226
rect 70730 46170 70798 46226
rect 70854 46170 70922 46226
rect 70978 46170 71046 46226
rect 71102 46170 71198 46226
rect 70578 46102 71198 46170
rect 70578 46046 70674 46102
rect 70730 46046 70798 46102
rect 70854 46046 70922 46102
rect 70978 46046 71046 46102
rect 71102 46046 71198 46102
rect 80220 46116 80276 77420
rect 80332 71428 80388 71438
rect 80332 54180 80388 71372
rect 80332 54114 80388 54124
rect 80444 68852 80500 68862
rect 80444 46788 80500 68796
rect 81452 50260 81508 91644
rect 81452 50194 81508 50204
rect 81564 72996 81620 73006
rect 81564 50148 81620 72940
rect 81564 50082 81620 50092
rect 82012 47460 82068 101052
rect 97578 94350 98198 111922
rect 117168 112350 117488 112384
rect 117168 112294 117238 112350
rect 117294 112294 117362 112350
rect 117418 112294 117488 112350
rect 117168 112226 117488 112294
rect 117168 112170 117238 112226
rect 117294 112170 117362 112226
rect 117418 112170 117488 112226
rect 117168 112102 117488 112170
rect 117168 112046 117238 112102
rect 117294 112046 117362 112102
rect 117418 112046 117488 112102
rect 117168 111978 117488 112046
rect 117168 111922 117238 111978
rect 117294 111922 117362 111978
rect 117418 111922 117488 111978
rect 117168 111888 117488 111922
rect 128298 112350 128918 129922
rect 128298 112294 128394 112350
rect 128450 112294 128518 112350
rect 128574 112294 128642 112350
rect 128698 112294 128766 112350
rect 128822 112294 128918 112350
rect 128298 112226 128918 112294
rect 128298 112170 128394 112226
rect 128450 112170 128518 112226
rect 128574 112170 128642 112226
rect 128698 112170 128766 112226
rect 128822 112170 128918 112226
rect 128298 112102 128918 112170
rect 128298 112046 128394 112102
rect 128450 112046 128518 112102
rect 128574 112046 128642 112102
rect 128698 112046 128766 112102
rect 128822 112046 128918 112102
rect 128298 111978 128918 112046
rect 128298 111922 128394 111978
rect 128450 111922 128518 111978
rect 128574 111922 128642 111978
rect 128698 111922 128766 111978
rect 128822 111922 128918 111978
rect 102844 101668 102900 101678
rect 97578 94294 97674 94350
rect 97730 94294 97798 94350
rect 97854 94294 97922 94350
rect 97978 94294 98046 94350
rect 98102 94294 98198 94350
rect 97578 94226 98198 94294
rect 97578 94170 97674 94226
rect 97730 94170 97798 94226
rect 97854 94170 97922 94226
rect 97978 94170 98046 94226
rect 98102 94170 98198 94226
rect 97578 94102 98198 94170
rect 97578 94046 97674 94102
rect 97730 94046 97798 94102
rect 97854 94046 97922 94102
rect 97978 94046 98046 94102
rect 98102 94046 98198 94102
rect 97578 93978 98198 94046
rect 97578 93922 97674 93978
rect 97730 93922 97798 93978
rect 97854 93922 97922 93978
rect 97978 93922 98046 93978
rect 98102 93922 98198 93978
rect 97578 76350 98198 93922
rect 97578 76294 97674 76350
rect 97730 76294 97798 76350
rect 97854 76294 97922 76350
rect 97978 76294 98046 76350
rect 98102 76294 98198 76350
rect 97578 76226 98198 76294
rect 97578 76170 97674 76226
rect 97730 76170 97798 76226
rect 97854 76170 97922 76226
rect 97978 76170 98046 76226
rect 98102 76170 98198 76226
rect 97578 76102 98198 76170
rect 97578 76046 97674 76102
rect 97730 76046 97798 76102
rect 97854 76046 97922 76102
rect 97978 76046 98046 76102
rect 98102 76046 98198 76102
rect 97578 75978 98198 76046
rect 97578 75922 97674 75978
rect 97730 75922 97798 75978
rect 97854 75922 97922 75978
rect 97978 75922 98046 75978
rect 98102 75922 98198 75978
rect 82348 75236 82404 75246
rect 82348 68852 82404 75180
rect 82348 68786 82404 68796
rect 86448 58350 86768 58384
rect 86448 58294 86518 58350
rect 86574 58294 86642 58350
rect 86698 58294 86768 58350
rect 86448 58226 86768 58294
rect 86448 58170 86518 58226
rect 86574 58170 86642 58226
rect 86698 58170 86768 58226
rect 86448 58102 86768 58170
rect 86448 58046 86518 58102
rect 86574 58046 86642 58102
rect 86698 58046 86768 58102
rect 86448 57978 86768 58046
rect 86448 57922 86518 57978
rect 86574 57922 86642 57978
rect 86698 57922 86768 57978
rect 86448 57888 86768 57922
rect 97578 58350 98198 75922
rect 101298 100350 101918 101364
rect 102844 100772 102900 101612
rect 102844 100706 102900 100716
rect 101298 100294 101394 100350
rect 101450 100294 101518 100350
rect 101574 100294 101642 100350
rect 101698 100294 101766 100350
rect 101822 100294 101918 100350
rect 101298 100226 101918 100294
rect 101298 100170 101394 100226
rect 101450 100170 101518 100226
rect 101574 100170 101642 100226
rect 101698 100170 101766 100226
rect 101822 100170 101918 100226
rect 101298 100102 101918 100170
rect 101298 100046 101394 100102
rect 101450 100046 101518 100102
rect 101574 100046 101642 100102
rect 101698 100046 101766 100102
rect 101822 100046 101918 100102
rect 101298 99978 101918 100046
rect 101298 99922 101394 99978
rect 101450 99922 101518 99978
rect 101574 99922 101642 99978
rect 101698 99922 101766 99978
rect 101822 99922 101918 99978
rect 101298 82350 101918 99922
rect 128298 94350 128918 111922
rect 128298 94294 128394 94350
rect 128450 94294 128518 94350
rect 128574 94294 128642 94350
rect 128698 94294 128766 94350
rect 128822 94294 128918 94350
rect 128298 94226 128918 94294
rect 128298 94170 128394 94226
rect 128450 94170 128518 94226
rect 128574 94170 128642 94226
rect 128698 94170 128766 94226
rect 128822 94170 128918 94226
rect 128298 94102 128918 94170
rect 128298 94046 128394 94102
rect 128450 94046 128518 94102
rect 128574 94046 128642 94102
rect 128698 94046 128766 94102
rect 128822 94046 128918 94102
rect 128298 93978 128918 94046
rect 128298 93922 128394 93978
rect 128450 93922 128518 93978
rect 128574 93922 128642 93978
rect 128698 93922 128766 93978
rect 128822 93922 128918 93978
rect 101298 82294 101394 82350
rect 101450 82294 101518 82350
rect 101574 82294 101642 82350
rect 101698 82294 101766 82350
rect 101822 82294 101918 82350
rect 101298 82226 101918 82294
rect 101298 82170 101394 82226
rect 101450 82170 101518 82226
rect 101574 82170 101642 82226
rect 101698 82170 101766 82226
rect 101822 82170 101918 82226
rect 101298 82102 101918 82170
rect 101298 82046 101394 82102
rect 101450 82046 101518 82102
rect 101574 82046 101642 82102
rect 101698 82046 101766 82102
rect 101822 82046 101918 82102
rect 101298 81978 101918 82046
rect 101298 81922 101394 81978
rect 101450 81922 101518 81978
rect 101574 81922 101642 81978
rect 101698 81922 101766 81978
rect 101822 81922 101918 81978
rect 101298 69788 101918 81922
rect 126812 84868 126868 84878
rect 101808 64350 102128 64384
rect 101808 64294 101878 64350
rect 101934 64294 102002 64350
rect 102058 64294 102128 64350
rect 101808 64226 102128 64294
rect 101808 64170 101878 64226
rect 101934 64170 102002 64226
rect 102058 64170 102128 64226
rect 101808 64102 102128 64170
rect 101808 64046 101878 64102
rect 101934 64046 102002 64102
rect 102058 64046 102128 64102
rect 101808 63978 102128 64046
rect 101808 63922 101878 63978
rect 101934 63922 102002 63978
rect 102058 63922 102128 63978
rect 101808 63888 102128 63922
rect 97578 58294 97674 58350
rect 97730 58294 97798 58350
rect 97854 58294 97922 58350
rect 97978 58294 98046 58350
rect 98102 58294 98198 58350
rect 97578 58226 98198 58294
rect 97578 58170 97674 58226
rect 97730 58170 97798 58226
rect 97854 58170 97922 58226
rect 97978 58170 98046 58226
rect 98102 58170 98198 58226
rect 97578 58102 98198 58170
rect 97578 58046 97674 58102
rect 97730 58046 97798 58102
rect 97854 58046 97922 58102
rect 97978 58046 98046 58102
rect 98102 58046 98198 58102
rect 97578 57978 98198 58046
rect 97578 57922 97674 57978
rect 97730 57922 97798 57978
rect 97854 57922 97922 57978
rect 97978 57922 98046 57978
rect 98102 57922 98198 57978
rect 82572 56308 82628 56318
rect 82684 56278 82740 56288
rect 82628 56252 82684 56278
rect 82572 56222 82684 56252
rect 82684 56212 82740 56222
rect 97578 50558 98198 57922
rect 117168 58350 117488 58384
rect 117168 58294 117238 58350
rect 117294 58294 117362 58350
rect 117418 58294 117488 58350
rect 117168 58226 117488 58294
rect 117168 58170 117238 58226
rect 117294 58170 117362 58226
rect 117418 58170 117488 58226
rect 117168 58102 117488 58170
rect 117168 58046 117238 58102
rect 117294 58046 117362 58102
rect 117418 58046 117488 58102
rect 117168 57978 117488 58046
rect 117168 57922 117238 57978
rect 117294 57922 117362 57978
rect 117418 57922 117488 57978
rect 117168 57888 117488 57922
rect 126812 50820 126868 84812
rect 128298 76350 128918 93922
rect 132018 208350 132638 225922
rect 132018 208294 132114 208350
rect 132170 208294 132238 208350
rect 132294 208294 132362 208350
rect 132418 208294 132486 208350
rect 132542 208294 132638 208350
rect 132018 208226 132638 208294
rect 132018 208170 132114 208226
rect 132170 208170 132238 208226
rect 132294 208170 132362 208226
rect 132418 208170 132486 208226
rect 132542 208170 132638 208226
rect 132018 208102 132638 208170
rect 132018 208046 132114 208102
rect 132170 208046 132238 208102
rect 132294 208046 132362 208102
rect 132418 208046 132486 208102
rect 132542 208046 132638 208102
rect 132018 207978 132638 208046
rect 132018 207922 132114 207978
rect 132170 207922 132238 207978
rect 132294 207922 132362 207978
rect 132418 207922 132486 207978
rect 132542 207922 132638 207978
rect 132018 190350 132638 207922
rect 140588 232596 140644 232606
rect 132018 190294 132114 190350
rect 132170 190294 132238 190350
rect 132294 190294 132362 190350
rect 132418 190294 132486 190350
rect 132542 190294 132638 190350
rect 132018 190226 132638 190294
rect 132018 190170 132114 190226
rect 132170 190170 132238 190226
rect 132294 190170 132362 190226
rect 132418 190170 132486 190226
rect 132542 190170 132638 190226
rect 132018 190102 132638 190170
rect 132018 190046 132114 190102
rect 132170 190046 132238 190102
rect 132294 190046 132362 190102
rect 132418 190046 132486 190102
rect 132542 190046 132638 190102
rect 132018 189978 132638 190046
rect 132018 189922 132114 189978
rect 132170 189922 132238 189978
rect 132294 189922 132362 189978
rect 132418 189922 132486 189978
rect 132542 189922 132638 189978
rect 132018 172350 132638 189922
rect 134428 192178 134484 192188
rect 134428 188468 134484 192122
rect 134428 188402 134484 188412
rect 140588 187796 140644 232540
rect 140700 231476 140756 231486
rect 140700 198548 140756 231420
rect 140700 198482 140756 198492
rect 140812 230356 140868 230366
rect 140812 192500 140868 230300
rect 140812 192434 140868 192444
rect 140924 229796 140980 229806
rect 140924 188468 140980 229740
rect 144060 224308 144116 224318
rect 144060 208628 144116 224252
rect 144060 208562 144116 208572
rect 159018 220350 159638 237922
rect 159018 220294 159114 220350
rect 159170 220294 159238 220350
rect 159294 220294 159362 220350
rect 159418 220294 159486 220350
rect 159542 220294 159638 220350
rect 159018 220226 159638 220294
rect 159018 220170 159114 220226
rect 159170 220170 159238 220226
rect 159294 220170 159362 220226
rect 159418 220170 159486 220226
rect 159542 220170 159638 220226
rect 159018 220102 159638 220170
rect 159018 220046 159114 220102
rect 159170 220046 159238 220102
rect 159294 220046 159362 220102
rect 159418 220046 159486 220102
rect 159542 220046 159638 220102
rect 159018 219978 159638 220046
rect 159018 219922 159114 219978
rect 159170 219922 159238 219978
rect 159294 219922 159362 219978
rect 159418 219922 159486 219978
rect 159542 219922 159638 219978
rect 148448 202350 148768 202384
rect 148448 202294 148518 202350
rect 148574 202294 148642 202350
rect 148698 202294 148768 202350
rect 148448 202226 148768 202294
rect 148448 202170 148518 202226
rect 148574 202170 148642 202226
rect 148698 202170 148768 202226
rect 148448 202102 148768 202170
rect 148448 202046 148518 202102
rect 148574 202046 148642 202102
rect 148698 202046 148768 202102
rect 148448 201978 148768 202046
rect 148448 201922 148518 201978
rect 148574 201922 148642 201978
rect 148698 201922 148768 201978
rect 148448 201888 148768 201922
rect 159018 202350 159638 219922
rect 162738 262052 163358 262098
rect 162738 261996 162834 262052
rect 162890 261996 162958 262052
rect 163014 261996 163082 262052
rect 163138 261996 163206 262052
rect 163262 261996 163358 262052
rect 162738 261928 163358 261996
rect 162738 261872 162834 261928
rect 162890 261872 162958 261928
rect 163014 261872 163082 261928
rect 163138 261872 163206 261928
rect 163262 261872 163358 261928
rect 163808 262046 163878 262102
rect 163934 262046 164002 262102
rect 164058 262046 164128 262102
rect 163808 261978 164128 262046
rect 163808 261922 163878 261978
rect 163934 261922 164002 261978
rect 164058 261922 164128 261978
rect 163808 261888 164128 261922
rect 162738 244350 163358 261872
rect 188972 259028 189028 289100
rect 189196 263732 189252 290220
rect 189738 274350 190358 291922
rect 189738 274294 189834 274350
rect 189890 274294 189958 274350
rect 190014 274294 190082 274350
rect 190138 274294 190206 274350
rect 190262 274294 190358 274350
rect 189738 274226 190358 274294
rect 189738 274170 189834 274226
rect 189890 274170 189958 274226
rect 190014 274170 190082 274226
rect 190138 274170 190206 274226
rect 190262 274170 190358 274226
rect 189738 274102 190358 274170
rect 189738 274046 189834 274102
rect 189890 274046 189958 274102
rect 190014 274046 190082 274102
rect 190138 274046 190206 274102
rect 190262 274046 190358 274102
rect 189738 273978 190358 274046
rect 189738 273922 189834 273978
rect 189890 273922 189958 273978
rect 190014 273922 190082 273978
rect 190138 273922 190206 273978
rect 190262 273922 190358 273978
rect 189532 268436 189588 268446
rect 189532 266644 189588 268380
rect 189532 266578 189588 266588
rect 189532 266420 189588 266430
rect 189532 264898 189588 266364
rect 189532 264832 189588 264842
rect 189196 263666 189252 263676
rect 188972 258962 189028 258972
rect 179168 256350 179488 256384
rect 179168 256294 179238 256350
rect 179294 256294 179362 256350
rect 179418 256294 179488 256350
rect 179168 256226 179488 256294
rect 179168 256170 179238 256226
rect 179294 256170 179362 256226
rect 179418 256170 179488 256226
rect 179168 256102 179488 256170
rect 179168 256046 179238 256102
rect 179294 256046 179362 256102
rect 179418 256046 179488 256102
rect 179168 255978 179488 256046
rect 179168 255922 179238 255978
rect 179294 255922 179362 255978
rect 179418 255922 179488 255978
rect 179168 255888 179488 255922
rect 189738 256350 190358 273922
rect 189738 256294 189834 256350
rect 189890 256294 189958 256350
rect 190014 256294 190082 256350
rect 190138 256294 190206 256350
rect 190262 256294 190358 256350
rect 189738 256226 190358 256294
rect 189738 256170 189834 256226
rect 189890 256170 189958 256226
rect 190014 256170 190082 256226
rect 190138 256170 190206 256226
rect 190262 256170 190358 256226
rect 189738 256102 190358 256170
rect 189738 256046 189834 256102
rect 189890 256046 189958 256102
rect 190014 256046 190082 256102
rect 190138 256046 190206 256102
rect 190262 256046 190358 256102
rect 189738 255978 190358 256046
rect 189738 255922 189834 255978
rect 189890 255922 189958 255978
rect 190014 255922 190082 255978
rect 190138 255922 190206 255978
rect 190262 255922 190358 255978
rect 162738 244294 162834 244350
rect 162890 244294 162958 244350
rect 163014 244294 163082 244350
rect 163138 244294 163206 244350
rect 163262 244294 163358 244350
rect 162738 244226 163358 244294
rect 162738 244170 162834 244226
rect 162890 244170 162958 244226
rect 163014 244170 163082 244226
rect 163138 244170 163206 244226
rect 163262 244170 163358 244226
rect 162738 244102 163358 244170
rect 162738 244046 162834 244102
rect 162890 244046 162958 244102
rect 163014 244046 163082 244102
rect 163138 244046 163206 244102
rect 163262 244046 163358 244102
rect 162738 243978 163358 244046
rect 162738 243922 162834 243978
rect 162890 243922 162958 243978
rect 163014 243922 163082 243978
rect 163138 243922 163206 243978
rect 163262 243922 163358 243978
rect 162738 226350 163358 243922
rect 189738 238350 190358 255922
rect 189738 238294 189834 238350
rect 189890 238294 189958 238350
rect 190014 238294 190082 238350
rect 190138 238294 190206 238350
rect 190262 238294 190358 238350
rect 189738 238226 190358 238294
rect 189738 238170 189834 238226
rect 189890 238170 189958 238226
rect 190014 238170 190082 238226
rect 190138 238170 190206 238226
rect 190262 238170 190358 238226
rect 189738 238102 190358 238170
rect 189738 238046 189834 238102
rect 189890 238046 189958 238102
rect 190014 238046 190082 238102
rect 190138 238046 190206 238102
rect 190262 238046 190358 238102
rect 189738 237978 190358 238046
rect 189738 237922 189834 237978
rect 189890 237922 189958 237978
rect 190014 237922 190082 237978
rect 190138 237922 190206 237978
rect 190262 237922 190358 237978
rect 189196 228116 189252 228126
rect 162738 226294 162834 226350
rect 162890 226294 162958 226350
rect 163014 226294 163082 226350
rect 163138 226294 163206 226350
rect 163262 226294 163358 226350
rect 162738 226226 163358 226294
rect 162738 226170 162834 226226
rect 162890 226170 162958 226226
rect 163014 226170 163082 226226
rect 163138 226170 163206 226226
rect 163262 226170 163358 226226
rect 162738 226102 163358 226170
rect 162738 226046 162834 226102
rect 162890 226046 162958 226102
rect 163014 226046 163082 226102
rect 163138 226046 163206 226102
rect 163262 226046 163358 226102
rect 162738 225978 163358 226046
rect 162738 225922 162834 225978
rect 162890 225922 162958 225978
rect 163014 225922 163082 225978
rect 163138 225922 163206 225978
rect 163262 225922 163358 225978
rect 160188 212884 160244 212894
rect 160188 212660 160244 212828
rect 160188 212594 160244 212604
rect 159018 202294 159114 202350
rect 159170 202294 159238 202350
rect 159294 202294 159362 202350
rect 159418 202294 159486 202350
rect 159542 202294 159638 202350
rect 159018 202226 159638 202294
rect 159018 202170 159114 202226
rect 159170 202170 159238 202226
rect 159294 202170 159362 202226
rect 159418 202170 159486 202226
rect 159542 202170 159638 202226
rect 159018 202102 159638 202170
rect 159018 202046 159114 202102
rect 159170 202046 159238 202102
rect 159294 202046 159362 202102
rect 159418 202046 159486 202102
rect 159542 202046 159638 202102
rect 159018 201978 159638 202046
rect 159018 201922 159114 201978
rect 159170 201922 159238 201978
rect 159294 201922 159362 201978
rect 159418 201922 159486 201978
rect 159542 201922 159638 201978
rect 141036 199892 141092 199902
rect 141036 199018 141092 199836
rect 141036 198952 141092 198962
rect 140924 188402 140980 188412
rect 140588 187730 140644 187740
rect 148448 184350 148768 184384
rect 148448 184294 148518 184350
rect 148574 184294 148642 184350
rect 148698 184294 148768 184350
rect 148448 184226 148768 184294
rect 148448 184170 148518 184226
rect 148574 184170 148642 184226
rect 148698 184170 148768 184226
rect 148448 184102 148768 184170
rect 148448 184046 148518 184102
rect 148574 184046 148642 184102
rect 148698 184046 148768 184102
rect 148448 183978 148768 184046
rect 148448 183922 148518 183978
rect 148574 183922 148642 183978
rect 148698 183922 148768 183978
rect 148448 183888 148768 183922
rect 159018 184350 159638 201922
rect 162738 208350 163358 225922
rect 188972 227556 189028 227566
rect 162738 208294 162834 208350
rect 162890 208294 162958 208350
rect 163014 208294 163082 208350
rect 163138 208294 163206 208350
rect 163262 208294 163358 208350
rect 162738 208226 163358 208294
rect 162738 208170 162834 208226
rect 162890 208170 162958 208226
rect 163014 208170 163082 208226
rect 163138 208170 163206 208226
rect 163262 208170 163358 208226
rect 162738 208102 163358 208170
rect 162738 208046 162834 208102
rect 162890 208046 162958 208102
rect 163014 208046 163082 208102
rect 163138 208046 163206 208102
rect 163262 208046 163358 208102
rect 162738 207978 163358 208046
rect 162738 207922 162834 207978
rect 162890 207922 162958 207978
rect 163014 207922 163082 207978
rect 163138 207922 163206 207978
rect 163262 207922 163358 207978
rect 162738 193966 163358 207922
rect 163808 208350 164128 208384
rect 163808 208294 163878 208350
rect 163934 208294 164002 208350
rect 164058 208294 164128 208350
rect 163808 208226 164128 208294
rect 163808 208170 163878 208226
rect 163934 208170 164002 208226
rect 164058 208170 164128 208226
rect 163808 208102 164128 208170
rect 163808 208046 163878 208102
rect 163934 208046 164002 208102
rect 164058 208046 164128 208102
rect 163808 207978 164128 208046
rect 163808 207922 163878 207978
rect 163934 207922 164002 207978
rect 164058 207922 164128 207978
rect 163808 207888 164128 207922
rect 179168 202350 179488 202384
rect 179168 202294 179238 202350
rect 179294 202294 179362 202350
rect 179418 202294 179488 202350
rect 179168 202226 179488 202294
rect 179168 202170 179238 202226
rect 179294 202170 179362 202226
rect 179418 202170 179488 202226
rect 179168 202102 179488 202170
rect 179168 202046 179238 202102
rect 179294 202046 179362 202102
rect 179418 202046 179488 202102
rect 179168 201978 179488 202046
rect 179168 201922 179238 201978
rect 179294 201922 179362 201978
rect 179418 201922 179488 201978
rect 179168 201888 179488 201922
rect 187292 196678 187348 196688
rect 169708 193978 169764 193988
rect 163808 190350 164128 190384
rect 163808 190294 163878 190350
rect 163934 190294 164002 190350
rect 164058 190294 164128 190350
rect 163808 190226 164128 190294
rect 163808 190170 163878 190226
rect 163934 190170 164002 190226
rect 164058 190170 164128 190226
rect 163808 190102 164128 190170
rect 163808 190046 163878 190102
rect 163934 190046 164002 190102
rect 164058 190046 164128 190102
rect 163808 189978 164128 190046
rect 163808 189922 163878 189978
rect 163934 189922 164002 189978
rect 164058 189922 164128 189978
rect 163808 189888 164128 189922
rect 169708 189658 169764 193922
rect 169708 189592 169764 189602
rect 187292 187498 187348 196622
rect 188076 195238 188132 195248
rect 188076 189478 188132 195182
rect 188972 193172 189028 227500
rect 189196 195188 189252 228060
rect 189738 220350 190358 237922
rect 193458 316350 194078 333922
rect 197372 328916 197428 347822
rect 197372 328850 197428 328860
rect 193458 316294 193554 316350
rect 193610 316294 193678 316350
rect 193734 316294 193802 316350
rect 193858 316294 193926 316350
rect 193982 316294 194078 316350
rect 193458 316226 194078 316294
rect 193458 316170 193554 316226
rect 193610 316170 193678 316226
rect 193734 316170 193802 316226
rect 193858 316170 193926 316226
rect 193982 316170 194078 316226
rect 193458 316102 194078 316170
rect 193458 316046 193554 316102
rect 193610 316046 193678 316102
rect 193734 316046 193802 316102
rect 193858 316046 193926 316102
rect 193982 316046 194078 316102
rect 193458 315978 194078 316046
rect 193458 315922 193554 315978
rect 193610 315922 193678 315978
rect 193734 315922 193802 315978
rect 193858 315922 193926 315978
rect 193982 315922 194078 315978
rect 193458 298350 194078 315922
rect 198156 313348 198212 313358
rect 198156 309316 198212 313292
rect 198156 309250 198212 309260
rect 193458 298294 193554 298350
rect 193610 298294 193678 298350
rect 193734 298294 193802 298350
rect 193858 298294 193926 298350
rect 193982 298294 194078 298350
rect 193458 298226 194078 298294
rect 193458 298170 193554 298226
rect 193610 298170 193678 298226
rect 193734 298170 193802 298226
rect 193858 298170 193926 298226
rect 193982 298170 194078 298226
rect 193458 298102 194078 298170
rect 193458 298046 193554 298102
rect 193610 298046 193678 298102
rect 193734 298046 193802 298102
rect 193858 298046 193926 298102
rect 193982 298046 194078 298102
rect 193458 297978 194078 298046
rect 193458 297922 193554 297978
rect 193610 297922 193678 297978
rect 193734 297922 193802 297978
rect 193858 297922 193926 297978
rect 193982 297922 194078 297978
rect 193458 280350 194078 297922
rect 193458 280294 193554 280350
rect 193610 280294 193678 280350
rect 193734 280294 193802 280350
rect 193858 280294 193926 280350
rect 193982 280294 194078 280350
rect 193458 280226 194078 280294
rect 193458 280170 193554 280226
rect 193610 280170 193678 280226
rect 193734 280170 193802 280226
rect 193858 280170 193926 280226
rect 193982 280170 194078 280226
rect 193458 280102 194078 280170
rect 193458 280046 193554 280102
rect 193610 280046 193678 280102
rect 193734 280046 193802 280102
rect 193858 280046 193926 280102
rect 193982 280046 194078 280102
rect 193458 279978 194078 280046
rect 193458 279922 193554 279978
rect 193610 279922 193678 279978
rect 193734 279922 193802 279978
rect 193858 279922 193926 279978
rect 193982 279922 194078 279978
rect 193458 262350 194078 279922
rect 200732 288036 200788 288046
rect 195692 278218 195748 278228
rect 194908 271558 194964 271568
rect 194908 270118 194964 271502
rect 194908 270052 194964 270062
rect 195692 267058 195748 278162
rect 195692 266992 195748 267002
rect 198268 268858 198324 268868
rect 198268 264538 198324 268802
rect 198268 264472 198324 264482
rect 199836 266644 199892 266654
rect 193458 262294 193554 262350
rect 193610 262294 193678 262350
rect 193734 262294 193802 262350
rect 193858 262294 193926 262350
rect 193982 262294 194078 262350
rect 193458 262226 194078 262294
rect 193458 262170 193554 262226
rect 193610 262170 193678 262226
rect 193734 262170 193802 262226
rect 193858 262170 193926 262226
rect 193982 262170 194078 262226
rect 193458 262102 194078 262170
rect 193458 262046 193554 262102
rect 193610 262046 193678 262102
rect 193734 262046 193802 262102
rect 193858 262046 193926 262102
rect 193982 262046 194078 262102
rect 193458 261978 194078 262046
rect 193458 261922 193554 261978
rect 193610 261922 193678 261978
rect 193734 261922 193802 261978
rect 193858 261922 193926 261978
rect 193982 261922 194078 261978
rect 193458 244350 194078 261922
rect 194908 262052 194964 262062
rect 194908 258418 194964 261996
rect 199836 260218 199892 266588
rect 200732 260372 200788 287980
rect 200732 260306 200788 260316
rect 199836 260152 199892 260162
rect 194908 258352 194964 258362
rect 193458 244294 193554 244350
rect 193610 244294 193678 244350
rect 193734 244294 193802 244350
rect 193858 244294 193926 244350
rect 193982 244294 194078 244350
rect 193458 244226 194078 244294
rect 193458 244170 193554 244226
rect 193610 244170 193678 244226
rect 193734 244170 193802 244226
rect 193858 244170 193926 244226
rect 193982 244170 194078 244226
rect 193458 244102 194078 244170
rect 193458 244046 193554 244102
rect 193610 244046 193678 244102
rect 193734 244046 193802 244102
rect 193858 244046 193926 244102
rect 193982 244046 194078 244102
rect 193458 243978 194078 244046
rect 193458 243922 193554 243978
rect 193610 243922 193678 243978
rect 193734 243922 193802 243978
rect 193858 243922 193926 243978
rect 193982 243922 194078 243978
rect 193458 226350 194078 243922
rect 193458 226294 193554 226350
rect 193610 226294 193678 226350
rect 193734 226294 193802 226350
rect 193858 226294 193926 226350
rect 193982 226294 194078 226350
rect 193458 226226 194078 226294
rect 193458 226170 193554 226226
rect 193610 226170 193678 226226
rect 193734 226170 193802 226226
rect 193858 226170 193926 226226
rect 193982 226170 194078 226226
rect 193458 226102 194078 226170
rect 193458 226046 193554 226102
rect 193610 226046 193678 226102
rect 193734 226046 193802 226102
rect 193858 226046 193926 226102
rect 193982 226046 194078 226102
rect 193458 225978 194078 226046
rect 193458 225922 193554 225978
rect 193610 225922 193678 225978
rect 193734 225922 193802 225978
rect 193858 225922 193926 225978
rect 193982 225922 194078 225978
rect 189738 220294 189834 220350
rect 189890 220294 189958 220350
rect 190014 220294 190082 220350
rect 190138 220294 190206 220350
rect 190262 220294 190358 220350
rect 189738 220226 190358 220294
rect 189738 220170 189834 220226
rect 189890 220170 189958 220226
rect 190014 220170 190082 220226
rect 190138 220170 190206 220226
rect 190262 220170 190358 220226
rect 189738 220102 190358 220170
rect 189738 220046 189834 220102
rect 189890 220046 189958 220102
rect 190014 220046 190082 220102
rect 190138 220046 190206 220102
rect 190262 220046 190358 220102
rect 189738 219978 190358 220046
rect 189738 219922 189834 219978
rect 189890 219922 189958 219978
rect 190014 219922 190082 219978
rect 190138 219922 190206 219978
rect 190262 219922 190358 219978
rect 189738 202350 190358 219922
rect 189738 202294 189834 202350
rect 189890 202294 189958 202350
rect 190014 202294 190082 202350
rect 190138 202294 190206 202350
rect 190262 202294 190358 202350
rect 189738 202226 190358 202294
rect 189738 202170 189834 202226
rect 189890 202170 189958 202226
rect 190014 202170 190082 202226
rect 190138 202170 190206 202226
rect 190262 202170 190358 202226
rect 189738 202102 190358 202170
rect 189738 202046 189834 202102
rect 189890 202046 189958 202102
rect 190014 202046 190082 202102
rect 190138 202046 190206 202102
rect 190262 202046 190358 202102
rect 189738 201978 190358 202046
rect 189738 201922 189834 201978
rect 189890 201922 189958 201978
rect 190014 201922 190082 201978
rect 190138 201922 190206 201978
rect 190262 201922 190358 201978
rect 189532 196498 189588 196508
rect 189532 195860 189588 196442
rect 189532 195794 189588 195804
rect 189196 195122 189252 195132
rect 188972 193106 189028 193116
rect 189532 192388 189588 192398
rect 189532 189812 189588 192332
rect 189532 189746 189588 189756
rect 188076 189412 188132 189422
rect 187292 187432 187348 187442
rect 169708 187318 169764 187328
rect 169708 186058 169764 187262
rect 169708 185992 169764 186002
rect 159018 184294 159114 184350
rect 159170 184294 159238 184350
rect 159294 184294 159362 184350
rect 159418 184294 159486 184350
rect 159542 184294 159638 184350
rect 159018 184226 159638 184294
rect 159018 184170 159114 184226
rect 159170 184170 159238 184226
rect 159294 184170 159362 184226
rect 159418 184170 159486 184226
rect 159542 184170 159638 184226
rect 159018 184102 159638 184170
rect 159018 184046 159114 184102
rect 159170 184046 159238 184102
rect 159294 184046 159362 184102
rect 159418 184046 159486 184102
rect 159542 184046 159638 184102
rect 159018 183978 159638 184046
rect 159018 183922 159114 183978
rect 159170 183922 159238 183978
rect 159294 183922 159362 183978
rect 159418 183922 159486 183978
rect 159542 183922 159638 183978
rect 132018 172294 132114 172350
rect 132170 172294 132238 172350
rect 132294 172294 132362 172350
rect 132418 172294 132486 172350
rect 132542 172294 132638 172350
rect 132018 172226 132638 172294
rect 132018 172170 132114 172226
rect 132170 172170 132238 172226
rect 132294 172170 132362 172226
rect 132418 172170 132486 172226
rect 132542 172170 132638 172226
rect 132018 172102 132638 172170
rect 132018 172046 132114 172102
rect 132170 172046 132238 172102
rect 132294 172046 132362 172102
rect 132418 172046 132486 172102
rect 132542 172046 132638 172102
rect 132018 171978 132638 172046
rect 132018 171922 132114 171978
rect 132170 171922 132238 171978
rect 132294 171922 132362 171978
rect 132418 171922 132486 171978
rect 132542 171922 132638 171978
rect 132018 154350 132638 171922
rect 132018 154294 132114 154350
rect 132170 154294 132238 154350
rect 132294 154294 132362 154350
rect 132418 154294 132486 154350
rect 132542 154294 132638 154350
rect 132018 154226 132638 154294
rect 132018 154170 132114 154226
rect 132170 154170 132238 154226
rect 132294 154170 132362 154226
rect 132418 154170 132486 154226
rect 132542 154170 132638 154226
rect 132018 154102 132638 154170
rect 132018 154046 132114 154102
rect 132170 154046 132238 154102
rect 132294 154046 132362 154102
rect 132418 154046 132486 154102
rect 132542 154046 132638 154102
rect 132018 153978 132638 154046
rect 132018 153922 132114 153978
rect 132170 153922 132238 153978
rect 132294 153922 132362 153978
rect 132418 153922 132486 153978
rect 132542 153922 132638 153978
rect 132018 136350 132638 153922
rect 140812 173796 140868 173806
rect 132018 136294 132114 136350
rect 132170 136294 132238 136350
rect 132294 136294 132362 136350
rect 132418 136294 132486 136350
rect 132542 136294 132638 136350
rect 132018 136226 132638 136294
rect 132018 136170 132114 136226
rect 132170 136170 132238 136226
rect 132294 136170 132362 136226
rect 132418 136170 132486 136226
rect 132542 136170 132638 136226
rect 132018 136102 132638 136170
rect 132018 136046 132114 136102
rect 132170 136046 132238 136102
rect 132294 136046 132362 136102
rect 132418 136046 132486 136102
rect 132542 136046 132638 136102
rect 132018 135978 132638 136046
rect 132018 135922 132114 135978
rect 132170 135922 132238 135978
rect 132294 135922 132362 135978
rect 132418 135922 132486 135978
rect 132542 135922 132638 135978
rect 132018 118350 132638 135922
rect 136892 139748 136948 139758
rect 136892 118580 136948 139692
rect 138572 132958 138628 132968
rect 138572 125938 138628 132902
rect 138572 125872 138628 125882
rect 140812 124628 140868 173740
rect 159018 166350 159638 183922
rect 159018 166294 159114 166350
rect 159170 166294 159238 166350
rect 159294 166294 159362 166350
rect 159418 166294 159486 166350
rect 159542 166294 159638 166350
rect 159018 166226 159638 166294
rect 159018 166170 159114 166226
rect 159170 166170 159238 166226
rect 159294 166170 159362 166226
rect 159418 166170 159486 166226
rect 159542 166170 159638 166226
rect 159018 166102 159638 166170
rect 159018 166046 159114 166102
rect 159170 166046 159238 166102
rect 159294 166046 159362 166102
rect 159418 166046 159486 166102
rect 159542 166046 159638 166102
rect 159018 165978 159638 166046
rect 159018 165922 159114 165978
rect 159170 165922 159238 165978
rect 159294 165922 159362 165978
rect 159418 165922 159486 165978
rect 159542 165922 159638 165978
rect 159018 148350 159638 165922
rect 159018 148294 159114 148350
rect 159170 148294 159238 148350
rect 159294 148294 159362 148350
rect 159418 148294 159486 148350
rect 159542 148294 159638 148350
rect 159018 148226 159638 148294
rect 159018 148170 159114 148226
rect 159170 148170 159238 148226
rect 159294 148170 159362 148226
rect 159418 148170 159486 148226
rect 159542 148170 159638 148226
rect 159018 148102 159638 148170
rect 159018 148046 159114 148102
rect 159170 148046 159238 148102
rect 159294 148046 159362 148102
rect 159418 148046 159486 148102
rect 159542 148046 159638 148102
rect 159018 147978 159638 148046
rect 159018 147922 159114 147978
rect 159170 147922 159238 147978
rect 159294 147922 159362 147978
rect 159418 147922 159486 147978
rect 159542 147922 159638 147978
rect 142828 144116 142884 144126
rect 142044 139636 142100 139646
rect 140812 124562 140868 124572
rect 140924 139412 140980 139422
rect 140924 123956 140980 139356
rect 141932 137818 141988 137828
rect 141036 127988 141092 127998
rect 141036 127738 141092 127932
rect 141036 127672 141092 127682
rect 140924 123890 140980 123900
rect 136892 118514 136948 118524
rect 141036 122724 141092 122734
rect 132018 118294 132114 118350
rect 132170 118294 132238 118350
rect 132294 118294 132362 118350
rect 132418 118294 132486 118350
rect 132542 118294 132638 118350
rect 132018 118226 132638 118294
rect 132018 118170 132114 118226
rect 132170 118170 132238 118226
rect 132294 118170 132362 118226
rect 132418 118170 132486 118226
rect 132542 118170 132638 118226
rect 132018 118102 132638 118170
rect 132018 118046 132114 118102
rect 132170 118046 132238 118102
rect 132294 118046 132362 118102
rect 132418 118046 132486 118102
rect 132542 118046 132638 118102
rect 132018 117978 132638 118046
rect 132018 117922 132114 117978
rect 132170 117922 132238 117978
rect 132294 117922 132362 117978
rect 132418 117922 132486 117978
rect 132542 117922 132638 117978
rect 132018 100350 132638 117922
rect 141036 116564 141092 122668
rect 141932 118468 141988 137762
rect 142044 122724 142100 139580
rect 142828 139412 142884 144060
rect 142828 139346 142884 139356
rect 143612 139860 143668 139870
rect 142044 122658 142100 122668
rect 141932 118402 141988 118412
rect 143612 117236 143668 139804
rect 148448 130350 148768 130384
rect 148448 130294 148518 130350
rect 148574 130294 148642 130350
rect 148698 130294 148768 130350
rect 148448 130226 148768 130294
rect 148448 130170 148518 130226
rect 148574 130170 148642 130226
rect 148698 130170 148768 130226
rect 148448 130102 148768 130170
rect 148448 130046 148518 130102
rect 148574 130046 148642 130102
rect 148698 130046 148768 130102
rect 148448 129978 148768 130046
rect 148448 129922 148518 129978
rect 148574 129922 148642 129978
rect 148698 129922 148768 129978
rect 148448 129888 148768 129922
rect 159018 130350 159638 147922
rect 159018 130294 159114 130350
rect 159170 130294 159238 130350
rect 159294 130294 159362 130350
rect 159418 130294 159486 130350
rect 159542 130294 159638 130350
rect 159018 130226 159638 130294
rect 159018 130170 159114 130226
rect 159170 130170 159238 130226
rect 159294 130170 159362 130226
rect 159418 130170 159486 130226
rect 159542 130170 159638 130226
rect 159018 130102 159638 130170
rect 159018 130046 159114 130102
rect 159170 130046 159238 130102
rect 159294 130046 159362 130102
rect 159418 130046 159486 130102
rect 159542 130046 159638 130102
rect 159018 129978 159638 130046
rect 159018 129922 159114 129978
rect 159170 129922 159238 129978
rect 159294 129922 159362 129978
rect 159418 129922 159486 129978
rect 159542 129922 159638 129978
rect 144060 128098 144116 128108
rect 144060 127988 144116 128042
rect 144060 127922 144116 127932
rect 143612 117170 143668 117180
rect 141036 116498 141092 116508
rect 148448 112350 148768 112384
rect 148448 112294 148518 112350
rect 148574 112294 148642 112350
rect 148698 112294 148768 112350
rect 148448 112226 148768 112294
rect 148448 112170 148518 112226
rect 148574 112170 148642 112226
rect 148698 112170 148768 112226
rect 148448 112102 148768 112170
rect 148448 112046 148518 112102
rect 148574 112046 148642 112102
rect 148698 112046 148768 112102
rect 148448 111978 148768 112046
rect 148448 111922 148518 111978
rect 148574 111922 148642 111978
rect 148698 111922 148768 111978
rect 148448 111888 148768 111922
rect 159018 112350 159638 129922
rect 162738 172350 163358 184626
rect 179168 184350 179488 184384
rect 179168 184294 179238 184350
rect 179294 184294 179362 184350
rect 179418 184294 179488 184350
rect 179168 184226 179488 184294
rect 179168 184170 179238 184226
rect 179294 184170 179362 184226
rect 179418 184170 179488 184226
rect 179168 184102 179488 184170
rect 179168 184046 179238 184102
rect 179294 184046 179362 184102
rect 179418 184046 179488 184102
rect 179168 183978 179488 184046
rect 179168 183922 179238 183978
rect 179294 183922 179362 183978
rect 179418 183922 179488 183978
rect 179168 183888 179488 183922
rect 189738 184350 190358 201922
rect 192332 222628 192388 222638
rect 191548 195058 191604 195068
rect 191548 186058 191604 195002
rect 192332 193844 192388 222572
rect 192332 193778 192388 193788
rect 193458 208350 194078 225922
rect 193458 208294 193554 208350
rect 193610 208294 193678 208350
rect 193734 208294 193802 208350
rect 193858 208294 193926 208350
rect 193982 208294 194078 208350
rect 193458 208226 194078 208294
rect 193458 208170 193554 208226
rect 193610 208170 193678 208226
rect 193734 208170 193802 208226
rect 193858 208170 193926 208226
rect 193982 208170 194078 208226
rect 193458 208102 194078 208170
rect 193458 208046 193554 208102
rect 193610 208046 193678 208102
rect 193734 208046 193802 208102
rect 193858 208046 193926 208102
rect 193982 208046 194078 208102
rect 193458 207978 194078 208046
rect 193458 207922 193554 207978
rect 193610 207922 193678 207978
rect 193734 207922 193802 207978
rect 193858 207922 193926 207978
rect 193982 207922 194078 207978
rect 191548 185992 191604 186002
rect 193458 190350 194078 207922
rect 197372 226436 197428 226446
rect 197372 197204 197428 226380
rect 197372 197138 197428 197148
rect 196588 196858 196644 196868
rect 196588 196532 196644 196802
rect 196588 196466 196644 196476
rect 197484 196678 197540 196688
rect 193458 190294 193554 190350
rect 193610 190294 193678 190350
rect 193734 190294 193802 190350
rect 193858 190294 193926 190350
rect 193982 190294 194078 190350
rect 193458 190226 194078 190294
rect 193458 190170 193554 190226
rect 193610 190170 193678 190226
rect 193734 190170 193802 190226
rect 193858 190170 193926 190226
rect 193982 190170 194078 190226
rect 193458 190102 194078 190170
rect 193458 190046 193554 190102
rect 193610 190046 193678 190102
rect 193734 190046 193802 190102
rect 193858 190046 193926 190102
rect 193982 190046 194078 190102
rect 193458 189978 194078 190046
rect 193458 189922 193554 189978
rect 193610 189922 193678 189978
rect 193734 189922 193802 189978
rect 193858 189922 193926 189978
rect 193982 189922 194078 189978
rect 189738 184294 189834 184350
rect 189890 184294 189958 184350
rect 190014 184294 190082 184350
rect 190138 184294 190206 184350
rect 190262 184294 190358 184350
rect 189738 184226 190358 184294
rect 189738 184170 189834 184226
rect 189890 184170 189958 184226
rect 190014 184170 190082 184226
rect 190138 184170 190206 184226
rect 190262 184170 190358 184226
rect 189738 184102 190358 184170
rect 189738 184046 189834 184102
rect 189890 184046 189958 184102
rect 190014 184046 190082 184102
rect 190138 184046 190206 184102
rect 190262 184046 190358 184102
rect 189738 183978 190358 184046
rect 189738 183922 189834 183978
rect 189890 183922 189958 183978
rect 190014 183922 190082 183978
rect 190138 183922 190206 183978
rect 190262 183922 190358 183978
rect 162738 172294 162834 172350
rect 162890 172294 162958 172350
rect 163014 172294 163082 172350
rect 163138 172294 163206 172350
rect 163262 172294 163358 172350
rect 162738 172226 163358 172294
rect 162738 172170 162834 172226
rect 162890 172170 162958 172226
rect 163014 172170 163082 172226
rect 163138 172170 163206 172226
rect 163262 172170 163358 172226
rect 162738 172102 163358 172170
rect 162738 172046 162834 172102
rect 162890 172046 162958 172102
rect 163014 172046 163082 172102
rect 163138 172046 163206 172102
rect 163262 172046 163358 172102
rect 162738 171978 163358 172046
rect 162738 171922 162834 171978
rect 162890 171922 162958 171978
rect 163014 171922 163082 171978
rect 163138 171922 163206 171978
rect 163262 171922 163358 171978
rect 162738 154350 163358 171922
rect 162738 154294 162834 154350
rect 162890 154294 162958 154350
rect 163014 154294 163082 154350
rect 163138 154294 163206 154350
rect 163262 154294 163358 154350
rect 162738 154226 163358 154294
rect 162738 154170 162834 154226
rect 162890 154170 162958 154226
rect 163014 154170 163082 154226
rect 163138 154170 163206 154226
rect 163262 154170 163358 154226
rect 162738 154102 163358 154170
rect 162738 154046 162834 154102
rect 162890 154046 162958 154102
rect 163014 154046 163082 154102
rect 163138 154046 163206 154102
rect 163262 154046 163358 154102
rect 162738 153978 163358 154046
rect 162738 153922 162834 153978
rect 162890 153922 162958 153978
rect 163014 153922 163082 153978
rect 163138 153922 163206 153978
rect 163262 153922 163358 153978
rect 162738 136350 163358 153922
rect 188972 169876 189028 169886
rect 162738 136294 162834 136350
rect 162890 136294 162958 136350
rect 163014 136294 163082 136350
rect 163138 136294 163206 136350
rect 163262 136294 163358 136350
rect 162738 136226 163358 136294
rect 162738 136170 162834 136226
rect 162890 136170 162958 136226
rect 163014 136170 163082 136226
rect 163138 136170 163206 136226
rect 163262 136170 163358 136226
rect 162738 136102 163358 136170
rect 162738 136046 162834 136102
rect 162890 136046 162958 136102
rect 163014 136046 163082 136102
rect 163138 136046 163206 136102
rect 163262 136046 163358 136102
rect 162738 135978 163358 136046
rect 162738 135922 162834 135978
rect 162890 135922 162958 135978
rect 163014 135922 163082 135978
rect 163138 135922 163206 135978
rect 163262 135922 163358 135978
rect 162738 125678 163358 135922
rect 163808 136350 164128 136384
rect 163808 136294 163878 136350
rect 163934 136294 164002 136350
rect 164058 136294 164128 136350
rect 163808 136226 164128 136294
rect 163808 136170 163878 136226
rect 163934 136170 164002 136226
rect 164058 136170 164128 136226
rect 163808 136102 164128 136170
rect 163808 136046 163878 136102
rect 163934 136046 164002 136102
rect 164058 136046 164128 136102
rect 163808 135978 164128 136046
rect 163808 135922 163878 135978
rect 163934 135922 164002 135978
rect 164058 135922 164128 135978
rect 163808 135888 164128 135922
rect 179168 130350 179488 130384
rect 179168 130294 179238 130350
rect 179294 130294 179362 130350
rect 179418 130294 179488 130350
rect 179168 130226 179488 130294
rect 179168 130170 179238 130226
rect 179294 130170 179362 130226
rect 179418 130170 179488 130226
rect 179168 130102 179488 130170
rect 179168 130046 179238 130102
rect 179294 130046 179362 130102
rect 179418 130046 179488 130102
rect 179168 129978 179488 130046
rect 179168 129922 179238 129978
rect 179294 129922 179362 129978
rect 179418 129922 179488 129978
rect 179168 129888 179488 129922
rect 188972 124628 189028 169820
rect 189738 166350 190358 183922
rect 189738 166294 189834 166350
rect 189890 166294 189958 166350
rect 190014 166294 190082 166350
rect 190138 166294 190206 166350
rect 190262 166294 190358 166350
rect 189738 166226 190358 166294
rect 189738 166170 189834 166226
rect 189890 166170 189958 166226
rect 190014 166170 190082 166226
rect 190138 166170 190206 166226
rect 190262 166170 190358 166226
rect 189738 166102 190358 166170
rect 189738 166046 189834 166102
rect 189890 166046 189958 166102
rect 190014 166046 190082 166102
rect 190138 166046 190206 166102
rect 190262 166046 190358 166102
rect 189738 165978 190358 166046
rect 189738 165922 189834 165978
rect 189890 165922 189958 165978
rect 190014 165922 190082 165978
rect 190138 165922 190206 165978
rect 190262 165922 190358 165978
rect 189738 148350 190358 165922
rect 193458 172350 194078 189922
rect 197484 187796 197540 196622
rect 197484 187730 197540 187740
rect 193458 172294 193554 172350
rect 193610 172294 193678 172350
rect 193734 172294 193802 172350
rect 193858 172294 193926 172350
rect 193982 172294 194078 172350
rect 193458 172226 194078 172294
rect 193458 172170 193554 172226
rect 193610 172170 193678 172226
rect 193734 172170 193802 172226
rect 193858 172170 193926 172226
rect 193982 172170 194078 172226
rect 193458 172102 194078 172170
rect 193458 172046 193554 172102
rect 193610 172046 193678 172102
rect 193734 172046 193802 172102
rect 193858 172046 193926 172102
rect 193982 172046 194078 172102
rect 193458 171978 194078 172046
rect 193458 171922 193554 171978
rect 193610 171922 193678 171978
rect 193734 171922 193802 171978
rect 193858 171922 193926 171978
rect 193982 171922 194078 171978
rect 189738 148294 189834 148350
rect 189890 148294 189958 148350
rect 190014 148294 190082 148350
rect 190138 148294 190206 148350
rect 190262 148294 190358 148350
rect 189738 148226 190358 148294
rect 189738 148170 189834 148226
rect 189890 148170 189958 148226
rect 190014 148170 190082 148226
rect 190138 148170 190206 148226
rect 190262 148170 190358 148226
rect 189738 148102 190358 148170
rect 189738 148046 189834 148102
rect 189890 148046 189958 148102
rect 190014 148046 190082 148102
rect 190138 148046 190206 148102
rect 190262 148046 190358 148102
rect 189738 147978 190358 148046
rect 189738 147922 189834 147978
rect 189890 147922 189958 147978
rect 190014 147922 190082 147978
rect 190138 147922 190206 147978
rect 190262 147922 190358 147978
rect 188972 124562 189028 124572
rect 189084 138628 189140 138638
rect 189084 121268 189140 138572
rect 189738 130350 190358 147922
rect 189738 130294 189834 130350
rect 189890 130294 189958 130350
rect 190014 130294 190082 130350
rect 190138 130294 190206 130350
rect 190262 130294 190358 130350
rect 189738 130226 190358 130294
rect 189738 130170 189834 130226
rect 189890 130170 189958 130226
rect 190014 130170 190082 130226
rect 190138 130170 190206 130226
rect 190262 130170 190358 130226
rect 189738 130102 190358 130170
rect 189738 130046 189834 130102
rect 189890 130046 189958 130102
rect 190014 130046 190082 130102
rect 190138 130046 190206 130102
rect 190262 130046 190358 130102
rect 189738 129978 190358 130046
rect 189738 129922 189834 129978
rect 189890 129922 189958 129978
rect 190014 129922 190082 129978
rect 190138 129922 190206 129978
rect 190262 129922 190358 129978
rect 189084 121202 189140 121212
rect 189532 121268 189588 121278
rect 159018 112294 159114 112350
rect 159170 112294 159238 112350
rect 159294 112294 159362 112350
rect 159418 112294 159486 112350
rect 159542 112294 159638 112350
rect 159018 112226 159638 112294
rect 159018 112170 159114 112226
rect 159170 112170 159238 112226
rect 159294 112170 159362 112226
rect 159418 112170 159486 112226
rect 159542 112170 159638 112226
rect 159018 112102 159638 112170
rect 159018 112046 159114 112102
rect 159170 112046 159238 112102
rect 159294 112046 159362 112102
rect 159418 112046 159486 112102
rect 159542 112046 159638 112102
rect 159018 111978 159638 112046
rect 159018 111922 159114 111978
rect 159170 111922 159238 111978
rect 159294 111922 159362 111978
rect 159418 111922 159486 111978
rect 159542 111922 159638 111978
rect 132018 100294 132114 100350
rect 132170 100294 132238 100350
rect 132294 100294 132362 100350
rect 132418 100294 132486 100350
rect 132542 100294 132638 100350
rect 132018 100226 132638 100294
rect 132018 100170 132114 100226
rect 132170 100170 132238 100226
rect 132294 100170 132362 100226
rect 132418 100170 132486 100226
rect 132542 100170 132638 100226
rect 132018 100102 132638 100170
rect 132018 100046 132114 100102
rect 132170 100046 132238 100102
rect 132294 100046 132362 100102
rect 132418 100046 132486 100102
rect 132542 100046 132638 100102
rect 132018 99978 132638 100046
rect 132018 99922 132114 99978
rect 132170 99922 132238 99978
rect 132294 99922 132362 99978
rect 132418 99922 132486 99978
rect 132542 99922 132638 99978
rect 132018 82350 132638 99922
rect 132018 82294 132114 82350
rect 132170 82294 132238 82350
rect 132294 82294 132362 82350
rect 132418 82294 132486 82350
rect 132542 82294 132638 82350
rect 132018 82226 132638 82294
rect 132018 82170 132114 82226
rect 132170 82170 132238 82226
rect 132294 82170 132362 82226
rect 132418 82170 132486 82226
rect 132542 82170 132638 82226
rect 132018 82102 132638 82170
rect 132018 82046 132114 82102
rect 132170 82046 132238 82102
rect 132294 82046 132362 82102
rect 132418 82046 132486 82102
rect 132542 82046 132638 82102
rect 132018 81978 132638 82046
rect 132018 81922 132114 81978
rect 132170 81922 132238 81978
rect 132294 81922 132362 81978
rect 132418 81922 132486 81978
rect 132542 81922 132638 81978
rect 128298 76294 128394 76350
rect 128450 76294 128518 76350
rect 128574 76294 128642 76350
rect 128698 76294 128766 76350
rect 128822 76294 128918 76350
rect 128298 76226 128918 76294
rect 128298 76170 128394 76226
rect 128450 76170 128518 76226
rect 128574 76170 128642 76226
rect 128698 76170 128766 76226
rect 128822 76170 128918 76226
rect 128298 76102 128918 76170
rect 128298 76046 128394 76102
rect 128450 76046 128518 76102
rect 128574 76046 128642 76102
rect 128698 76046 128766 76102
rect 128822 76046 128918 76102
rect 128298 75978 128918 76046
rect 128298 75922 128394 75978
rect 128450 75922 128518 75978
rect 128574 75922 128642 75978
rect 128698 75922 128766 75978
rect 128822 75922 128918 75978
rect 126924 69748 126980 69758
rect 126924 54180 126980 69692
rect 126924 54114 126980 54124
rect 128298 58350 128918 75922
rect 128298 58294 128394 58350
rect 128450 58294 128518 58350
rect 128574 58294 128642 58350
rect 128698 58294 128766 58350
rect 128822 58294 128918 58350
rect 128298 58226 128918 58294
rect 128298 58170 128394 58226
rect 128450 58170 128518 58226
rect 128574 58170 128642 58226
rect 128698 58170 128766 58226
rect 128822 58170 128918 58226
rect 128298 58102 128918 58170
rect 128298 58046 128394 58102
rect 128450 58046 128518 58102
rect 128574 58046 128642 58102
rect 128698 58046 128766 58102
rect 128822 58046 128918 58102
rect 128298 57978 128918 58046
rect 128298 57922 128394 57978
rect 128450 57922 128518 57978
rect 128574 57922 128642 57978
rect 128698 57922 128766 57978
rect 128822 57922 128918 57978
rect 126812 50754 126868 50764
rect 127596 50596 127652 50606
rect 82012 47394 82068 47404
rect 80444 46722 80500 46732
rect 80220 46050 80276 46060
rect 101808 46350 102128 46384
rect 101808 46294 101878 46350
rect 101934 46294 102002 46350
rect 102058 46294 102128 46350
rect 101808 46226 102128 46294
rect 101808 46170 101878 46226
rect 101934 46170 102002 46226
rect 102058 46170 102128 46226
rect 101808 46102 102128 46170
rect 70578 45978 71198 46046
rect 70578 45922 70674 45978
rect 70730 45922 70798 45978
rect 70854 45922 70922 45978
rect 70978 45922 71046 45978
rect 71102 45922 71198 45978
rect 66858 40294 66954 40350
rect 67010 40294 67078 40350
rect 67134 40294 67202 40350
rect 67258 40294 67326 40350
rect 67382 40294 67478 40350
rect 66858 40226 67478 40294
rect 66858 40170 66954 40226
rect 67010 40170 67078 40226
rect 67134 40170 67202 40226
rect 67258 40170 67326 40226
rect 67382 40170 67478 40226
rect 66858 40102 67478 40170
rect 66858 40046 66954 40102
rect 67010 40046 67078 40102
rect 67134 40046 67202 40102
rect 67258 40046 67326 40102
rect 67382 40046 67478 40102
rect 66858 39978 67478 40046
rect 66858 39922 66954 39978
rect 67010 39922 67078 39978
rect 67134 39922 67202 39978
rect 67258 39922 67326 39978
rect 67382 39922 67478 39978
rect 36138 22294 36234 22350
rect 36290 22294 36358 22350
rect 36414 22294 36482 22350
rect 36538 22294 36606 22350
rect 36662 22294 36758 22350
rect 36138 22226 36758 22294
rect 36138 22170 36234 22226
rect 36290 22170 36358 22226
rect 36414 22170 36482 22226
rect 36538 22170 36606 22226
rect 36662 22170 36758 22226
rect 36138 22102 36758 22170
rect 36138 22046 36234 22102
rect 36290 22046 36358 22102
rect 36414 22046 36482 22102
rect 36538 22046 36606 22102
rect 36662 22046 36758 22102
rect 36138 21978 36758 22046
rect 36138 21922 36234 21978
rect 36290 21922 36358 21978
rect 36414 21922 36482 21978
rect 36538 21922 36606 21978
rect 36662 21922 36758 21978
rect 9138 -1176 9234 -1120
rect 9290 -1176 9358 -1120
rect 9414 -1176 9482 -1120
rect 9538 -1176 9606 -1120
rect 9662 -1176 9758 -1120
rect 9138 -1244 9758 -1176
rect 9138 -1300 9234 -1244
rect 9290 -1300 9358 -1244
rect 9414 -1300 9482 -1244
rect 9538 -1300 9606 -1244
rect 9662 -1300 9758 -1244
rect 9138 -1368 9758 -1300
rect 9138 -1424 9234 -1368
rect 9290 -1424 9358 -1368
rect 9414 -1424 9482 -1368
rect 9538 -1424 9606 -1368
rect 9662 -1424 9758 -1368
rect 9138 -1492 9758 -1424
rect 9138 -1548 9234 -1492
rect 9290 -1548 9358 -1492
rect 9414 -1548 9482 -1492
rect 9538 -1548 9606 -1492
rect 9662 -1548 9758 -1492
rect 9138 -1644 9758 -1548
rect 36138 4350 36758 21922
rect 36138 4294 36234 4350
rect 36290 4294 36358 4350
rect 36414 4294 36482 4350
rect 36538 4294 36606 4350
rect 36662 4294 36758 4350
rect 36138 4226 36758 4294
rect 36138 4170 36234 4226
rect 36290 4170 36358 4226
rect 36414 4170 36482 4226
rect 36538 4170 36606 4226
rect 36662 4170 36758 4226
rect 36138 4102 36758 4170
rect 36138 4046 36234 4102
rect 36290 4046 36358 4102
rect 36414 4046 36482 4102
rect 36538 4046 36606 4102
rect 36662 4046 36758 4102
rect 36138 3978 36758 4046
rect 36138 3922 36234 3978
rect 36290 3922 36358 3978
rect 36414 3922 36482 3978
rect 36538 3922 36606 3978
rect 36662 3922 36758 3978
rect 36138 -160 36758 3922
rect 36138 -216 36234 -160
rect 36290 -216 36358 -160
rect 36414 -216 36482 -160
rect 36538 -216 36606 -160
rect 36662 -216 36758 -160
rect 36138 -284 36758 -216
rect 36138 -340 36234 -284
rect 36290 -340 36358 -284
rect 36414 -340 36482 -284
rect 36538 -340 36606 -284
rect 36662 -340 36758 -284
rect 36138 -408 36758 -340
rect 36138 -464 36234 -408
rect 36290 -464 36358 -408
rect 36414 -464 36482 -408
rect 36538 -464 36606 -408
rect 36662 -464 36758 -408
rect 36138 -532 36758 -464
rect 36138 -588 36234 -532
rect 36290 -588 36358 -532
rect 36414 -588 36482 -532
rect 36538 -588 36606 -532
rect 36662 -588 36758 -532
rect 36138 -1644 36758 -588
rect 39858 28350 40478 30164
rect 39858 28294 39954 28350
rect 40010 28294 40078 28350
rect 40134 28294 40202 28350
rect 40258 28294 40326 28350
rect 40382 28294 40478 28350
rect 39858 28226 40478 28294
rect 39858 28170 39954 28226
rect 40010 28170 40078 28226
rect 40134 28170 40202 28226
rect 40258 28170 40326 28226
rect 40382 28170 40478 28226
rect 39858 28102 40478 28170
rect 39858 28046 39954 28102
rect 40010 28046 40078 28102
rect 40134 28046 40202 28102
rect 40258 28046 40326 28102
rect 40382 28046 40478 28102
rect 39858 27978 40478 28046
rect 39858 27922 39954 27978
rect 40010 27922 40078 27978
rect 40134 27922 40202 27978
rect 40258 27922 40326 27978
rect 40382 27922 40478 27978
rect 39858 10350 40478 27922
rect 39858 10294 39954 10350
rect 40010 10294 40078 10350
rect 40134 10294 40202 10350
rect 40258 10294 40326 10350
rect 40382 10294 40478 10350
rect 39858 10226 40478 10294
rect 39858 10170 39954 10226
rect 40010 10170 40078 10226
rect 40134 10170 40202 10226
rect 40258 10170 40326 10226
rect 40382 10170 40478 10226
rect 39858 10102 40478 10170
rect 39858 10046 39954 10102
rect 40010 10046 40078 10102
rect 40134 10046 40202 10102
rect 40258 10046 40326 10102
rect 40382 10046 40478 10102
rect 39858 9978 40478 10046
rect 39858 9922 39954 9978
rect 40010 9922 40078 9978
rect 40134 9922 40202 9978
rect 40258 9922 40326 9978
rect 40382 9922 40478 9978
rect 39858 -1120 40478 9922
rect 39858 -1176 39954 -1120
rect 40010 -1176 40078 -1120
rect 40134 -1176 40202 -1120
rect 40258 -1176 40326 -1120
rect 40382 -1176 40478 -1120
rect 39858 -1244 40478 -1176
rect 39858 -1300 39954 -1244
rect 40010 -1300 40078 -1244
rect 40134 -1300 40202 -1244
rect 40258 -1300 40326 -1244
rect 40382 -1300 40478 -1244
rect 39858 -1368 40478 -1300
rect 39858 -1424 39954 -1368
rect 40010 -1424 40078 -1368
rect 40134 -1424 40202 -1368
rect 40258 -1424 40326 -1368
rect 40382 -1424 40478 -1368
rect 39858 -1492 40478 -1424
rect 39858 -1548 39954 -1492
rect 40010 -1548 40078 -1492
rect 40134 -1548 40202 -1492
rect 40258 -1548 40326 -1492
rect 40382 -1548 40478 -1492
rect 39858 -1644 40478 -1548
rect 66858 22350 67478 39922
rect 66858 22294 66954 22350
rect 67010 22294 67078 22350
rect 67134 22294 67202 22350
rect 67258 22294 67326 22350
rect 67382 22294 67478 22350
rect 66858 22226 67478 22294
rect 66858 22170 66954 22226
rect 67010 22170 67078 22226
rect 67134 22170 67202 22226
rect 67258 22170 67326 22226
rect 67382 22170 67478 22226
rect 66858 22102 67478 22170
rect 66858 22046 66954 22102
rect 67010 22046 67078 22102
rect 67134 22046 67202 22102
rect 67258 22046 67326 22102
rect 67382 22046 67478 22102
rect 66858 21978 67478 22046
rect 66858 21922 66954 21978
rect 67010 21922 67078 21978
rect 67134 21922 67202 21978
rect 67258 21922 67326 21978
rect 67382 21922 67478 21978
rect 66858 4350 67478 21922
rect 66858 4294 66954 4350
rect 67010 4294 67078 4350
rect 67134 4294 67202 4350
rect 67258 4294 67326 4350
rect 67382 4294 67478 4350
rect 66858 4226 67478 4294
rect 66858 4170 66954 4226
rect 67010 4170 67078 4226
rect 67134 4170 67202 4226
rect 67258 4170 67326 4226
rect 67382 4170 67478 4226
rect 66858 4102 67478 4170
rect 66858 4046 66954 4102
rect 67010 4046 67078 4102
rect 67134 4046 67202 4102
rect 67258 4046 67326 4102
rect 67382 4046 67478 4102
rect 66858 3978 67478 4046
rect 66858 3922 66954 3978
rect 67010 3922 67078 3978
rect 67134 3922 67202 3978
rect 67258 3922 67326 3978
rect 67382 3922 67478 3978
rect 66858 -160 67478 3922
rect 66858 -216 66954 -160
rect 67010 -216 67078 -160
rect 67134 -216 67202 -160
rect 67258 -216 67326 -160
rect 67382 -216 67478 -160
rect 66858 -284 67478 -216
rect 66858 -340 66954 -284
rect 67010 -340 67078 -284
rect 67134 -340 67202 -284
rect 67258 -340 67326 -284
rect 67382 -340 67478 -284
rect 66858 -408 67478 -340
rect 66858 -464 66954 -408
rect 67010 -464 67078 -408
rect 67134 -464 67202 -408
rect 67258 -464 67326 -408
rect 67382 -464 67478 -408
rect 66858 -532 67478 -464
rect 66858 -588 66954 -532
rect 67010 -588 67078 -532
rect 67134 -588 67202 -532
rect 67258 -588 67326 -532
rect 67382 -588 67478 -532
rect 66858 -1644 67478 -588
rect 70578 28350 71198 45922
rect 101808 46046 101878 46102
rect 101934 46046 102002 46102
rect 102058 46046 102128 46102
rect 127596 46116 127652 50540
rect 127596 46050 127652 46060
rect 101808 45978 102128 46046
rect 101808 45922 101878 45978
rect 101934 45922 102002 45978
rect 102058 45922 102128 45978
rect 101808 45888 102128 45922
rect 86448 40350 86768 40384
rect 86448 40294 86518 40350
rect 86574 40294 86642 40350
rect 86698 40294 86768 40350
rect 86448 40226 86768 40294
rect 86448 40170 86518 40226
rect 86574 40170 86642 40226
rect 86698 40170 86768 40226
rect 86448 40102 86768 40170
rect 86448 40046 86518 40102
rect 86574 40046 86642 40102
rect 86698 40046 86768 40102
rect 86448 39978 86768 40046
rect 86448 39922 86518 39978
rect 86574 39922 86642 39978
rect 86698 39922 86768 39978
rect 86448 39888 86768 39922
rect 97578 40350 98198 44578
rect 97578 40294 97674 40350
rect 97730 40294 97798 40350
rect 97854 40294 97922 40350
rect 97978 40294 98046 40350
rect 98102 40294 98198 40350
rect 97578 40226 98198 40294
rect 97578 40170 97674 40226
rect 97730 40170 97798 40226
rect 97854 40170 97922 40226
rect 97978 40170 98046 40226
rect 98102 40170 98198 40226
rect 97578 40102 98198 40170
rect 97578 40046 97674 40102
rect 97730 40046 97798 40102
rect 97854 40046 97922 40102
rect 97978 40046 98046 40102
rect 98102 40046 98198 40102
rect 97578 39978 98198 40046
rect 97578 39922 97674 39978
rect 97730 39922 97798 39978
rect 97854 39922 97922 39978
rect 97978 39922 98046 39978
rect 98102 39922 98198 39978
rect 70578 28294 70674 28350
rect 70730 28294 70798 28350
rect 70854 28294 70922 28350
rect 70978 28294 71046 28350
rect 71102 28294 71198 28350
rect 70578 28226 71198 28294
rect 70578 28170 70674 28226
rect 70730 28170 70798 28226
rect 70854 28170 70922 28226
rect 70978 28170 71046 28226
rect 71102 28170 71198 28226
rect 70578 28102 71198 28170
rect 70578 28046 70674 28102
rect 70730 28046 70798 28102
rect 70854 28046 70922 28102
rect 70978 28046 71046 28102
rect 71102 28046 71198 28102
rect 70578 27978 71198 28046
rect 70578 27922 70674 27978
rect 70730 27922 70798 27978
rect 70854 27922 70922 27978
rect 70978 27922 71046 27978
rect 71102 27922 71198 27978
rect 70578 10350 71198 27922
rect 70578 10294 70674 10350
rect 70730 10294 70798 10350
rect 70854 10294 70922 10350
rect 70978 10294 71046 10350
rect 71102 10294 71198 10350
rect 70578 10226 71198 10294
rect 70578 10170 70674 10226
rect 70730 10170 70798 10226
rect 70854 10170 70922 10226
rect 70978 10170 71046 10226
rect 71102 10170 71198 10226
rect 70578 10102 71198 10170
rect 70578 10046 70674 10102
rect 70730 10046 70798 10102
rect 70854 10046 70922 10102
rect 70978 10046 71046 10102
rect 71102 10046 71198 10102
rect 70578 9978 71198 10046
rect 70578 9922 70674 9978
rect 70730 9922 70798 9978
rect 70854 9922 70922 9978
rect 70978 9922 71046 9978
rect 71102 9922 71198 9978
rect 70578 -1120 71198 9922
rect 70578 -1176 70674 -1120
rect 70730 -1176 70798 -1120
rect 70854 -1176 70922 -1120
rect 70978 -1176 71046 -1120
rect 71102 -1176 71198 -1120
rect 70578 -1244 71198 -1176
rect 70578 -1300 70674 -1244
rect 70730 -1300 70798 -1244
rect 70854 -1300 70922 -1244
rect 70978 -1300 71046 -1244
rect 71102 -1300 71198 -1244
rect 70578 -1368 71198 -1300
rect 70578 -1424 70674 -1368
rect 70730 -1424 70798 -1368
rect 70854 -1424 70922 -1368
rect 70978 -1424 71046 -1368
rect 71102 -1424 71198 -1368
rect 70578 -1492 71198 -1424
rect 70578 -1548 70674 -1492
rect 70730 -1548 70798 -1492
rect 70854 -1548 70922 -1492
rect 70978 -1548 71046 -1492
rect 71102 -1548 71198 -1492
rect 70578 -1644 71198 -1548
rect 97578 22350 98198 39922
rect 117168 40350 117488 40384
rect 117168 40294 117238 40350
rect 117294 40294 117362 40350
rect 117418 40294 117488 40350
rect 117168 40226 117488 40294
rect 117168 40170 117238 40226
rect 117294 40170 117362 40226
rect 117418 40170 117488 40226
rect 117168 40102 117488 40170
rect 117168 40046 117238 40102
rect 117294 40046 117362 40102
rect 117418 40046 117488 40102
rect 117168 39978 117488 40046
rect 117168 39922 117238 39978
rect 117294 39922 117362 39978
rect 117418 39922 117488 39978
rect 117168 39888 117488 39922
rect 128298 40350 128918 57922
rect 130172 78036 130228 78046
rect 130172 50596 130228 77980
rect 130172 50530 130228 50540
rect 132018 64350 132638 81922
rect 132018 64294 132114 64350
rect 132170 64294 132238 64350
rect 132294 64294 132362 64350
rect 132418 64294 132486 64350
rect 132542 64294 132638 64350
rect 132018 64226 132638 64294
rect 132018 64170 132114 64226
rect 132170 64170 132238 64226
rect 132294 64170 132362 64226
rect 132418 64170 132486 64226
rect 132542 64170 132638 64226
rect 132018 64102 132638 64170
rect 132018 64046 132114 64102
rect 132170 64046 132238 64102
rect 132294 64046 132362 64102
rect 132418 64046 132486 64102
rect 132542 64046 132638 64102
rect 132018 63978 132638 64046
rect 132018 63922 132114 63978
rect 132170 63922 132238 63978
rect 132294 63922 132362 63978
rect 132418 63922 132486 63978
rect 132542 63922 132638 63978
rect 128298 40294 128394 40350
rect 128450 40294 128518 40350
rect 128574 40294 128642 40350
rect 128698 40294 128766 40350
rect 128822 40294 128918 40350
rect 128298 40226 128918 40294
rect 128298 40170 128394 40226
rect 128450 40170 128518 40226
rect 128574 40170 128642 40226
rect 128698 40170 128766 40226
rect 128822 40170 128918 40226
rect 128298 40102 128918 40170
rect 128298 40046 128394 40102
rect 128450 40046 128518 40102
rect 128574 40046 128642 40102
rect 128698 40046 128766 40102
rect 128822 40046 128918 40102
rect 128298 39978 128918 40046
rect 128298 39922 128394 39978
rect 128450 39922 128518 39978
rect 128574 39922 128642 39978
rect 128698 39922 128766 39978
rect 128822 39922 128918 39978
rect 97578 22294 97674 22350
rect 97730 22294 97798 22350
rect 97854 22294 97922 22350
rect 97978 22294 98046 22350
rect 98102 22294 98198 22350
rect 97578 22226 98198 22294
rect 97578 22170 97674 22226
rect 97730 22170 97798 22226
rect 97854 22170 97922 22226
rect 97978 22170 98046 22226
rect 98102 22170 98198 22226
rect 97578 22102 98198 22170
rect 97578 22046 97674 22102
rect 97730 22046 97798 22102
rect 97854 22046 97922 22102
rect 97978 22046 98046 22102
rect 98102 22046 98198 22102
rect 97578 21978 98198 22046
rect 97578 21922 97674 21978
rect 97730 21922 97798 21978
rect 97854 21922 97922 21978
rect 97978 21922 98046 21978
rect 98102 21922 98198 21978
rect 97578 4350 98198 21922
rect 97578 4294 97674 4350
rect 97730 4294 97798 4350
rect 97854 4294 97922 4350
rect 97978 4294 98046 4350
rect 98102 4294 98198 4350
rect 97578 4226 98198 4294
rect 97578 4170 97674 4226
rect 97730 4170 97798 4226
rect 97854 4170 97922 4226
rect 97978 4170 98046 4226
rect 98102 4170 98198 4226
rect 97578 4102 98198 4170
rect 97578 4046 97674 4102
rect 97730 4046 97798 4102
rect 97854 4046 97922 4102
rect 97978 4046 98046 4102
rect 98102 4046 98198 4102
rect 97578 3978 98198 4046
rect 97578 3922 97674 3978
rect 97730 3922 97798 3978
rect 97854 3922 97922 3978
rect 97978 3922 98046 3978
rect 98102 3922 98198 3978
rect 97578 -160 98198 3922
rect 97578 -216 97674 -160
rect 97730 -216 97798 -160
rect 97854 -216 97922 -160
rect 97978 -216 98046 -160
rect 98102 -216 98198 -160
rect 97578 -284 98198 -216
rect 97578 -340 97674 -284
rect 97730 -340 97798 -284
rect 97854 -340 97922 -284
rect 97978 -340 98046 -284
rect 98102 -340 98198 -284
rect 97578 -408 98198 -340
rect 97578 -464 97674 -408
rect 97730 -464 97798 -408
rect 97854 -464 97922 -408
rect 97978 -464 98046 -408
rect 98102 -464 98198 -408
rect 97578 -532 98198 -464
rect 97578 -588 97674 -532
rect 97730 -588 97798 -532
rect 97854 -588 97922 -532
rect 97978 -588 98046 -532
rect 98102 -588 98198 -532
rect 97578 -1644 98198 -588
rect 101298 28350 101918 30164
rect 101298 28294 101394 28350
rect 101450 28294 101518 28350
rect 101574 28294 101642 28350
rect 101698 28294 101766 28350
rect 101822 28294 101918 28350
rect 101298 28226 101918 28294
rect 101298 28170 101394 28226
rect 101450 28170 101518 28226
rect 101574 28170 101642 28226
rect 101698 28170 101766 28226
rect 101822 28170 101918 28226
rect 101298 28102 101918 28170
rect 101298 28046 101394 28102
rect 101450 28046 101518 28102
rect 101574 28046 101642 28102
rect 101698 28046 101766 28102
rect 101822 28046 101918 28102
rect 101298 27978 101918 28046
rect 101298 27922 101394 27978
rect 101450 27922 101518 27978
rect 101574 27922 101642 27978
rect 101698 27922 101766 27978
rect 101822 27922 101918 27978
rect 101298 10350 101918 27922
rect 101298 10294 101394 10350
rect 101450 10294 101518 10350
rect 101574 10294 101642 10350
rect 101698 10294 101766 10350
rect 101822 10294 101918 10350
rect 101298 10226 101918 10294
rect 101298 10170 101394 10226
rect 101450 10170 101518 10226
rect 101574 10170 101642 10226
rect 101698 10170 101766 10226
rect 101822 10170 101918 10226
rect 101298 10102 101918 10170
rect 101298 10046 101394 10102
rect 101450 10046 101518 10102
rect 101574 10046 101642 10102
rect 101698 10046 101766 10102
rect 101822 10046 101918 10102
rect 101298 9978 101918 10046
rect 101298 9922 101394 9978
rect 101450 9922 101518 9978
rect 101574 9922 101642 9978
rect 101698 9922 101766 9978
rect 101822 9922 101918 9978
rect 101298 -1120 101918 9922
rect 101298 -1176 101394 -1120
rect 101450 -1176 101518 -1120
rect 101574 -1176 101642 -1120
rect 101698 -1176 101766 -1120
rect 101822 -1176 101918 -1120
rect 101298 -1244 101918 -1176
rect 101298 -1300 101394 -1244
rect 101450 -1300 101518 -1244
rect 101574 -1300 101642 -1244
rect 101698 -1300 101766 -1244
rect 101822 -1300 101918 -1244
rect 101298 -1368 101918 -1300
rect 101298 -1424 101394 -1368
rect 101450 -1424 101518 -1368
rect 101574 -1424 101642 -1368
rect 101698 -1424 101766 -1368
rect 101822 -1424 101918 -1368
rect 101298 -1492 101918 -1424
rect 101298 -1548 101394 -1492
rect 101450 -1548 101518 -1492
rect 101574 -1548 101642 -1492
rect 101698 -1548 101766 -1492
rect 101822 -1548 101918 -1492
rect 101298 -1644 101918 -1548
rect 128298 22350 128918 39922
rect 128298 22294 128394 22350
rect 128450 22294 128518 22350
rect 128574 22294 128642 22350
rect 128698 22294 128766 22350
rect 128822 22294 128918 22350
rect 128298 22226 128918 22294
rect 128298 22170 128394 22226
rect 128450 22170 128518 22226
rect 128574 22170 128642 22226
rect 128698 22170 128766 22226
rect 128822 22170 128918 22226
rect 128298 22102 128918 22170
rect 128298 22046 128394 22102
rect 128450 22046 128518 22102
rect 128574 22046 128642 22102
rect 128698 22046 128766 22102
rect 128822 22046 128918 22102
rect 128298 21978 128918 22046
rect 128298 21922 128394 21978
rect 128450 21922 128518 21978
rect 128574 21922 128642 21978
rect 128698 21922 128766 21978
rect 128822 21922 128918 21978
rect 128298 4350 128918 21922
rect 128298 4294 128394 4350
rect 128450 4294 128518 4350
rect 128574 4294 128642 4350
rect 128698 4294 128766 4350
rect 128822 4294 128918 4350
rect 128298 4226 128918 4294
rect 128298 4170 128394 4226
rect 128450 4170 128518 4226
rect 128574 4170 128642 4226
rect 128698 4170 128766 4226
rect 128822 4170 128918 4226
rect 128298 4102 128918 4170
rect 128298 4046 128394 4102
rect 128450 4046 128518 4102
rect 128574 4046 128642 4102
rect 128698 4046 128766 4102
rect 128822 4046 128918 4102
rect 128298 3978 128918 4046
rect 128298 3922 128394 3978
rect 128450 3922 128518 3978
rect 128574 3922 128642 3978
rect 128698 3922 128766 3978
rect 128822 3922 128918 3978
rect 128298 -160 128918 3922
rect 128298 -216 128394 -160
rect 128450 -216 128518 -160
rect 128574 -216 128642 -160
rect 128698 -216 128766 -160
rect 128822 -216 128918 -160
rect 128298 -284 128918 -216
rect 128298 -340 128394 -284
rect 128450 -340 128518 -284
rect 128574 -340 128642 -284
rect 128698 -340 128766 -284
rect 128822 -340 128918 -284
rect 128298 -408 128918 -340
rect 128298 -464 128394 -408
rect 128450 -464 128518 -408
rect 128574 -464 128642 -408
rect 128698 -464 128766 -408
rect 128822 -464 128918 -408
rect 128298 -532 128918 -464
rect 128298 -588 128394 -532
rect 128450 -588 128518 -532
rect 128574 -588 128642 -532
rect 128698 -588 128766 -532
rect 128822 -588 128918 -532
rect 128298 -1644 128918 -588
rect 132018 46350 132638 63922
rect 133532 103348 133588 103358
rect 133532 49476 133588 103292
rect 136892 101668 136948 101678
rect 133532 49410 133588 49420
rect 135212 74116 135268 74126
rect 135212 47124 135268 74060
rect 136892 50148 136948 101612
rect 143612 101556 143668 101566
rect 138572 99988 138628 99998
rect 138572 66276 138628 99932
rect 142716 96740 142772 96750
rect 141932 88340 141988 88350
rect 140588 85316 140644 85326
rect 138572 66210 138628 66220
rect 138684 73108 138740 73118
rect 138684 55524 138740 73052
rect 138684 55458 138740 55468
rect 136892 50082 136948 50092
rect 135212 47058 135268 47068
rect 132018 46294 132114 46350
rect 132170 46294 132238 46350
rect 132294 46294 132362 46350
rect 132418 46294 132486 46350
rect 132542 46294 132638 46350
rect 132018 46226 132638 46294
rect 132018 46170 132114 46226
rect 132170 46170 132238 46226
rect 132294 46170 132362 46226
rect 132418 46170 132486 46226
rect 132542 46170 132638 46226
rect 132018 46102 132638 46170
rect 132018 46046 132114 46102
rect 132170 46046 132238 46102
rect 132294 46046 132362 46102
rect 132418 46046 132486 46102
rect 132542 46046 132638 46102
rect 140588 46116 140644 85260
rect 140924 83636 140980 83646
rect 140812 70420 140868 70430
rect 140700 68852 140756 68862
rect 140700 53508 140756 68796
rect 140812 54180 140868 70364
rect 140812 54114 140868 54124
rect 140700 53442 140756 53452
rect 140588 46050 140644 46060
rect 132018 45978 132638 46046
rect 132018 45922 132114 45978
rect 132170 45922 132238 45978
rect 132294 45922 132362 45978
rect 132418 45922 132486 45978
rect 132542 45922 132638 45978
rect 132018 28350 132638 45922
rect 140924 45444 140980 83580
rect 141036 56278 141092 56288
rect 141036 56196 141092 56222
rect 141036 56130 141092 56140
rect 141932 54852 141988 88284
rect 141932 54786 141988 54796
rect 142044 81396 142100 81406
rect 142044 49252 142100 81340
rect 142604 80276 142660 80286
rect 142604 52836 142660 80220
rect 142716 65604 142772 96684
rect 142716 65538 142772 65548
rect 143612 56308 143668 101500
rect 159018 94350 159638 111922
rect 162738 118350 163358 120034
rect 162738 118294 162834 118350
rect 162890 118294 162958 118350
rect 163014 118294 163082 118350
rect 163138 118294 163206 118350
rect 163262 118294 163358 118350
rect 162738 118226 163358 118294
rect 162738 118170 162834 118226
rect 162890 118170 162958 118226
rect 163014 118170 163082 118226
rect 163138 118170 163206 118226
rect 163262 118170 163358 118226
rect 162738 118102 163358 118170
rect 162738 118046 162834 118102
rect 162890 118046 162958 118102
rect 163014 118046 163082 118102
rect 163138 118046 163206 118102
rect 163262 118046 163358 118102
rect 162738 117978 163358 118046
rect 162738 117922 162834 117978
rect 162890 117922 162958 117978
rect 163014 117922 163082 117978
rect 163138 117922 163206 117978
rect 163262 117922 163358 117978
rect 160860 101780 160916 101790
rect 160860 100996 160916 101724
rect 160860 100930 160916 100940
rect 159018 94294 159114 94350
rect 159170 94294 159238 94350
rect 159294 94294 159362 94350
rect 159418 94294 159486 94350
rect 159542 94294 159638 94350
rect 159018 94226 159638 94294
rect 159018 94170 159114 94226
rect 159170 94170 159238 94226
rect 159294 94170 159362 94226
rect 159418 94170 159486 94226
rect 159542 94170 159638 94226
rect 159018 94102 159638 94170
rect 159018 94046 159114 94102
rect 159170 94046 159238 94102
rect 159294 94046 159362 94102
rect 159418 94046 159486 94102
rect 159542 94046 159638 94102
rect 159018 93978 159638 94046
rect 159018 93922 159114 93978
rect 159170 93922 159238 93978
rect 159294 93922 159362 93978
rect 159418 93922 159486 93978
rect 159542 93922 159638 93978
rect 146972 83076 147028 83086
rect 145292 82516 145348 82526
rect 144060 79716 144116 79726
rect 144060 67228 144116 79660
rect 143612 56242 143668 56252
rect 143948 67172 144116 67228
rect 144284 78260 144340 78270
rect 143948 55468 144004 67172
rect 144060 56278 144116 56288
rect 144060 56196 144116 56222
rect 144060 56130 144116 56140
rect 143948 55412 144116 55468
rect 142604 52770 142660 52780
rect 144060 49476 144116 55412
rect 144284 50148 144340 78204
rect 145292 68852 145348 82460
rect 146972 70420 147028 83020
rect 146972 70354 147028 70364
rect 159018 76350 159638 93922
rect 159018 76294 159114 76350
rect 159170 76294 159238 76350
rect 159294 76294 159362 76350
rect 159418 76294 159486 76350
rect 159542 76294 159638 76350
rect 159018 76226 159638 76294
rect 159018 76170 159114 76226
rect 159170 76170 159238 76226
rect 159294 76170 159362 76226
rect 159418 76170 159486 76226
rect 159542 76170 159638 76226
rect 159018 76102 159638 76170
rect 159018 76046 159114 76102
rect 159170 76046 159238 76102
rect 159294 76046 159362 76102
rect 159418 76046 159486 76102
rect 159542 76046 159638 76102
rect 159018 75978 159638 76046
rect 159018 75922 159114 75978
rect 159170 75922 159238 75978
rect 159294 75922 159362 75978
rect 159418 75922 159486 75978
rect 159542 75922 159638 75978
rect 145292 68786 145348 68796
rect 148448 58350 148768 58384
rect 148448 58294 148518 58350
rect 148574 58294 148642 58350
rect 148698 58294 148768 58350
rect 148448 58226 148768 58294
rect 148448 58170 148518 58226
rect 148574 58170 148642 58226
rect 148698 58170 148768 58226
rect 148448 58102 148768 58170
rect 148448 58046 148518 58102
rect 148574 58046 148642 58102
rect 148698 58046 148768 58102
rect 148448 57978 148768 58046
rect 148448 57922 148518 57978
rect 148574 57922 148642 57978
rect 148698 57922 148768 57978
rect 148448 57888 148768 57922
rect 159018 58350 159638 75922
rect 159018 58294 159114 58350
rect 159170 58294 159238 58350
rect 159294 58294 159362 58350
rect 159418 58294 159486 58350
rect 159542 58294 159638 58350
rect 159018 58226 159638 58294
rect 159018 58170 159114 58226
rect 159170 58170 159238 58226
rect 159294 58170 159362 58226
rect 159418 58170 159486 58226
rect 159542 58170 159638 58226
rect 159018 58102 159638 58170
rect 159018 58046 159114 58102
rect 159170 58046 159238 58102
rect 159294 58046 159362 58102
rect 159418 58046 159486 58102
rect 159542 58046 159638 58102
rect 159018 57978 159638 58046
rect 159018 57922 159114 57978
rect 159170 57922 159238 57978
rect 159294 57922 159362 57978
rect 159418 57922 159486 57978
rect 159542 57922 159638 57978
rect 144284 50082 144340 50092
rect 144060 49410 144116 49420
rect 142044 49186 142100 49196
rect 140924 45378 140980 45388
rect 148448 40350 148768 40384
rect 148448 40294 148518 40350
rect 148574 40294 148642 40350
rect 148698 40294 148768 40350
rect 148448 40226 148768 40294
rect 148448 40170 148518 40226
rect 148574 40170 148642 40226
rect 148698 40170 148768 40226
rect 148448 40102 148768 40170
rect 148448 40046 148518 40102
rect 148574 40046 148642 40102
rect 148698 40046 148768 40102
rect 148448 39978 148768 40046
rect 148448 39922 148518 39978
rect 148574 39922 148642 39978
rect 148698 39922 148768 39978
rect 148448 39888 148768 39922
rect 159018 40350 159638 57922
rect 162738 100350 163358 117922
rect 163808 118350 164128 118384
rect 163808 118294 163878 118350
rect 163934 118294 164002 118350
rect 164058 118294 164128 118350
rect 163808 118226 164128 118294
rect 163808 118170 163878 118226
rect 163934 118170 164002 118226
rect 164058 118170 164128 118226
rect 163808 118102 164128 118170
rect 163808 118046 163878 118102
rect 163934 118046 164002 118102
rect 164058 118046 164128 118102
rect 163808 117978 164128 118046
rect 163808 117922 163878 117978
rect 163934 117922 164002 117978
rect 164058 117922 164128 117978
rect 163808 117888 164128 117922
rect 189532 117908 189588 121212
rect 189532 117842 189588 117852
rect 179168 112350 179488 112384
rect 179168 112294 179238 112350
rect 179294 112294 179362 112350
rect 179418 112294 179488 112350
rect 179168 112226 179488 112294
rect 179168 112170 179238 112226
rect 179294 112170 179362 112226
rect 179418 112170 179488 112226
rect 179168 112102 179488 112170
rect 179168 112046 179238 112102
rect 179294 112046 179362 112102
rect 179418 112046 179488 112102
rect 179168 111978 179488 112046
rect 179168 111922 179238 111978
rect 179294 111922 179362 111978
rect 179418 111922 179488 111978
rect 179168 111888 179488 111922
rect 189738 112350 190358 129922
rect 192332 162148 192388 162158
rect 192332 125300 192388 162092
rect 192332 125234 192388 125244
rect 193458 154350 194078 171922
rect 197372 167636 197428 167646
rect 193458 154294 193554 154350
rect 193610 154294 193678 154350
rect 193734 154294 193802 154350
rect 193858 154294 193926 154350
rect 193982 154294 194078 154350
rect 193458 154226 194078 154294
rect 193458 154170 193554 154226
rect 193610 154170 193678 154226
rect 193734 154170 193802 154226
rect 193858 154170 193926 154226
rect 193982 154170 194078 154226
rect 193458 154102 194078 154170
rect 193458 154046 193554 154102
rect 193610 154046 193678 154102
rect 193734 154046 193802 154102
rect 193858 154046 193926 154102
rect 193982 154046 194078 154102
rect 193458 153978 194078 154046
rect 193458 153922 193554 153978
rect 193610 153922 193678 153978
rect 193734 153922 193802 153978
rect 193858 153922 193926 153978
rect 193982 153922 194078 153978
rect 193458 136350 194078 153922
rect 193458 136294 193554 136350
rect 193610 136294 193678 136350
rect 193734 136294 193802 136350
rect 193858 136294 193926 136350
rect 193982 136294 194078 136350
rect 193458 136226 194078 136294
rect 193458 136170 193554 136226
rect 193610 136170 193678 136226
rect 193734 136170 193802 136226
rect 193858 136170 193926 136226
rect 193982 136170 194078 136226
rect 193458 136102 194078 136170
rect 193458 136046 193554 136102
rect 193610 136046 193678 136102
rect 193734 136046 193802 136102
rect 193858 136046 193926 136102
rect 193982 136046 194078 136102
rect 193458 135978 194078 136046
rect 193458 135922 193554 135978
rect 193610 135922 193678 135978
rect 193734 135922 193802 135978
rect 193858 135922 193926 135978
rect 193982 135922 194078 135978
rect 189738 112294 189834 112350
rect 189890 112294 189958 112350
rect 190014 112294 190082 112350
rect 190138 112294 190206 112350
rect 190262 112294 190358 112350
rect 189738 112226 190358 112294
rect 189738 112170 189834 112226
rect 189890 112170 189958 112226
rect 190014 112170 190082 112226
rect 190138 112170 190206 112226
rect 190262 112170 190358 112226
rect 189738 112102 190358 112170
rect 189738 112046 189834 112102
rect 189890 112046 189958 112102
rect 190014 112046 190082 112102
rect 190138 112046 190206 112102
rect 190262 112046 190358 112102
rect 189738 111978 190358 112046
rect 189738 111922 189834 111978
rect 189890 111922 189958 111978
rect 190014 111922 190082 111978
rect 190138 111922 190206 111978
rect 190262 111922 190358 111978
rect 162738 100294 162834 100350
rect 162890 100294 162958 100350
rect 163014 100294 163082 100350
rect 163138 100294 163206 100350
rect 163262 100294 163358 100350
rect 162738 100226 163358 100294
rect 162738 100170 162834 100226
rect 162890 100170 162958 100226
rect 163014 100170 163082 100226
rect 163138 100170 163206 100226
rect 163262 100170 163358 100226
rect 162738 100102 163358 100170
rect 162738 100046 162834 100102
rect 162890 100046 162958 100102
rect 163014 100046 163082 100102
rect 163138 100046 163206 100102
rect 163262 100046 163358 100102
rect 162738 99978 163358 100046
rect 162738 99922 162834 99978
rect 162890 99922 162958 99978
rect 163014 99922 163082 99978
rect 163138 99922 163206 99978
rect 163262 99922 163358 99978
rect 162738 82350 163358 99922
rect 189738 94350 190358 111922
rect 189738 94294 189834 94350
rect 189890 94294 189958 94350
rect 190014 94294 190082 94350
rect 190138 94294 190206 94350
rect 190262 94294 190358 94350
rect 189738 94226 190358 94294
rect 189738 94170 189834 94226
rect 189890 94170 189958 94226
rect 190014 94170 190082 94226
rect 190138 94170 190206 94226
rect 190262 94170 190358 94226
rect 189738 94102 190358 94170
rect 189738 94046 189834 94102
rect 189890 94046 189958 94102
rect 190014 94046 190082 94102
rect 190138 94046 190206 94102
rect 190262 94046 190358 94102
rect 189738 93978 190358 94046
rect 189738 93922 189834 93978
rect 189890 93922 189958 93978
rect 190014 93922 190082 93978
rect 190138 93922 190206 93978
rect 190262 93922 190358 93978
rect 162738 82294 162834 82350
rect 162890 82294 162958 82350
rect 163014 82294 163082 82350
rect 163138 82294 163206 82350
rect 163262 82294 163358 82350
rect 162738 82226 163358 82294
rect 162738 82170 162834 82226
rect 162890 82170 162958 82226
rect 163014 82170 163082 82226
rect 163138 82170 163206 82226
rect 163262 82170 163358 82226
rect 162738 82102 163358 82170
rect 162738 82046 162834 82102
rect 162890 82046 162958 82102
rect 163014 82046 163082 82102
rect 163138 82046 163206 82102
rect 163262 82046 163358 82102
rect 162738 81978 163358 82046
rect 162738 81922 162834 81978
rect 162890 81922 162958 81978
rect 163014 81922 163082 81978
rect 163138 81922 163206 81978
rect 163262 81922 163358 81978
rect 162738 64350 163358 81922
rect 188972 91924 189028 91934
rect 188076 76916 188132 76926
rect 188076 71428 188132 76860
rect 188076 71362 188132 71372
rect 162738 64294 162834 64350
rect 162890 64294 162958 64350
rect 163014 64294 163082 64350
rect 163138 64294 163206 64350
rect 163262 64294 163358 64350
rect 162738 64226 163358 64294
rect 162738 64170 162834 64226
rect 162890 64170 162958 64226
rect 163014 64170 163082 64226
rect 163138 64170 163206 64226
rect 163262 64170 163358 64226
rect 162738 64102 163358 64170
rect 162738 64046 162834 64102
rect 162890 64046 162958 64102
rect 163014 64046 163082 64102
rect 163138 64046 163206 64102
rect 163262 64046 163358 64102
rect 162738 63978 163358 64046
rect 162738 63922 162834 63978
rect 162890 63922 162958 63978
rect 163014 63922 163082 63978
rect 163138 63922 163206 63978
rect 163262 63922 163358 63978
rect 162738 53358 163358 63922
rect 163808 64350 164128 64384
rect 163808 64294 163878 64350
rect 163934 64294 164002 64350
rect 164058 64294 164128 64350
rect 163808 64226 164128 64294
rect 163808 64170 163878 64226
rect 163934 64170 164002 64226
rect 164058 64170 164128 64226
rect 163808 64102 164128 64170
rect 163808 64046 163878 64102
rect 163934 64046 164002 64102
rect 164058 64046 164128 64102
rect 163808 63978 164128 64046
rect 163808 63922 163878 63978
rect 163934 63922 164002 63978
rect 164058 63922 164128 63978
rect 163808 63888 164128 63922
rect 179168 58350 179488 58384
rect 179168 58294 179238 58350
rect 179294 58294 179362 58350
rect 179418 58294 179488 58350
rect 179168 58226 179488 58294
rect 179168 58170 179238 58226
rect 179294 58170 179362 58226
rect 179418 58170 179488 58226
rect 179168 58102 179488 58170
rect 179168 58046 179238 58102
rect 179294 58046 179362 58102
rect 179418 58046 179488 58102
rect 179168 57978 179488 58046
rect 179168 57922 179238 57978
rect 179294 57922 179362 57978
rect 179418 57922 179488 57978
rect 179168 57888 179488 57922
rect 188972 54180 189028 91868
rect 189738 76350 190358 93922
rect 189738 76294 189834 76350
rect 189890 76294 189958 76350
rect 190014 76294 190082 76350
rect 190138 76294 190206 76350
rect 190262 76294 190358 76350
rect 189738 76226 190358 76294
rect 189738 76170 189834 76226
rect 189890 76170 189958 76226
rect 190014 76170 190082 76226
rect 190138 76170 190206 76226
rect 190262 76170 190358 76226
rect 189738 76102 190358 76170
rect 189738 76046 189834 76102
rect 189890 76046 189958 76102
rect 190014 76046 190082 76102
rect 190138 76046 190206 76102
rect 190262 76046 190358 76102
rect 189738 75978 190358 76046
rect 189738 75922 189834 75978
rect 189890 75922 189958 75978
rect 190014 75922 190082 75978
rect 190138 75922 190206 75978
rect 190262 75922 190358 75978
rect 188972 54114 189028 54124
rect 189084 73220 189140 73230
rect 189084 49476 189140 73164
rect 189420 71540 189476 71550
rect 189196 71428 189252 71438
rect 189196 52164 189252 71372
rect 189308 69860 189364 69870
rect 189308 54852 189364 69804
rect 189420 65604 189476 71484
rect 189420 65538 189476 65548
rect 189308 54786 189364 54796
rect 189738 58350 190358 75922
rect 189738 58294 189834 58350
rect 189890 58294 189958 58350
rect 190014 58294 190082 58350
rect 190138 58294 190206 58350
rect 190262 58294 190358 58350
rect 189738 58226 190358 58294
rect 189738 58170 189834 58226
rect 189890 58170 189958 58226
rect 190014 58170 190082 58226
rect 190138 58170 190206 58226
rect 190262 58170 190358 58226
rect 189738 58102 190358 58170
rect 189738 58046 189834 58102
rect 189890 58046 189958 58102
rect 190014 58046 190082 58102
rect 190138 58046 190206 58102
rect 190262 58046 190358 58102
rect 189738 57978 190358 58046
rect 189738 57922 189834 57978
rect 189890 57922 189958 57978
rect 190014 57922 190082 57978
rect 190138 57922 190206 57978
rect 190262 57922 190358 57978
rect 189196 52098 189252 52108
rect 189084 49410 189140 49420
rect 189532 48692 189588 48702
rect 159018 40294 159114 40350
rect 159170 40294 159238 40350
rect 159294 40294 159362 40350
rect 159418 40294 159486 40350
rect 159542 40294 159638 40350
rect 159018 40226 159638 40294
rect 159018 40170 159114 40226
rect 159170 40170 159238 40226
rect 159294 40170 159362 40226
rect 159418 40170 159486 40226
rect 159542 40170 159638 40226
rect 159018 40102 159638 40170
rect 159018 40046 159114 40102
rect 159170 40046 159238 40102
rect 159294 40046 159362 40102
rect 159418 40046 159486 40102
rect 159542 40046 159638 40102
rect 159018 39978 159638 40046
rect 159018 39922 159114 39978
rect 159170 39922 159238 39978
rect 159294 39922 159362 39978
rect 159418 39922 159486 39978
rect 159542 39922 159638 39978
rect 132018 28294 132114 28350
rect 132170 28294 132238 28350
rect 132294 28294 132362 28350
rect 132418 28294 132486 28350
rect 132542 28294 132638 28350
rect 132018 28226 132638 28294
rect 132018 28170 132114 28226
rect 132170 28170 132238 28226
rect 132294 28170 132362 28226
rect 132418 28170 132486 28226
rect 132542 28170 132638 28226
rect 132018 28102 132638 28170
rect 132018 28046 132114 28102
rect 132170 28046 132238 28102
rect 132294 28046 132362 28102
rect 132418 28046 132486 28102
rect 132542 28046 132638 28102
rect 132018 27978 132638 28046
rect 132018 27922 132114 27978
rect 132170 27922 132238 27978
rect 132294 27922 132362 27978
rect 132418 27922 132486 27978
rect 132542 27922 132638 27978
rect 132018 10350 132638 27922
rect 132018 10294 132114 10350
rect 132170 10294 132238 10350
rect 132294 10294 132362 10350
rect 132418 10294 132486 10350
rect 132542 10294 132638 10350
rect 132018 10226 132638 10294
rect 132018 10170 132114 10226
rect 132170 10170 132238 10226
rect 132294 10170 132362 10226
rect 132418 10170 132486 10226
rect 132542 10170 132638 10226
rect 132018 10102 132638 10170
rect 132018 10046 132114 10102
rect 132170 10046 132238 10102
rect 132294 10046 132362 10102
rect 132418 10046 132486 10102
rect 132542 10046 132638 10102
rect 132018 9978 132638 10046
rect 132018 9922 132114 9978
rect 132170 9922 132238 9978
rect 132294 9922 132362 9978
rect 132418 9922 132486 9978
rect 132542 9922 132638 9978
rect 132018 -1120 132638 9922
rect 132018 -1176 132114 -1120
rect 132170 -1176 132238 -1120
rect 132294 -1176 132362 -1120
rect 132418 -1176 132486 -1120
rect 132542 -1176 132638 -1120
rect 132018 -1244 132638 -1176
rect 132018 -1300 132114 -1244
rect 132170 -1300 132238 -1244
rect 132294 -1300 132362 -1244
rect 132418 -1300 132486 -1244
rect 132542 -1300 132638 -1244
rect 132018 -1368 132638 -1300
rect 132018 -1424 132114 -1368
rect 132170 -1424 132238 -1368
rect 132294 -1424 132362 -1368
rect 132418 -1424 132486 -1368
rect 132542 -1424 132638 -1368
rect 132018 -1492 132638 -1424
rect 132018 -1548 132114 -1492
rect 132170 -1548 132238 -1492
rect 132294 -1548 132362 -1492
rect 132418 -1548 132486 -1492
rect 132542 -1548 132638 -1492
rect 132018 -1644 132638 -1548
rect 159018 22350 159638 39922
rect 159018 22294 159114 22350
rect 159170 22294 159238 22350
rect 159294 22294 159362 22350
rect 159418 22294 159486 22350
rect 159542 22294 159638 22350
rect 159018 22226 159638 22294
rect 159018 22170 159114 22226
rect 159170 22170 159238 22226
rect 159294 22170 159362 22226
rect 159418 22170 159486 22226
rect 159542 22170 159638 22226
rect 159018 22102 159638 22170
rect 159018 22046 159114 22102
rect 159170 22046 159238 22102
rect 159294 22046 159362 22102
rect 159418 22046 159486 22102
rect 159542 22046 159638 22102
rect 159018 21978 159638 22046
rect 159018 21922 159114 21978
rect 159170 21922 159238 21978
rect 159294 21922 159362 21978
rect 159418 21922 159486 21978
rect 159542 21922 159638 21978
rect 159018 4350 159638 21922
rect 159018 4294 159114 4350
rect 159170 4294 159238 4350
rect 159294 4294 159362 4350
rect 159418 4294 159486 4350
rect 159542 4294 159638 4350
rect 159018 4226 159638 4294
rect 159018 4170 159114 4226
rect 159170 4170 159238 4226
rect 159294 4170 159362 4226
rect 159418 4170 159486 4226
rect 159542 4170 159638 4226
rect 159018 4102 159638 4170
rect 159018 4046 159114 4102
rect 159170 4046 159238 4102
rect 159294 4046 159362 4102
rect 159418 4046 159486 4102
rect 159542 4046 159638 4102
rect 159018 3978 159638 4046
rect 159018 3922 159114 3978
rect 159170 3922 159238 3978
rect 159294 3922 159362 3978
rect 159418 3922 159486 3978
rect 159542 3922 159638 3978
rect 159018 -160 159638 3922
rect 159018 -216 159114 -160
rect 159170 -216 159238 -160
rect 159294 -216 159362 -160
rect 159418 -216 159486 -160
rect 159542 -216 159638 -160
rect 159018 -284 159638 -216
rect 159018 -340 159114 -284
rect 159170 -340 159238 -284
rect 159294 -340 159362 -284
rect 159418 -340 159486 -284
rect 159542 -340 159638 -284
rect 159018 -408 159638 -340
rect 159018 -464 159114 -408
rect 159170 -464 159238 -408
rect 159294 -464 159362 -408
rect 159418 -464 159486 -408
rect 159542 -464 159638 -408
rect 159018 -532 159638 -464
rect 159018 -588 159114 -532
rect 159170 -588 159238 -532
rect 159294 -588 159362 -532
rect 159418 -588 159486 -532
rect 159542 -588 159638 -532
rect 159018 -1644 159638 -588
rect 162738 46350 163358 48274
rect 162738 46294 162834 46350
rect 162890 46294 162958 46350
rect 163014 46294 163082 46350
rect 163138 46294 163206 46350
rect 163262 46294 163358 46350
rect 162738 46226 163358 46294
rect 162738 46170 162834 46226
rect 162890 46170 162958 46226
rect 163014 46170 163082 46226
rect 163138 46170 163206 46226
rect 163262 46170 163358 46226
rect 162738 46102 163358 46170
rect 162738 46046 162834 46102
rect 162890 46046 162958 46102
rect 163014 46046 163082 46102
rect 163138 46046 163206 46102
rect 163262 46046 163358 46102
rect 162738 45978 163358 46046
rect 162738 45922 162834 45978
rect 162890 45922 162958 45978
rect 163014 45922 163082 45978
rect 163138 45922 163206 45978
rect 163262 45922 163358 45978
rect 162738 28350 163358 45922
rect 163808 46350 164128 46384
rect 163808 46294 163878 46350
rect 163934 46294 164002 46350
rect 164058 46294 164128 46350
rect 163808 46226 164128 46294
rect 163808 46170 163878 46226
rect 163934 46170 164002 46226
rect 164058 46170 164128 46226
rect 163808 46102 164128 46170
rect 163808 46046 163878 46102
rect 163934 46046 164002 46102
rect 164058 46046 164128 46102
rect 189532 46116 189588 48636
rect 189532 46050 189588 46060
rect 163808 45978 164128 46046
rect 163808 45922 163878 45978
rect 163934 45922 164002 45978
rect 164058 45922 164128 45978
rect 163808 45888 164128 45922
rect 179168 40350 179488 40384
rect 179168 40294 179238 40350
rect 179294 40294 179362 40350
rect 179418 40294 179488 40350
rect 179168 40226 179488 40294
rect 179168 40170 179238 40226
rect 179294 40170 179362 40226
rect 179418 40170 179488 40226
rect 179168 40102 179488 40170
rect 179168 40046 179238 40102
rect 179294 40046 179362 40102
rect 179418 40046 179488 40102
rect 179168 39978 179488 40046
rect 179168 39922 179238 39978
rect 179294 39922 179362 39978
rect 179418 39922 179488 39978
rect 179168 39888 179488 39922
rect 189738 40350 190358 57922
rect 189738 40294 189834 40350
rect 189890 40294 189958 40350
rect 190014 40294 190082 40350
rect 190138 40294 190206 40350
rect 190262 40294 190358 40350
rect 189738 40226 190358 40294
rect 189738 40170 189834 40226
rect 189890 40170 189958 40226
rect 190014 40170 190082 40226
rect 190138 40170 190206 40226
rect 190262 40170 190358 40226
rect 189738 40102 190358 40170
rect 189738 40046 189834 40102
rect 189890 40046 189958 40102
rect 190014 40046 190082 40102
rect 190138 40046 190206 40102
rect 190262 40046 190358 40102
rect 189738 39978 190358 40046
rect 189738 39922 189834 39978
rect 189890 39922 189958 39978
rect 190014 39922 190082 39978
rect 190138 39922 190206 39978
rect 190262 39922 190358 39978
rect 162738 28294 162834 28350
rect 162890 28294 162958 28350
rect 163014 28294 163082 28350
rect 163138 28294 163206 28350
rect 163262 28294 163358 28350
rect 162738 28226 163358 28294
rect 162738 28170 162834 28226
rect 162890 28170 162958 28226
rect 163014 28170 163082 28226
rect 163138 28170 163206 28226
rect 163262 28170 163358 28226
rect 162738 28102 163358 28170
rect 162738 28046 162834 28102
rect 162890 28046 162958 28102
rect 163014 28046 163082 28102
rect 163138 28046 163206 28102
rect 163262 28046 163358 28102
rect 162738 27978 163358 28046
rect 162738 27922 162834 27978
rect 162890 27922 162958 27978
rect 163014 27922 163082 27978
rect 163138 27922 163206 27978
rect 163262 27922 163358 27978
rect 162738 10350 163358 27922
rect 162738 10294 162834 10350
rect 162890 10294 162958 10350
rect 163014 10294 163082 10350
rect 163138 10294 163206 10350
rect 163262 10294 163358 10350
rect 162738 10226 163358 10294
rect 162738 10170 162834 10226
rect 162890 10170 162958 10226
rect 163014 10170 163082 10226
rect 163138 10170 163206 10226
rect 163262 10170 163358 10226
rect 162738 10102 163358 10170
rect 162738 10046 162834 10102
rect 162890 10046 162958 10102
rect 163014 10046 163082 10102
rect 163138 10046 163206 10102
rect 163262 10046 163358 10102
rect 162738 9978 163358 10046
rect 162738 9922 162834 9978
rect 162890 9922 162958 9978
rect 163014 9922 163082 9978
rect 163138 9922 163206 9978
rect 163262 9922 163358 9978
rect 162738 -1120 163358 9922
rect 162738 -1176 162834 -1120
rect 162890 -1176 162958 -1120
rect 163014 -1176 163082 -1120
rect 163138 -1176 163206 -1120
rect 163262 -1176 163358 -1120
rect 162738 -1244 163358 -1176
rect 162738 -1300 162834 -1244
rect 162890 -1300 162958 -1244
rect 163014 -1300 163082 -1244
rect 163138 -1300 163206 -1244
rect 163262 -1300 163358 -1244
rect 162738 -1368 163358 -1300
rect 162738 -1424 162834 -1368
rect 162890 -1424 162958 -1368
rect 163014 -1424 163082 -1368
rect 163138 -1424 163206 -1368
rect 163262 -1424 163358 -1368
rect 162738 -1492 163358 -1424
rect 162738 -1548 162834 -1492
rect 162890 -1548 162958 -1492
rect 163014 -1548 163082 -1492
rect 163138 -1548 163206 -1492
rect 163262 -1548 163358 -1492
rect 162738 -1644 163358 -1548
rect 189738 22350 190358 39922
rect 189738 22294 189834 22350
rect 189890 22294 189958 22350
rect 190014 22294 190082 22350
rect 190138 22294 190206 22350
rect 190262 22294 190358 22350
rect 189738 22226 190358 22294
rect 189738 22170 189834 22226
rect 189890 22170 189958 22226
rect 190014 22170 190082 22226
rect 190138 22170 190206 22226
rect 190262 22170 190358 22226
rect 189738 22102 190358 22170
rect 189738 22046 189834 22102
rect 189890 22046 189958 22102
rect 190014 22046 190082 22102
rect 190138 22046 190206 22102
rect 190262 22046 190358 22102
rect 189738 21978 190358 22046
rect 189738 21922 189834 21978
rect 189890 21922 189958 21978
rect 190014 21922 190082 21978
rect 190138 21922 190206 21978
rect 190262 21922 190358 21978
rect 189738 4350 190358 21922
rect 189738 4294 189834 4350
rect 189890 4294 189958 4350
rect 190014 4294 190082 4350
rect 190138 4294 190206 4350
rect 190262 4294 190358 4350
rect 189738 4226 190358 4294
rect 189738 4170 189834 4226
rect 189890 4170 189958 4226
rect 190014 4170 190082 4226
rect 190138 4170 190206 4226
rect 190262 4170 190358 4226
rect 189738 4102 190358 4170
rect 189738 4046 189834 4102
rect 189890 4046 189958 4102
rect 190014 4046 190082 4102
rect 190138 4046 190206 4102
rect 190262 4046 190358 4102
rect 189738 3978 190358 4046
rect 189738 3922 189834 3978
rect 189890 3922 189958 3978
rect 190014 3922 190082 3978
rect 190138 3922 190206 3978
rect 190262 3922 190358 3978
rect 189738 -160 190358 3922
rect 189738 -216 189834 -160
rect 189890 -216 189958 -160
rect 190014 -216 190082 -160
rect 190138 -216 190206 -160
rect 190262 -216 190358 -160
rect 189738 -284 190358 -216
rect 189738 -340 189834 -284
rect 189890 -340 189958 -284
rect 190014 -340 190082 -284
rect 190138 -340 190206 -284
rect 190262 -340 190358 -284
rect 189738 -408 190358 -340
rect 189738 -464 189834 -408
rect 189890 -464 189958 -408
rect 190014 -464 190082 -408
rect 190138 -464 190206 -408
rect 190262 -464 190358 -408
rect 189738 -532 190358 -464
rect 189738 -588 189834 -532
rect 189890 -588 189958 -532
rect 190014 -588 190082 -532
rect 190138 -588 190206 -532
rect 190262 -588 190358 -532
rect 189738 -1644 190358 -588
rect 193458 118350 194078 135922
rect 195692 163828 195748 163838
rect 195692 125972 195748 163772
rect 195692 125906 195748 125916
rect 195804 139076 195860 139086
rect 193458 118294 193554 118350
rect 193610 118294 193678 118350
rect 193734 118294 193802 118350
rect 193858 118294 193926 118350
rect 193982 118294 194078 118350
rect 193458 118226 194078 118294
rect 193458 118170 193554 118226
rect 193610 118170 193678 118226
rect 193734 118170 193802 118226
rect 193858 118170 193926 118226
rect 193982 118170 194078 118226
rect 193458 118102 194078 118170
rect 193458 118046 193554 118102
rect 193610 118046 193678 118102
rect 193734 118046 193802 118102
rect 193858 118046 193926 118102
rect 193982 118046 194078 118102
rect 193458 117978 194078 118046
rect 193458 117922 193554 117978
rect 193610 117922 193678 117978
rect 193734 117922 193802 117978
rect 193858 117922 193926 117978
rect 193982 117922 194078 117978
rect 193458 100350 194078 117922
rect 195804 117236 195860 139020
rect 197372 119364 197428 167580
rect 199052 167076 199108 167086
rect 197484 142212 197540 142222
rect 197484 121268 197540 142156
rect 199052 126644 199108 167020
rect 199052 126578 199108 126588
rect 199164 143556 199220 143566
rect 199164 122724 199220 143500
rect 199164 122658 199220 122668
rect 199276 139188 199332 139198
rect 197484 121202 197540 121212
rect 199276 120596 199332 139132
rect 199276 120530 199332 120540
rect 197372 119298 197428 119308
rect 195804 117170 195860 117180
rect 193458 100294 193554 100350
rect 193610 100294 193678 100350
rect 193734 100294 193802 100350
rect 193858 100294 193926 100350
rect 193982 100294 194078 100350
rect 193458 100226 194078 100294
rect 193458 100170 193554 100226
rect 193610 100170 193678 100226
rect 193734 100170 193802 100226
rect 193858 100170 193926 100226
rect 193982 100170 194078 100226
rect 193458 100102 194078 100170
rect 193458 100046 193554 100102
rect 193610 100046 193678 100102
rect 193734 100046 193802 100102
rect 193858 100046 193926 100102
rect 193982 100046 194078 100102
rect 193458 99978 194078 100046
rect 193458 99922 193554 99978
rect 193610 99922 193678 99978
rect 193734 99922 193802 99978
rect 193858 99922 193926 99978
rect 193982 99922 194078 99978
rect 193458 82350 194078 99922
rect 193458 82294 193554 82350
rect 193610 82294 193678 82350
rect 193734 82294 193802 82350
rect 193858 82294 193926 82350
rect 193982 82294 194078 82350
rect 193458 82226 194078 82294
rect 193458 82170 193554 82226
rect 193610 82170 193678 82226
rect 193734 82170 193802 82226
rect 193858 82170 193926 82226
rect 193982 82170 194078 82226
rect 193458 82102 194078 82170
rect 193458 82046 193554 82102
rect 193610 82046 193678 82102
rect 193734 82046 193802 82102
rect 193858 82046 193926 82102
rect 193982 82046 194078 82102
rect 193458 81978 194078 82046
rect 193458 81922 193554 81978
rect 193610 81922 193678 81978
rect 193734 81922 193802 81978
rect 193858 81922 193926 81978
rect 193982 81922 194078 81978
rect 193458 64350 194078 81922
rect 193458 64294 193554 64350
rect 193610 64294 193678 64350
rect 193734 64294 193802 64350
rect 193858 64294 193926 64350
rect 193982 64294 194078 64350
rect 193458 64226 194078 64294
rect 193458 64170 193554 64226
rect 193610 64170 193678 64226
rect 193734 64170 193802 64226
rect 193858 64170 193926 64226
rect 193982 64170 194078 64226
rect 193458 64102 194078 64170
rect 193458 64046 193554 64102
rect 193610 64046 193678 64102
rect 193734 64046 193802 64102
rect 193858 64046 193926 64102
rect 193982 64046 194078 64102
rect 193458 63978 194078 64046
rect 193458 63922 193554 63978
rect 193610 63922 193678 63978
rect 193734 63922 193802 63978
rect 193858 63922 193926 63978
rect 193982 63922 194078 63978
rect 193458 46350 194078 63922
rect 195692 103124 195748 103134
rect 195692 55524 195748 103068
rect 195692 55458 195748 55468
rect 197372 85876 197428 85886
rect 197372 47460 197428 85820
rect 199052 84196 199108 84206
rect 199052 48692 199108 84140
rect 199052 48626 199108 48636
rect 197372 47394 197428 47404
rect 193458 46294 193554 46350
rect 193610 46294 193678 46350
rect 193734 46294 193802 46350
rect 193858 46294 193926 46350
rect 193982 46294 194078 46350
rect 193458 46226 194078 46294
rect 193458 46170 193554 46226
rect 193610 46170 193678 46226
rect 193734 46170 193802 46226
rect 193858 46170 193926 46226
rect 193982 46170 194078 46226
rect 193458 46102 194078 46170
rect 193458 46046 193554 46102
rect 193610 46046 193678 46102
rect 193734 46046 193802 46102
rect 193858 46046 193926 46102
rect 193982 46046 194078 46102
rect 193458 45978 194078 46046
rect 193458 45922 193554 45978
rect 193610 45922 193678 45978
rect 193734 45922 193802 45978
rect 193858 45922 193926 45978
rect 193982 45922 194078 45978
rect 193458 28350 194078 45922
rect 193458 28294 193554 28350
rect 193610 28294 193678 28350
rect 193734 28294 193802 28350
rect 193858 28294 193926 28350
rect 193982 28294 194078 28350
rect 193458 28226 194078 28294
rect 193458 28170 193554 28226
rect 193610 28170 193678 28226
rect 193734 28170 193802 28226
rect 193858 28170 193926 28226
rect 193982 28170 194078 28226
rect 193458 28102 194078 28170
rect 193458 28046 193554 28102
rect 193610 28046 193678 28102
rect 193734 28046 193802 28102
rect 193858 28046 193926 28102
rect 193982 28046 194078 28102
rect 193458 27978 194078 28046
rect 193458 27922 193554 27978
rect 193610 27922 193678 27978
rect 193734 27922 193802 27978
rect 193858 27922 193926 27978
rect 193982 27922 194078 27978
rect 193458 10350 194078 27922
rect 193458 10294 193554 10350
rect 193610 10294 193678 10350
rect 193734 10294 193802 10350
rect 193858 10294 193926 10350
rect 193982 10294 194078 10350
rect 193458 10226 194078 10294
rect 193458 10170 193554 10226
rect 193610 10170 193678 10226
rect 193734 10170 193802 10226
rect 193858 10170 193926 10226
rect 193982 10170 194078 10226
rect 193458 10102 194078 10170
rect 193458 10046 193554 10102
rect 193610 10046 193678 10102
rect 193734 10046 193802 10102
rect 193858 10046 193926 10102
rect 193982 10046 194078 10102
rect 193458 9978 194078 10046
rect 193458 9922 193554 9978
rect 193610 9922 193678 9978
rect 193734 9922 193802 9978
rect 193858 9922 193926 9978
rect 193982 9922 194078 9978
rect 193458 -1120 194078 9922
rect 200844 8596 200900 571202
rect 210448 562350 210768 562384
rect 210448 562294 210518 562350
rect 210574 562294 210642 562350
rect 210698 562294 210768 562350
rect 210448 562226 210768 562294
rect 210448 562170 210518 562226
rect 210574 562170 210642 562226
rect 210698 562170 210768 562226
rect 210448 562102 210768 562170
rect 210448 562046 210518 562102
rect 210574 562046 210642 562102
rect 210698 562046 210768 562102
rect 210448 561978 210768 562046
rect 210448 561922 210518 561978
rect 210574 561922 210642 561978
rect 210698 561922 210768 561978
rect 210448 561888 210768 561922
rect 220458 562350 221078 579922
rect 220458 562294 220554 562350
rect 220610 562294 220678 562350
rect 220734 562294 220802 562350
rect 220858 562294 220926 562350
rect 220982 562294 221078 562350
rect 220458 562226 221078 562294
rect 220458 562170 220554 562226
rect 220610 562170 220678 562226
rect 220734 562170 220802 562226
rect 220858 562170 220926 562226
rect 220982 562170 221078 562226
rect 220458 562102 221078 562170
rect 220458 562046 220554 562102
rect 220610 562046 220678 562102
rect 220734 562046 220802 562102
rect 220858 562046 220926 562102
rect 220982 562046 221078 562102
rect 220458 561978 221078 562046
rect 220458 561922 220554 561978
rect 220610 561922 220678 561978
rect 220734 561922 220802 561978
rect 220858 561922 220926 561978
rect 220982 561922 221078 561978
rect 201628 555238 201684 555248
rect 201628 554596 201684 555182
rect 201628 554530 201684 554540
rect 204876 552580 204932 552590
rect 203196 551908 203252 551918
rect 203084 544516 203140 544526
rect 203084 544078 203140 544460
rect 203196 544404 203252 551852
rect 203196 544338 203252 544348
rect 204092 544404 204148 544414
rect 203084 544022 203252 544078
rect 203084 543844 203140 543854
rect 203084 523572 203140 543788
rect 203084 523506 203140 523516
rect 203196 501508 203252 544022
rect 203196 501442 203252 501452
rect 204092 496916 204148 544348
rect 204876 533458 204932 552524
rect 204876 533392 204932 533402
rect 205772 550004 205828 550014
rect 205772 529956 205828 549948
rect 210448 544350 210768 544384
rect 210448 544294 210518 544350
rect 210574 544294 210642 544350
rect 210698 544294 210768 544350
rect 210448 544226 210768 544294
rect 210448 544170 210518 544226
rect 210574 544170 210642 544226
rect 210698 544170 210768 544226
rect 210448 544102 210768 544170
rect 210448 544046 210518 544102
rect 210574 544046 210642 544102
rect 210698 544046 210768 544102
rect 210448 543978 210768 544046
rect 210448 543922 210518 543978
rect 210574 543922 210642 543978
rect 210698 543922 210768 543978
rect 210448 543888 210768 543922
rect 220458 544350 221078 561922
rect 224178 598172 224798 598268
rect 224178 598116 224274 598172
rect 224330 598116 224398 598172
rect 224454 598116 224522 598172
rect 224578 598116 224646 598172
rect 224702 598116 224798 598172
rect 224178 598048 224798 598116
rect 224178 597992 224274 598048
rect 224330 597992 224398 598048
rect 224454 597992 224522 598048
rect 224578 597992 224646 598048
rect 224702 597992 224798 598048
rect 224178 597924 224798 597992
rect 224178 597868 224274 597924
rect 224330 597868 224398 597924
rect 224454 597868 224522 597924
rect 224578 597868 224646 597924
rect 224702 597868 224798 597924
rect 224178 597800 224798 597868
rect 224178 597744 224274 597800
rect 224330 597744 224398 597800
rect 224454 597744 224522 597800
rect 224578 597744 224646 597800
rect 224702 597744 224798 597800
rect 224178 586350 224798 597744
rect 224178 586294 224274 586350
rect 224330 586294 224398 586350
rect 224454 586294 224522 586350
rect 224578 586294 224646 586350
rect 224702 586294 224798 586350
rect 224178 586226 224798 586294
rect 224178 586170 224274 586226
rect 224330 586170 224398 586226
rect 224454 586170 224522 586226
rect 224578 586170 224646 586226
rect 224702 586170 224798 586226
rect 224178 586102 224798 586170
rect 224178 586046 224274 586102
rect 224330 586046 224398 586102
rect 224454 586046 224522 586102
rect 224578 586046 224646 586102
rect 224702 586046 224798 586102
rect 224178 585978 224798 586046
rect 224178 585922 224274 585978
rect 224330 585922 224398 585978
rect 224454 585922 224522 585978
rect 224578 585922 224646 585978
rect 224702 585922 224798 585978
rect 224178 568350 224798 585922
rect 224178 568294 224274 568350
rect 224330 568294 224398 568350
rect 224454 568294 224522 568350
rect 224578 568294 224646 568350
rect 224702 568294 224798 568350
rect 224178 568226 224798 568294
rect 224178 568170 224274 568226
rect 224330 568170 224398 568226
rect 224454 568170 224522 568226
rect 224578 568170 224646 568226
rect 224702 568170 224798 568226
rect 224178 568102 224798 568170
rect 224178 568046 224274 568102
rect 224330 568046 224398 568102
rect 224454 568046 224522 568102
rect 224578 568046 224646 568102
rect 224702 568046 224798 568102
rect 224178 567978 224798 568046
rect 224178 567922 224274 567978
rect 224330 567922 224398 567978
rect 224454 567922 224522 567978
rect 224578 567922 224646 567978
rect 224702 567922 224798 567978
rect 224178 551870 224798 567922
rect 251178 597212 251798 598268
rect 251178 597156 251274 597212
rect 251330 597156 251398 597212
rect 251454 597156 251522 597212
rect 251578 597156 251646 597212
rect 251702 597156 251798 597212
rect 251178 597088 251798 597156
rect 251178 597032 251274 597088
rect 251330 597032 251398 597088
rect 251454 597032 251522 597088
rect 251578 597032 251646 597088
rect 251702 597032 251798 597088
rect 251178 596964 251798 597032
rect 251178 596908 251274 596964
rect 251330 596908 251398 596964
rect 251454 596908 251522 596964
rect 251578 596908 251646 596964
rect 251702 596908 251798 596964
rect 251178 596840 251798 596908
rect 251178 596784 251274 596840
rect 251330 596784 251398 596840
rect 251454 596784 251522 596840
rect 251578 596784 251646 596840
rect 251702 596784 251798 596840
rect 251178 580350 251798 596784
rect 251178 580294 251274 580350
rect 251330 580294 251398 580350
rect 251454 580294 251522 580350
rect 251578 580294 251646 580350
rect 251702 580294 251798 580350
rect 251178 580226 251798 580294
rect 251178 580170 251274 580226
rect 251330 580170 251398 580226
rect 251454 580170 251522 580226
rect 251578 580170 251646 580226
rect 251702 580170 251798 580226
rect 251178 580102 251798 580170
rect 251178 580046 251274 580102
rect 251330 580046 251398 580102
rect 251454 580046 251522 580102
rect 251578 580046 251646 580102
rect 251702 580046 251798 580102
rect 251178 579978 251798 580046
rect 251178 579922 251274 579978
rect 251330 579922 251398 579978
rect 251454 579922 251522 579978
rect 251578 579922 251646 579978
rect 251702 579922 251798 579978
rect 241168 562350 241488 562384
rect 241168 562294 241238 562350
rect 241294 562294 241362 562350
rect 241418 562294 241488 562350
rect 241168 562226 241488 562294
rect 241168 562170 241238 562226
rect 241294 562170 241362 562226
rect 241418 562170 241488 562226
rect 241168 562102 241488 562170
rect 241168 562046 241238 562102
rect 241294 562046 241362 562102
rect 241418 562046 241488 562102
rect 241168 561978 241488 562046
rect 241168 561922 241238 561978
rect 241294 561922 241362 561978
rect 241418 561922 241488 561978
rect 241168 561888 241488 561922
rect 251178 562350 251798 579922
rect 251178 562294 251274 562350
rect 251330 562294 251398 562350
rect 251454 562294 251522 562350
rect 251578 562294 251646 562350
rect 251702 562294 251798 562350
rect 251178 562226 251798 562294
rect 251178 562170 251274 562226
rect 251330 562170 251398 562226
rect 251454 562170 251522 562226
rect 251578 562170 251646 562226
rect 251702 562170 251798 562226
rect 251178 562102 251798 562170
rect 251178 562046 251274 562102
rect 251330 562046 251398 562102
rect 251454 562046 251522 562102
rect 251578 562046 251646 562102
rect 251702 562046 251798 562102
rect 251178 561978 251798 562046
rect 251178 561922 251274 561978
rect 251330 561922 251398 561978
rect 251454 561922 251522 561978
rect 251578 561922 251646 561978
rect 251702 561922 251798 561978
rect 225808 550350 226128 550384
rect 225808 550294 225878 550350
rect 225934 550294 226002 550350
rect 226058 550294 226128 550350
rect 225808 550226 226128 550294
rect 225808 550170 225878 550226
rect 225934 550170 226002 550226
rect 226058 550170 226128 550226
rect 225808 550102 226128 550170
rect 225808 550046 225878 550102
rect 225934 550046 226002 550102
rect 226058 550046 226128 550102
rect 225808 549978 226128 550046
rect 225808 549922 225878 549978
rect 225934 549922 226002 549978
rect 226058 549922 226128 549978
rect 225808 549888 226128 549922
rect 220458 544294 220554 544350
rect 220610 544294 220678 544350
rect 220734 544294 220802 544350
rect 220858 544294 220926 544350
rect 220982 544294 221078 544350
rect 220458 544226 221078 544294
rect 220458 544170 220554 544226
rect 220610 544170 220678 544226
rect 220734 544170 220802 544226
rect 220858 544170 220926 544226
rect 220982 544170 221078 544226
rect 220458 544102 221078 544170
rect 220458 544046 220554 544102
rect 220610 544046 220678 544102
rect 220734 544046 220802 544102
rect 220858 544046 220926 544102
rect 220982 544046 221078 544102
rect 220458 543978 221078 544046
rect 241168 544350 241488 544384
rect 241168 544294 241238 544350
rect 241294 544294 241362 544350
rect 241418 544294 241488 544350
rect 241168 544226 241488 544294
rect 241168 544170 241238 544226
rect 241294 544170 241362 544226
rect 241418 544170 241488 544226
rect 241168 544102 241488 544170
rect 241168 544046 241238 544102
rect 241294 544046 241362 544102
rect 241418 544046 241488 544102
rect 220458 543922 220554 543978
rect 220610 543922 220678 543978
rect 220734 543922 220802 543978
rect 220858 543922 220926 543978
rect 220982 543922 221078 543978
rect 205772 529890 205828 529900
rect 205996 530292 206052 530302
rect 205996 520996 206052 530236
rect 205996 520930 206052 520940
rect 220458 526350 221078 543922
rect 220458 526294 220554 526350
rect 220610 526294 220678 526350
rect 220734 526294 220802 526350
rect 220858 526294 220926 526350
rect 220982 526294 221078 526350
rect 220458 526226 221078 526294
rect 220458 526170 220554 526226
rect 220610 526170 220678 526226
rect 220734 526170 220802 526226
rect 220858 526170 220926 526226
rect 220982 526170 221078 526226
rect 220458 526102 221078 526170
rect 220458 526046 220554 526102
rect 220610 526046 220678 526102
rect 220734 526046 220802 526102
rect 220858 526046 220926 526102
rect 220982 526046 221078 526102
rect 220458 525978 221078 526046
rect 220458 525922 220554 525978
rect 220610 525922 220678 525978
rect 220734 525922 220802 525978
rect 220858 525922 220926 525978
rect 220982 525922 221078 525978
rect 204092 496850 204148 496860
rect 220458 508350 221078 525922
rect 220458 508294 220554 508350
rect 220610 508294 220678 508350
rect 220734 508294 220802 508350
rect 220858 508294 220926 508350
rect 220982 508294 221078 508350
rect 220458 508226 221078 508294
rect 220458 508170 220554 508226
rect 220610 508170 220678 508226
rect 220734 508170 220802 508226
rect 220858 508170 220926 508226
rect 220982 508170 221078 508226
rect 220458 508102 221078 508170
rect 220458 508046 220554 508102
rect 220610 508046 220678 508102
rect 220734 508046 220802 508102
rect 220858 508046 220926 508102
rect 220982 508046 221078 508102
rect 220458 507978 221078 508046
rect 220458 507922 220554 507978
rect 220610 507922 220678 507978
rect 220734 507922 220802 507978
rect 220858 507922 220926 507978
rect 220982 507922 221078 507978
rect 210448 490350 210768 490384
rect 210448 490294 210518 490350
rect 210574 490294 210642 490350
rect 210698 490294 210768 490350
rect 210448 490226 210768 490294
rect 210448 490170 210518 490226
rect 210574 490170 210642 490226
rect 210698 490170 210768 490226
rect 210448 490102 210768 490170
rect 210448 490046 210518 490102
rect 210574 490046 210642 490102
rect 210698 490046 210768 490102
rect 210448 489978 210768 490046
rect 210448 489922 210518 489978
rect 210574 489922 210642 489978
rect 210698 489922 210768 489978
rect 210448 489888 210768 489922
rect 220458 490350 221078 507922
rect 220458 490294 220554 490350
rect 220610 490294 220678 490350
rect 220734 490294 220802 490350
rect 220858 490294 220926 490350
rect 220982 490294 221078 490350
rect 220458 490226 221078 490294
rect 220458 490170 220554 490226
rect 220610 490170 220678 490226
rect 220734 490170 220802 490226
rect 220858 490170 220926 490226
rect 220982 490170 221078 490226
rect 220458 490102 221078 490170
rect 220458 490046 220554 490102
rect 220610 490046 220678 490102
rect 220734 490046 220802 490102
rect 220858 490046 220926 490102
rect 220982 490046 221078 490102
rect 220458 489978 221078 490046
rect 220458 489922 220554 489978
rect 220610 489922 220678 489978
rect 220734 489922 220802 489978
rect 220858 489922 220926 489978
rect 220982 489922 221078 489978
rect 201628 483364 201684 483374
rect 201628 483058 201684 483308
rect 201628 482992 201684 483002
rect 206668 482356 206724 482376
rect 206668 482272 206724 482282
rect 203196 481348 203252 481358
rect 203196 442036 203252 481292
rect 204204 479332 204260 479342
rect 203196 441970 203252 441980
rect 204092 467908 204148 467918
rect 204092 433636 204148 467852
rect 204204 458836 204260 479276
rect 206556 478660 206612 478670
rect 206556 474598 206612 478604
rect 206556 474532 206612 474542
rect 210448 472350 210768 472384
rect 210448 472294 210518 472350
rect 210574 472294 210642 472350
rect 210698 472294 210768 472350
rect 210448 472226 210768 472294
rect 210448 472170 210518 472226
rect 210574 472170 210642 472226
rect 210698 472170 210768 472226
rect 210448 472102 210768 472170
rect 210448 472046 210518 472102
rect 210574 472046 210642 472102
rect 210698 472046 210768 472102
rect 210448 471978 210768 472046
rect 210448 471922 210518 471978
rect 210574 471922 210642 471978
rect 210698 471922 210768 471978
rect 210448 471888 210768 471922
rect 220458 472350 221078 489922
rect 224178 532350 224798 543986
rect 241168 543978 241488 544046
rect 241168 543922 241238 543978
rect 241294 543922 241362 543978
rect 241418 543922 241488 543978
rect 241168 543888 241488 543922
rect 251178 544350 251798 561922
rect 254898 598172 255518 598268
rect 254898 598116 254994 598172
rect 255050 598116 255118 598172
rect 255174 598116 255242 598172
rect 255298 598116 255366 598172
rect 255422 598116 255518 598172
rect 254898 598048 255518 598116
rect 254898 597992 254994 598048
rect 255050 597992 255118 598048
rect 255174 597992 255242 598048
rect 255298 597992 255366 598048
rect 255422 597992 255518 598048
rect 254898 597924 255518 597992
rect 254898 597868 254994 597924
rect 255050 597868 255118 597924
rect 255174 597868 255242 597924
rect 255298 597868 255366 597924
rect 255422 597868 255518 597924
rect 254898 597800 255518 597868
rect 254898 597744 254994 597800
rect 255050 597744 255118 597800
rect 255174 597744 255242 597800
rect 255298 597744 255366 597800
rect 255422 597744 255518 597800
rect 254898 586350 255518 597744
rect 254898 586294 254994 586350
rect 255050 586294 255118 586350
rect 255174 586294 255242 586350
rect 255298 586294 255366 586350
rect 255422 586294 255518 586350
rect 254898 586226 255518 586294
rect 254898 586170 254994 586226
rect 255050 586170 255118 586226
rect 255174 586170 255242 586226
rect 255298 586170 255366 586226
rect 255422 586170 255518 586226
rect 254898 586102 255518 586170
rect 254898 586046 254994 586102
rect 255050 586046 255118 586102
rect 255174 586046 255242 586102
rect 255298 586046 255366 586102
rect 255422 586046 255518 586102
rect 254898 585978 255518 586046
rect 254898 585922 254994 585978
rect 255050 585922 255118 585978
rect 255174 585922 255242 585978
rect 255298 585922 255366 585978
rect 255422 585922 255518 585978
rect 254898 568350 255518 585922
rect 281898 597212 282518 598268
rect 281898 597156 281994 597212
rect 282050 597156 282118 597212
rect 282174 597156 282242 597212
rect 282298 597156 282366 597212
rect 282422 597156 282518 597212
rect 281898 597088 282518 597156
rect 281898 597032 281994 597088
rect 282050 597032 282118 597088
rect 282174 597032 282242 597088
rect 282298 597032 282366 597088
rect 282422 597032 282518 597088
rect 281898 596964 282518 597032
rect 281898 596908 281994 596964
rect 282050 596908 282118 596964
rect 282174 596908 282242 596964
rect 282298 596908 282366 596964
rect 282422 596908 282518 596964
rect 281898 596840 282518 596908
rect 281898 596784 281994 596840
rect 282050 596784 282118 596840
rect 282174 596784 282242 596840
rect 282298 596784 282366 596840
rect 282422 596784 282518 596840
rect 281898 580350 282518 596784
rect 281898 580294 281994 580350
rect 282050 580294 282118 580350
rect 282174 580294 282242 580350
rect 282298 580294 282366 580350
rect 282422 580294 282518 580350
rect 281898 580226 282518 580294
rect 281898 580170 281994 580226
rect 282050 580170 282118 580226
rect 282174 580170 282242 580226
rect 282298 580170 282366 580226
rect 282422 580170 282518 580226
rect 281898 580102 282518 580170
rect 281898 580046 281994 580102
rect 282050 580046 282118 580102
rect 282174 580046 282242 580102
rect 282298 580046 282366 580102
rect 282422 580046 282518 580102
rect 281898 579978 282518 580046
rect 281898 579922 281994 579978
rect 282050 579922 282118 579978
rect 282174 579922 282242 579978
rect 282298 579922 282366 579978
rect 282422 579922 282518 579978
rect 254898 568294 254994 568350
rect 255050 568294 255118 568350
rect 255174 568294 255242 568350
rect 255298 568294 255366 568350
rect 255422 568294 255518 568350
rect 254898 568226 255518 568294
rect 254898 568170 254994 568226
rect 255050 568170 255118 568226
rect 255174 568170 255242 568226
rect 255298 568170 255366 568226
rect 255422 568170 255518 568226
rect 254898 568102 255518 568170
rect 254898 568046 254994 568102
rect 255050 568046 255118 568102
rect 255174 568046 255242 568102
rect 255298 568046 255366 568102
rect 255422 568046 255518 568102
rect 254898 567978 255518 568046
rect 254898 567922 254994 567978
rect 255050 567922 255118 567978
rect 255174 567922 255242 567978
rect 255298 567922 255366 567978
rect 255422 567922 255518 567978
rect 252812 553924 252868 553934
rect 251178 544294 251274 544350
rect 251330 544294 251398 544350
rect 251454 544294 251522 544350
rect 251578 544294 251646 544350
rect 251702 544294 251798 544350
rect 251178 544226 251798 544294
rect 251178 544170 251274 544226
rect 251330 544170 251398 544226
rect 251454 544170 251522 544226
rect 251578 544170 251646 544226
rect 251702 544170 251798 544226
rect 251178 544102 251798 544170
rect 251178 544046 251274 544102
rect 251330 544046 251398 544102
rect 251454 544046 251522 544102
rect 251578 544046 251646 544102
rect 251702 544046 251798 544102
rect 251178 543978 251798 544046
rect 251178 543922 251274 543978
rect 251330 543922 251398 543978
rect 251454 543922 251522 543978
rect 251578 543922 251646 543978
rect 251702 543922 251798 543978
rect 224178 532294 224274 532350
rect 224330 532294 224398 532350
rect 224454 532294 224522 532350
rect 224578 532294 224646 532350
rect 224702 532294 224798 532350
rect 224178 532226 224798 532294
rect 224178 532170 224274 532226
rect 224330 532170 224398 532226
rect 224454 532170 224522 532226
rect 224578 532170 224646 532226
rect 224702 532170 224798 532226
rect 224178 532102 224798 532170
rect 224178 532046 224274 532102
rect 224330 532046 224398 532102
rect 224454 532046 224522 532102
rect 224578 532046 224646 532102
rect 224702 532046 224798 532102
rect 224178 531978 224798 532046
rect 224178 531922 224274 531978
rect 224330 531922 224398 531978
rect 224454 531922 224522 531978
rect 224578 531922 224646 531978
rect 224702 531922 224798 531978
rect 224178 514350 224798 531922
rect 225808 532350 226128 532384
rect 225808 532294 225878 532350
rect 225934 532294 226002 532350
rect 226058 532294 226128 532350
rect 225808 532226 226128 532294
rect 225808 532170 225878 532226
rect 225934 532170 226002 532226
rect 226058 532170 226128 532226
rect 225808 532102 226128 532170
rect 225808 532046 225878 532102
rect 225934 532046 226002 532102
rect 226058 532046 226128 532102
rect 225808 531978 226128 532046
rect 225808 531922 225878 531978
rect 225934 531922 226002 531978
rect 226058 531922 226128 531978
rect 225808 531888 226128 531922
rect 249452 526708 249508 526718
rect 224178 514294 224274 514350
rect 224330 514294 224398 514350
rect 224454 514294 224522 514350
rect 224578 514294 224646 514350
rect 224702 514294 224798 514350
rect 224178 514226 224798 514294
rect 224178 514170 224274 514226
rect 224330 514170 224398 514226
rect 224454 514170 224522 514226
rect 224578 514170 224646 514226
rect 224702 514170 224798 514226
rect 224178 514102 224798 514170
rect 224178 514046 224274 514102
rect 224330 514046 224398 514102
rect 224454 514046 224522 514102
rect 224578 514046 224646 514102
rect 224702 514046 224798 514102
rect 224178 513978 224798 514046
rect 224178 513922 224274 513978
rect 224330 513922 224398 513978
rect 224454 513922 224522 513978
rect 224578 513922 224646 513978
rect 224702 513922 224798 513978
rect 224178 496350 224798 513922
rect 224178 496294 224274 496350
rect 224330 496294 224398 496350
rect 224454 496294 224522 496350
rect 224578 496294 224646 496350
rect 224702 496294 224798 496350
rect 224178 496226 224798 496294
rect 224178 496170 224274 496226
rect 224330 496170 224398 496226
rect 224454 496170 224522 496226
rect 224578 496170 224646 496226
rect 224702 496170 224798 496226
rect 224178 496102 224798 496170
rect 224178 496046 224274 496102
rect 224330 496046 224398 496102
rect 224454 496046 224522 496102
rect 224578 496046 224646 496102
rect 224702 496046 224798 496102
rect 224178 495978 224798 496046
rect 224178 495922 224274 495978
rect 224330 495922 224398 495978
rect 224454 495922 224522 495978
rect 224578 495922 224646 495978
rect 224702 495922 224798 495978
rect 224178 483918 224798 495922
rect 246092 523572 246148 523582
rect 246092 495236 246148 523516
rect 247772 520100 247828 520110
rect 246876 501508 246932 501518
rect 246876 497588 246932 501452
rect 246876 497522 246932 497532
rect 246092 495170 246148 495180
rect 241168 490350 241488 490384
rect 241168 490294 241238 490350
rect 241294 490294 241362 490350
rect 241418 490294 241488 490350
rect 241168 490226 241488 490294
rect 241168 490170 241238 490226
rect 241294 490170 241362 490226
rect 241418 490170 241488 490226
rect 241168 490102 241488 490170
rect 241168 490046 241238 490102
rect 241294 490046 241362 490102
rect 241418 490046 241488 490102
rect 241168 489978 241488 490046
rect 241168 489922 241238 489978
rect 241294 489922 241362 489978
rect 241418 489922 241488 489978
rect 241168 489888 241488 489922
rect 247772 486836 247828 520044
rect 247884 511700 247940 511710
rect 247884 492996 247940 511644
rect 247884 492930 247940 492940
rect 247996 506772 248052 506782
rect 247996 490756 248052 506716
rect 247996 490690 248052 490700
rect 247772 486770 247828 486780
rect 249452 484596 249508 526652
rect 249452 484530 249508 484540
rect 251178 526350 251798 543922
rect 251178 526294 251274 526350
rect 251330 526294 251398 526350
rect 251454 526294 251522 526350
rect 251578 526294 251646 526350
rect 251702 526294 251798 526350
rect 251178 526226 251798 526294
rect 251178 526170 251274 526226
rect 251330 526170 251398 526226
rect 251454 526170 251522 526226
rect 251578 526170 251646 526226
rect 251702 526170 251798 526226
rect 251178 526102 251798 526170
rect 251178 526046 251274 526102
rect 251330 526046 251398 526102
rect 251454 526046 251522 526102
rect 251578 526046 251646 526102
rect 251702 526046 251798 526102
rect 251178 525978 251798 526046
rect 251178 525922 251274 525978
rect 251330 525922 251398 525978
rect 251454 525922 251522 525978
rect 251578 525922 251646 525978
rect 251702 525922 251798 525978
rect 251178 508350 251798 525922
rect 251916 547204 251972 547214
rect 251916 524356 251972 547148
rect 252812 533428 252868 553868
rect 254898 550350 255518 567922
rect 270284 568932 270340 568942
rect 270284 567812 270340 568876
rect 270284 567746 270340 567756
rect 271404 568932 271460 568942
rect 271404 567028 271460 568876
rect 272524 568932 272580 568942
rect 272524 567588 272580 568876
rect 272524 567522 272580 567532
rect 281898 567214 282518 579922
rect 285618 598172 286238 598268
rect 285618 598116 285714 598172
rect 285770 598116 285838 598172
rect 285894 598116 285962 598172
rect 286018 598116 286086 598172
rect 286142 598116 286238 598172
rect 285618 598048 286238 598116
rect 285618 597992 285714 598048
rect 285770 597992 285838 598048
rect 285894 597992 285962 598048
rect 286018 597992 286086 598048
rect 286142 597992 286238 598048
rect 285618 597924 286238 597992
rect 285618 597868 285714 597924
rect 285770 597868 285838 597924
rect 285894 597868 285962 597924
rect 286018 597868 286086 597924
rect 286142 597868 286238 597924
rect 285618 597800 286238 597868
rect 285618 597744 285714 597800
rect 285770 597744 285838 597800
rect 285894 597744 285962 597800
rect 286018 597744 286086 597800
rect 286142 597744 286238 597800
rect 285618 586350 286238 597744
rect 285618 586294 285714 586350
rect 285770 586294 285838 586350
rect 285894 586294 285962 586350
rect 286018 586294 286086 586350
rect 286142 586294 286238 586350
rect 285618 586226 286238 586294
rect 285618 586170 285714 586226
rect 285770 586170 285838 586226
rect 285894 586170 285962 586226
rect 286018 586170 286086 586226
rect 286142 586170 286238 586226
rect 285618 586102 286238 586170
rect 285618 586046 285714 586102
rect 285770 586046 285838 586102
rect 285894 586046 285962 586102
rect 286018 586046 286086 586102
rect 286142 586046 286238 586102
rect 285618 585978 286238 586046
rect 285618 585922 285714 585978
rect 285770 585922 285838 585978
rect 285894 585922 285962 585978
rect 286018 585922 286086 585978
rect 286142 585922 286238 585978
rect 285618 568350 286238 585922
rect 312618 597212 313238 598268
rect 312618 597156 312714 597212
rect 312770 597156 312838 597212
rect 312894 597156 312962 597212
rect 313018 597156 313086 597212
rect 313142 597156 313238 597212
rect 312618 597088 313238 597156
rect 312618 597032 312714 597088
rect 312770 597032 312838 597088
rect 312894 597032 312962 597088
rect 313018 597032 313086 597088
rect 313142 597032 313238 597088
rect 312618 596964 313238 597032
rect 312618 596908 312714 596964
rect 312770 596908 312838 596964
rect 312894 596908 312962 596964
rect 313018 596908 313086 596964
rect 313142 596908 313238 596964
rect 312618 596840 313238 596908
rect 312618 596784 312714 596840
rect 312770 596784 312838 596840
rect 312894 596784 312962 596840
rect 313018 596784 313086 596840
rect 313142 596784 313238 596840
rect 312618 580350 313238 596784
rect 312618 580294 312714 580350
rect 312770 580294 312838 580350
rect 312894 580294 312962 580350
rect 313018 580294 313086 580350
rect 313142 580294 313238 580350
rect 312618 580226 313238 580294
rect 312618 580170 312714 580226
rect 312770 580170 312838 580226
rect 312894 580170 312962 580226
rect 313018 580170 313086 580226
rect 313142 580170 313238 580226
rect 312618 580102 313238 580170
rect 312618 580046 312714 580102
rect 312770 580046 312838 580102
rect 312894 580046 312962 580102
rect 313018 580046 313086 580102
rect 313142 580046 313238 580102
rect 312618 579978 313238 580046
rect 312618 579922 312714 579978
rect 312770 579922 312838 579978
rect 312894 579922 312962 579978
rect 313018 579922 313086 579978
rect 313142 579922 313238 579978
rect 290444 569828 290500 569838
rect 290444 569638 290500 569772
rect 290444 569572 290500 569582
rect 303660 569604 303716 569614
rect 285618 568294 285714 568350
rect 285770 568294 285838 568350
rect 285894 568294 285962 568350
rect 286018 568294 286086 568350
rect 286142 568294 286238 568350
rect 285618 568226 286238 568294
rect 285618 568170 285714 568226
rect 285770 568170 285838 568226
rect 285894 568170 285962 568226
rect 286018 568170 286086 568226
rect 286142 568170 286238 568226
rect 285618 568102 286238 568170
rect 285618 568046 285714 568102
rect 285770 568046 285838 568102
rect 285894 568046 285962 568102
rect 286018 568046 286086 568102
rect 286142 568046 286238 568102
rect 285618 567978 286238 568046
rect 285618 567922 285714 567978
rect 285770 567922 285838 567978
rect 285894 567922 285962 567978
rect 286018 567922 286086 567978
rect 286142 567922 286238 567978
rect 285618 567214 286238 567922
rect 289324 568932 289380 568942
rect 271404 566962 271460 566972
rect 289324 566938 289380 568876
rect 300524 568932 300580 568942
rect 300524 567700 300580 568876
rect 300524 567634 300580 567644
rect 301644 568932 301700 568942
rect 301644 567364 301700 568876
rect 302764 568932 302820 568942
rect 302764 568708 302820 568876
rect 302764 568642 302820 568652
rect 303660 567476 303716 569548
rect 303660 567410 303716 567420
rect 301644 567298 301700 567308
rect 312618 567214 313238 579922
rect 316338 598172 316958 598268
rect 316338 598116 316434 598172
rect 316490 598116 316558 598172
rect 316614 598116 316682 598172
rect 316738 598116 316806 598172
rect 316862 598116 316958 598172
rect 316338 598048 316958 598116
rect 316338 597992 316434 598048
rect 316490 597992 316558 598048
rect 316614 597992 316682 598048
rect 316738 597992 316806 598048
rect 316862 597992 316958 598048
rect 316338 597924 316958 597992
rect 316338 597868 316434 597924
rect 316490 597868 316558 597924
rect 316614 597868 316682 597924
rect 316738 597868 316806 597924
rect 316862 597868 316958 597924
rect 316338 597800 316958 597868
rect 316338 597744 316434 597800
rect 316490 597744 316558 597800
rect 316614 597744 316682 597800
rect 316738 597744 316806 597800
rect 316862 597744 316958 597800
rect 316338 586350 316958 597744
rect 316338 586294 316434 586350
rect 316490 586294 316558 586350
rect 316614 586294 316682 586350
rect 316738 586294 316806 586350
rect 316862 586294 316958 586350
rect 316338 586226 316958 586294
rect 316338 586170 316434 586226
rect 316490 586170 316558 586226
rect 316614 586170 316682 586226
rect 316738 586170 316806 586226
rect 316862 586170 316958 586226
rect 316338 586102 316958 586170
rect 316338 586046 316434 586102
rect 316490 586046 316558 586102
rect 316614 586046 316682 586102
rect 316738 586046 316806 586102
rect 316862 586046 316958 586102
rect 316338 585978 316958 586046
rect 316338 585922 316434 585978
rect 316490 585922 316558 585978
rect 316614 585922 316682 585978
rect 316738 585922 316806 585978
rect 316862 585922 316958 585978
rect 315756 569604 315812 569614
rect 315756 567252 315812 569548
rect 316338 568350 316958 585922
rect 343338 597212 343958 598268
rect 343338 597156 343434 597212
rect 343490 597156 343558 597212
rect 343614 597156 343682 597212
rect 343738 597156 343806 597212
rect 343862 597156 343958 597212
rect 343338 597088 343958 597156
rect 343338 597032 343434 597088
rect 343490 597032 343558 597088
rect 343614 597032 343682 597088
rect 343738 597032 343806 597088
rect 343862 597032 343958 597088
rect 343338 596964 343958 597032
rect 343338 596908 343434 596964
rect 343490 596908 343558 596964
rect 343614 596908 343682 596964
rect 343738 596908 343806 596964
rect 343862 596908 343958 596964
rect 343338 596840 343958 596908
rect 343338 596784 343434 596840
rect 343490 596784 343558 596840
rect 343614 596784 343682 596840
rect 343738 596784 343806 596840
rect 343862 596784 343958 596840
rect 343338 580350 343958 596784
rect 343338 580294 343434 580350
rect 343490 580294 343558 580350
rect 343614 580294 343682 580350
rect 343738 580294 343806 580350
rect 343862 580294 343958 580350
rect 343338 580226 343958 580294
rect 343338 580170 343434 580226
rect 343490 580170 343558 580226
rect 343614 580170 343682 580226
rect 343738 580170 343806 580226
rect 343862 580170 343958 580226
rect 343338 580102 343958 580170
rect 343338 580046 343434 580102
rect 343490 580046 343558 580102
rect 343614 580046 343682 580102
rect 343738 580046 343806 580102
rect 343862 580046 343958 580102
rect 343338 579978 343958 580046
rect 343338 579922 343434 579978
rect 343490 579922 343558 579978
rect 343614 579922 343682 579978
rect 343738 579922 343806 579978
rect 343862 579922 343958 579978
rect 319116 571284 319172 571294
rect 317996 570052 318052 570062
rect 317996 569380 318052 569996
rect 317996 569314 318052 569324
rect 316338 568294 316434 568350
rect 316490 568294 316558 568350
rect 316614 568294 316682 568350
rect 316738 568294 316806 568350
rect 316862 568294 316958 568350
rect 316338 568226 316958 568294
rect 316338 568170 316434 568226
rect 316490 568170 316558 568226
rect 316614 568170 316682 568226
rect 316738 568170 316806 568226
rect 316862 568170 316958 568226
rect 316338 568102 316958 568170
rect 316338 568046 316434 568102
rect 316490 568046 316558 568102
rect 316614 568046 316682 568102
rect 316738 568046 316806 568102
rect 316862 568046 316958 568102
rect 316338 567978 316958 568046
rect 316338 567922 316434 567978
rect 316490 567922 316558 567978
rect 316614 567922 316682 567978
rect 316738 567922 316806 567978
rect 316862 567922 316958 567978
rect 316338 567214 316958 567922
rect 315756 567186 315812 567196
rect 319116 567140 319172 571228
rect 330764 571284 330820 571296
rect 330764 571192 330820 571202
rect 319116 567074 319172 567084
rect 333452 569638 333508 569648
rect 289324 566872 289380 566882
rect 272448 562350 272768 562384
rect 272448 562294 272518 562350
rect 272574 562294 272642 562350
rect 272698 562294 272768 562350
rect 272448 562226 272768 562294
rect 272448 562170 272518 562226
rect 272574 562170 272642 562226
rect 272698 562170 272768 562226
rect 272448 562102 272768 562170
rect 272448 562046 272518 562102
rect 272574 562046 272642 562102
rect 272698 562046 272768 562102
rect 272448 561978 272768 562046
rect 272448 561922 272518 561978
rect 272574 561922 272642 561978
rect 272698 561922 272768 561978
rect 272448 561888 272768 561922
rect 303168 562350 303488 562384
rect 303168 562294 303238 562350
rect 303294 562294 303362 562350
rect 303418 562294 303488 562350
rect 303168 562226 303488 562294
rect 303168 562170 303238 562226
rect 303294 562170 303362 562226
rect 303418 562170 303488 562226
rect 303168 562102 303488 562170
rect 303168 562046 303238 562102
rect 303294 562046 303362 562102
rect 303418 562046 303488 562102
rect 303168 561978 303488 562046
rect 303168 561922 303238 561978
rect 303294 561922 303362 561978
rect 303418 561922 303488 561978
rect 303168 561888 303488 561922
rect 254898 550294 254994 550350
rect 255050 550294 255118 550350
rect 255174 550294 255242 550350
rect 255298 550294 255366 550350
rect 255422 550294 255518 550350
rect 254898 550226 255518 550294
rect 254898 550170 254994 550226
rect 255050 550170 255118 550226
rect 255174 550170 255242 550226
rect 255298 550170 255366 550226
rect 255422 550170 255518 550226
rect 254898 550102 255518 550170
rect 254898 550046 254994 550102
rect 255050 550046 255118 550102
rect 255174 550046 255242 550102
rect 255298 550046 255366 550102
rect 255422 550046 255518 550102
rect 254898 549978 255518 550046
rect 254898 549922 254994 549978
rect 255050 549922 255118 549978
rect 255174 549922 255242 549978
rect 255298 549922 255366 549978
rect 255422 549922 255518 549978
rect 252812 533362 252868 533372
rect 254492 545860 254548 545870
rect 254492 531636 254548 545804
rect 254492 531570 254548 531580
rect 254898 532350 255518 549922
rect 261324 552580 261380 552590
rect 257852 548548 257908 548558
rect 254898 532294 254994 532350
rect 255050 532294 255118 532350
rect 255174 532294 255242 532350
rect 255298 532294 255366 532350
rect 255422 532294 255518 532350
rect 254898 532226 255518 532294
rect 254898 532170 254994 532226
rect 255050 532170 255118 532226
rect 255174 532170 255242 532226
rect 255298 532170 255366 532226
rect 255422 532170 255518 532226
rect 254898 532102 255518 532170
rect 254898 532046 254994 532102
rect 255050 532046 255118 532102
rect 255174 532046 255242 532102
rect 255298 532046 255366 532102
rect 255422 532046 255518 532102
rect 254898 531978 255518 532046
rect 254898 531922 254994 531978
rect 255050 531922 255118 531978
rect 255174 531922 255242 531978
rect 255298 531922 255366 531978
rect 255422 531922 255518 531978
rect 251916 524290 251972 524300
rect 252812 528052 252868 528062
rect 251178 508294 251274 508350
rect 251330 508294 251398 508350
rect 251454 508294 251522 508350
rect 251578 508294 251646 508350
rect 251702 508294 251798 508350
rect 251178 508226 251798 508294
rect 251178 508170 251274 508226
rect 251330 508170 251398 508226
rect 251454 508170 251522 508226
rect 251578 508170 251646 508226
rect 251702 508170 251798 508226
rect 251178 508102 251798 508170
rect 251178 508046 251274 508102
rect 251330 508046 251398 508102
rect 251454 508046 251522 508102
rect 251578 508046 251646 508102
rect 251702 508046 251798 508102
rect 251178 507978 251798 508046
rect 251178 507922 251274 507978
rect 251330 507922 251398 507978
rect 251454 507922 251522 507978
rect 251578 507922 251646 507978
rect 251702 507922 251798 507978
rect 251178 490350 251798 507922
rect 251178 490294 251274 490350
rect 251330 490294 251398 490350
rect 251454 490294 251522 490350
rect 251578 490294 251646 490350
rect 251702 490294 251798 490350
rect 251178 490226 251798 490294
rect 251178 490170 251274 490226
rect 251330 490170 251398 490226
rect 251454 490170 251522 490226
rect 251578 490170 251646 490226
rect 251702 490170 251798 490226
rect 251178 490102 251798 490170
rect 251178 490046 251274 490102
rect 251330 490046 251398 490102
rect 251454 490046 251522 490102
rect 251578 490046 251646 490102
rect 251702 490046 251798 490102
rect 251178 489978 251798 490046
rect 251178 489922 251274 489978
rect 251330 489922 251398 489978
rect 251454 489922 251522 489978
rect 251578 489922 251646 489978
rect 251702 489922 251798 489978
rect 247996 482338 248052 482348
rect 225808 478350 226128 478384
rect 225808 478294 225878 478350
rect 225934 478294 226002 478350
rect 226058 478294 226128 478350
rect 225808 478226 226128 478294
rect 225808 478170 225878 478226
rect 225934 478170 226002 478226
rect 226058 478170 226128 478226
rect 225808 478102 226128 478170
rect 225808 478046 225878 478102
rect 225934 478046 226002 478102
rect 226058 478046 226128 478102
rect 225808 477978 226128 478046
rect 225808 477922 225878 477978
rect 225934 477922 226002 477978
rect 226058 477922 226128 477978
rect 225808 477888 226128 477922
rect 223356 474598 223412 474608
rect 223356 473698 223412 474542
rect 223356 473632 223412 473642
rect 220458 472294 220554 472350
rect 220610 472294 220678 472350
rect 220734 472294 220802 472350
rect 220858 472294 220926 472350
rect 220982 472294 221078 472350
rect 220458 472226 221078 472294
rect 220458 472170 220554 472226
rect 220610 472170 220678 472226
rect 220734 472170 220802 472226
rect 220858 472170 220926 472226
rect 220982 472170 221078 472226
rect 220458 472102 221078 472170
rect 220458 472046 220554 472102
rect 220610 472046 220678 472102
rect 220734 472046 220802 472102
rect 220858 472046 220926 472102
rect 220982 472046 221078 472102
rect 220458 471978 221078 472046
rect 220458 471922 220554 471978
rect 220610 471922 220678 471978
rect 220734 471922 220802 471978
rect 220858 471922 220926 471978
rect 220982 471922 221078 471978
rect 204204 458770 204260 458780
rect 205772 461188 205828 461198
rect 205772 434756 205828 461132
rect 205772 434690 205828 434700
rect 220458 454350 221078 471922
rect 220458 454294 220554 454350
rect 220610 454294 220678 454350
rect 220734 454294 220802 454350
rect 220858 454294 220926 454350
rect 220982 454294 221078 454350
rect 220458 454226 221078 454294
rect 220458 454170 220554 454226
rect 220610 454170 220678 454226
rect 220734 454170 220802 454226
rect 220858 454170 220926 454226
rect 220982 454170 221078 454226
rect 220458 454102 221078 454170
rect 220458 454046 220554 454102
rect 220610 454046 220678 454102
rect 220734 454046 220802 454102
rect 220858 454046 220926 454102
rect 220982 454046 221078 454102
rect 220458 453978 221078 454046
rect 220458 453922 220554 453978
rect 220610 453922 220678 453978
rect 220734 453922 220802 453978
rect 220858 453922 220926 453978
rect 220982 453922 221078 453978
rect 220458 436350 221078 453922
rect 220458 436294 220554 436350
rect 220610 436294 220678 436350
rect 220734 436294 220802 436350
rect 220858 436294 220926 436350
rect 220982 436294 221078 436350
rect 220458 436226 221078 436294
rect 220458 436170 220554 436226
rect 220610 436170 220678 436226
rect 220734 436170 220802 436226
rect 220858 436170 220926 436226
rect 220982 436170 221078 436226
rect 220458 436102 221078 436170
rect 220458 436046 220554 436102
rect 220610 436046 220678 436102
rect 220734 436046 220802 436102
rect 220858 436046 220926 436102
rect 220982 436046 221078 436102
rect 220458 435978 221078 436046
rect 220458 435922 220554 435978
rect 220610 435922 220678 435978
rect 220734 435922 220802 435978
rect 220858 435922 220926 435978
rect 220982 435922 221078 435978
rect 204092 433570 204148 433580
rect 210448 418350 210768 418384
rect 210448 418294 210518 418350
rect 210574 418294 210642 418350
rect 210698 418294 210768 418350
rect 210448 418226 210768 418294
rect 210448 418170 210518 418226
rect 210574 418170 210642 418226
rect 210698 418170 210768 418226
rect 210448 418102 210768 418170
rect 210448 418046 210518 418102
rect 210574 418046 210642 418102
rect 210698 418046 210768 418102
rect 210448 417978 210768 418046
rect 210448 417922 210518 417978
rect 210574 417922 210642 417978
rect 210698 417922 210768 417978
rect 210448 417888 210768 417922
rect 220458 418350 221078 435922
rect 224178 460350 224798 473122
rect 241168 472350 241488 472384
rect 241168 472294 241238 472350
rect 241294 472294 241362 472350
rect 241418 472294 241488 472350
rect 241168 472226 241488 472294
rect 241168 472170 241238 472226
rect 241294 472170 241362 472226
rect 241418 472170 241488 472226
rect 241168 472102 241488 472170
rect 241168 472046 241238 472102
rect 241294 472046 241362 472102
rect 241418 472046 241488 472102
rect 241168 471978 241488 472046
rect 241168 471922 241238 471978
rect 241294 471922 241362 471978
rect 241418 471922 241488 471978
rect 241168 471888 241488 471922
rect 247996 471716 248052 482282
rect 251020 478660 251076 478670
rect 250908 477988 250964 477998
rect 250908 474852 250964 477932
rect 251020 476308 251076 478604
rect 251020 476242 251076 476252
rect 250908 474786 250964 474796
rect 247996 471650 248052 471660
rect 249452 473878 249508 473888
rect 249452 466228 249508 473822
rect 249452 466162 249508 466172
rect 251178 472350 251798 489922
rect 251916 503300 251972 503310
rect 251916 487396 251972 503244
rect 251916 487330 251972 487340
rect 252812 483476 252868 527996
rect 252812 483410 252868 483420
rect 254898 514350 255518 531922
rect 256284 544516 256340 544526
rect 254898 514294 254994 514350
rect 255050 514294 255118 514350
rect 255174 514294 255242 514350
rect 255298 514294 255366 514350
rect 255422 514294 255518 514350
rect 254898 514226 255518 514294
rect 254898 514170 254994 514226
rect 255050 514170 255118 514226
rect 255174 514170 255242 514226
rect 255298 514170 255366 514226
rect 255422 514170 255518 514226
rect 254898 514102 255518 514170
rect 254898 514046 254994 514102
rect 255050 514046 255118 514102
rect 255174 514046 255242 514102
rect 255298 514046 255366 514102
rect 255422 514046 255518 514102
rect 254898 513978 255518 514046
rect 254898 513922 254994 513978
rect 255050 513922 255118 513978
rect 255174 513922 255242 513978
rect 255298 513922 255366 513978
rect 255422 513922 255518 513978
rect 254898 496350 255518 513922
rect 254898 496294 254994 496350
rect 255050 496294 255118 496350
rect 255174 496294 255242 496350
rect 255298 496294 255366 496350
rect 255422 496294 255518 496350
rect 254898 496226 255518 496294
rect 254898 496170 254994 496226
rect 255050 496170 255118 496226
rect 255174 496170 255242 496226
rect 255298 496170 255366 496226
rect 255422 496170 255518 496226
rect 254898 496102 255518 496170
rect 254898 496046 254994 496102
rect 255050 496046 255118 496102
rect 255174 496046 255242 496102
rect 255298 496046 255366 496102
rect 255422 496046 255518 496102
rect 254898 495978 255518 496046
rect 254898 495922 254994 495978
rect 255050 495922 255118 495978
rect 255174 495922 255242 495978
rect 255298 495922 255366 495978
rect 255422 495922 255518 495978
rect 254898 478350 255518 495922
rect 254898 478294 254994 478350
rect 255050 478294 255118 478350
rect 255174 478294 255242 478350
rect 255298 478294 255366 478350
rect 255422 478294 255518 478350
rect 254898 478226 255518 478294
rect 254898 478170 254994 478226
rect 255050 478170 255118 478226
rect 255174 478170 255242 478226
rect 255298 478170 255366 478226
rect 255422 478170 255518 478226
rect 254898 478102 255518 478170
rect 254898 478046 254994 478102
rect 255050 478046 255118 478102
rect 255174 478046 255242 478102
rect 255298 478046 255366 478102
rect 255422 478046 255518 478102
rect 254898 477978 255518 478046
rect 254898 477922 254994 477978
rect 255050 477922 255118 477978
rect 255174 477922 255242 477978
rect 255298 477922 255366 477978
rect 255422 477922 255518 477978
rect 251178 472294 251274 472350
rect 251330 472294 251398 472350
rect 251454 472294 251522 472350
rect 251578 472294 251646 472350
rect 251702 472294 251798 472350
rect 251178 472226 251798 472294
rect 251178 472170 251274 472226
rect 251330 472170 251398 472226
rect 251454 472170 251522 472226
rect 251578 472170 251646 472226
rect 251702 472170 251798 472226
rect 251178 472102 251798 472170
rect 251178 472046 251274 472102
rect 251330 472046 251398 472102
rect 251454 472046 251522 472102
rect 251578 472046 251646 472102
rect 251702 472046 251798 472102
rect 251178 471978 251798 472046
rect 251178 471922 251274 471978
rect 251330 471922 251398 471978
rect 251454 471922 251522 471978
rect 251578 471922 251646 471978
rect 251702 471922 251798 471978
rect 249564 466138 249620 466148
rect 249564 462196 249620 466082
rect 249564 462130 249620 462140
rect 224178 460294 224274 460350
rect 224330 460294 224398 460350
rect 224454 460294 224522 460350
rect 224578 460294 224646 460350
rect 224702 460294 224798 460350
rect 224178 460226 224798 460294
rect 224178 460170 224274 460226
rect 224330 460170 224398 460226
rect 224454 460170 224522 460226
rect 224578 460170 224646 460226
rect 224702 460170 224798 460226
rect 224178 460102 224798 460170
rect 224178 460046 224274 460102
rect 224330 460046 224398 460102
rect 224454 460046 224522 460102
rect 224578 460046 224646 460102
rect 224702 460046 224798 460102
rect 224178 459978 224798 460046
rect 224178 459922 224274 459978
rect 224330 459922 224398 459978
rect 224454 459922 224522 459978
rect 224578 459922 224646 459978
rect 224702 459922 224798 459978
rect 224178 442350 224798 459922
rect 225808 460350 226128 460384
rect 225808 460294 225878 460350
rect 225934 460294 226002 460350
rect 226058 460294 226128 460350
rect 225808 460226 226128 460294
rect 225808 460170 225878 460226
rect 225934 460170 226002 460226
rect 226058 460170 226128 460226
rect 225808 460102 226128 460170
rect 225808 460046 225878 460102
rect 225934 460046 226002 460102
rect 226058 460046 226128 460102
rect 225808 459978 226128 460046
rect 225808 459922 225878 459978
rect 225934 459922 226002 459978
rect 226058 459922 226128 459978
rect 225808 459888 226128 459922
rect 230860 458164 230916 458174
rect 230860 456932 230916 458108
rect 230860 456866 230916 456876
rect 251178 454350 251798 471922
rect 251178 454294 251274 454350
rect 251330 454294 251398 454350
rect 251454 454294 251522 454350
rect 251578 454294 251646 454350
rect 251702 454294 251798 454350
rect 251178 454226 251798 454294
rect 251178 454170 251274 454226
rect 251330 454170 251398 454226
rect 251454 454170 251522 454226
rect 251578 454170 251646 454226
rect 251702 454170 251798 454226
rect 251178 454102 251798 454170
rect 251178 454046 251274 454102
rect 251330 454046 251398 454102
rect 251454 454046 251522 454102
rect 251578 454046 251646 454102
rect 251702 454046 251798 454102
rect 251178 453978 251798 454046
rect 251178 453922 251274 453978
rect 251330 453922 251398 453978
rect 251454 453922 251522 453978
rect 251578 453922 251646 453978
rect 251702 453922 251798 453978
rect 224178 442294 224274 442350
rect 224330 442294 224398 442350
rect 224454 442294 224522 442350
rect 224578 442294 224646 442350
rect 224702 442294 224798 442350
rect 224178 442226 224798 442294
rect 224178 442170 224274 442226
rect 224330 442170 224398 442226
rect 224454 442170 224522 442226
rect 224578 442170 224646 442226
rect 224702 442170 224798 442226
rect 224178 442102 224798 442170
rect 224178 442046 224274 442102
rect 224330 442046 224398 442102
rect 224454 442046 224522 442102
rect 224578 442046 224646 442102
rect 224702 442046 224798 442102
rect 224178 441978 224798 442046
rect 224178 441922 224274 441978
rect 224330 441922 224398 441978
rect 224454 441922 224522 441978
rect 224578 441922 224646 441978
rect 224702 441922 224798 441978
rect 222796 426468 222852 426478
rect 222796 426132 222852 426412
rect 222796 426066 222852 426076
rect 220458 418294 220554 418350
rect 220610 418294 220678 418350
rect 220734 418294 220802 418350
rect 220858 418294 220926 418350
rect 220982 418294 221078 418350
rect 220458 418226 221078 418294
rect 220458 418170 220554 418226
rect 220610 418170 220678 418226
rect 220734 418170 220802 418226
rect 220858 418170 220926 418226
rect 220982 418170 221078 418226
rect 220458 418102 221078 418170
rect 220458 418046 220554 418102
rect 220610 418046 220678 418102
rect 220734 418046 220802 418102
rect 220858 418046 220926 418102
rect 220982 418046 221078 418102
rect 220458 417978 221078 418046
rect 220458 417922 220554 417978
rect 220610 417922 220678 417978
rect 220734 417922 220802 417978
rect 220858 417922 220926 417978
rect 220982 417922 221078 417978
rect 206668 415044 206724 415056
rect 206668 414952 206724 414962
rect 201628 412498 201684 412508
rect 201628 412132 201684 412442
rect 201628 412066 201684 412076
rect 204764 411778 204820 411788
rect 203196 409444 203252 409454
rect 203196 383796 203252 409388
rect 204764 402052 204820 411722
rect 206108 408772 206164 408782
rect 204764 401986 204820 401996
rect 204876 408100 204932 408110
rect 203196 383730 203252 383740
rect 204876 380436 204932 408044
rect 204988 407098 205044 407108
rect 204988 405412 205044 407042
rect 204988 405346 205044 405356
rect 204988 404218 205044 404228
rect 204988 402958 205044 404162
rect 204988 402892 205044 402902
rect 204876 380370 204932 380380
rect 205772 395668 205828 395678
rect 205772 371476 205828 395612
rect 206108 381556 206164 408716
rect 210448 400350 210768 400384
rect 210448 400294 210518 400350
rect 210574 400294 210642 400350
rect 210698 400294 210768 400350
rect 210448 400226 210768 400294
rect 210448 400170 210518 400226
rect 210574 400170 210642 400226
rect 210698 400170 210768 400226
rect 210448 400102 210768 400170
rect 210448 400046 210518 400102
rect 210574 400046 210642 400102
rect 210698 400046 210768 400102
rect 210448 399978 210768 400046
rect 210448 399922 210518 399978
rect 210574 399922 210642 399978
rect 210698 399922 210768 399978
rect 210448 399888 210768 399922
rect 220458 400350 221078 417922
rect 220458 400294 220554 400350
rect 220610 400294 220678 400350
rect 220734 400294 220802 400350
rect 220858 400294 220926 400350
rect 220982 400294 221078 400350
rect 220458 400226 221078 400294
rect 220458 400170 220554 400226
rect 220610 400170 220678 400226
rect 220734 400170 220802 400226
rect 220858 400170 220926 400226
rect 220982 400170 221078 400226
rect 220458 400102 221078 400170
rect 220458 400046 220554 400102
rect 220610 400046 220678 400102
rect 220734 400046 220802 400102
rect 220858 400046 220926 400102
rect 220982 400046 221078 400102
rect 220458 399978 221078 400046
rect 220458 399922 220554 399978
rect 220610 399922 220678 399978
rect 220734 399922 220802 399978
rect 220858 399922 220926 399978
rect 220982 399922 221078 399978
rect 206108 381490 206164 381500
rect 220458 382350 221078 399922
rect 220458 382294 220554 382350
rect 220610 382294 220678 382350
rect 220734 382294 220802 382350
rect 220858 382294 220926 382350
rect 220982 382294 221078 382350
rect 220458 382226 221078 382294
rect 220458 382170 220554 382226
rect 220610 382170 220678 382226
rect 220734 382170 220802 382226
rect 220858 382170 220926 382226
rect 220982 382170 221078 382226
rect 220458 382102 221078 382170
rect 220458 382046 220554 382102
rect 220610 382046 220678 382102
rect 220734 382046 220802 382102
rect 220858 382046 220926 382102
rect 220982 382046 221078 382102
rect 220458 381978 221078 382046
rect 220458 381922 220554 381978
rect 220610 381922 220678 381978
rect 220734 381922 220802 381978
rect 220858 381922 220926 381978
rect 220982 381922 221078 381978
rect 205772 371410 205828 371420
rect 220458 364350 221078 381922
rect 220458 364294 220554 364350
rect 220610 364294 220678 364350
rect 220734 364294 220802 364350
rect 220858 364294 220926 364350
rect 220982 364294 221078 364350
rect 220458 364226 221078 364294
rect 220458 364170 220554 364226
rect 220610 364170 220678 364226
rect 220734 364170 220802 364226
rect 220858 364170 220926 364226
rect 220982 364170 221078 364226
rect 220458 364102 221078 364170
rect 220458 364046 220554 364102
rect 220610 364046 220678 364102
rect 220734 364046 220802 364102
rect 220858 364046 220926 364102
rect 220982 364046 221078 364102
rect 220458 363978 221078 364046
rect 220458 363922 220554 363978
rect 220610 363922 220678 363978
rect 220734 363922 220802 363978
rect 220858 363922 220926 363978
rect 220982 363922 221078 363978
rect 205660 356916 205716 356926
rect 204764 354116 204820 354126
rect 202972 352660 203028 352670
rect 202860 351092 202916 351102
rect 201292 341218 201348 341228
rect 201292 341012 201348 341162
rect 201292 340946 201348 340956
rect 200956 339668 201012 339678
rect 200956 312676 201012 339612
rect 202860 329588 202916 351036
rect 202972 333620 203028 352604
rect 202972 333554 203028 333564
rect 203084 348598 203140 348608
rect 203084 330932 203140 348542
rect 203084 330866 203140 330876
rect 204092 338548 204148 338558
rect 202860 329522 202916 329532
rect 204092 316036 204148 338492
rect 204764 332948 204820 354060
rect 205660 351092 205716 356860
rect 206668 355796 206724 355806
rect 205660 351026 205716 351036
rect 206220 354228 206276 354238
rect 205996 349498 206052 349508
rect 204764 332882 204820 332892
rect 204876 336308 204932 336318
rect 204876 324118 204932 336252
rect 204876 324052 204932 324062
rect 205772 332276 205828 332286
rect 204988 318388 205044 318398
rect 204988 317044 205044 318332
rect 204988 316978 205044 316988
rect 204092 315970 204148 315980
rect 205772 313684 205828 332220
rect 205996 330708 206052 349442
rect 205996 330642 206052 330652
rect 206108 338324 206164 338334
rect 206108 325558 206164 338268
rect 206220 334292 206276 354172
rect 206668 352660 206724 355740
rect 206668 352594 206724 352604
rect 210448 346350 210768 346384
rect 210448 346294 210518 346350
rect 210574 346294 210642 346350
rect 210698 346294 210768 346350
rect 210448 346226 210768 346294
rect 210448 346170 210518 346226
rect 210574 346170 210642 346226
rect 210698 346170 210768 346226
rect 210448 346102 210768 346170
rect 210448 346046 210518 346102
rect 210574 346046 210642 346102
rect 210698 346046 210768 346102
rect 210448 345978 210768 346046
rect 210448 345922 210518 345978
rect 210574 345922 210642 345978
rect 210698 345922 210768 345978
rect 210448 345888 210768 345922
rect 220458 346350 221078 363922
rect 220458 346294 220554 346350
rect 220610 346294 220678 346350
rect 220734 346294 220802 346350
rect 220858 346294 220926 346350
rect 220982 346294 221078 346350
rect 220458 346226 221078 346294
rect 220458 346170 220554 346226
rect 220610 346170 220678 346226
rect 220734 346170 220802 346226
rect 220858 346170 220926 346226
rect 220982 346170 221078 346226
rect 220458 346102 221078 346170
rect 220458 346046 220554 346102
rect 220610 346046 220678 346102
rect 220734 346046 220802 346102
rect 220858 346046 220926 346102
rect 220982 346046 221078 346102
rect 220458 345978 221078 346046
rect 220458 345922 220554 345978
rect 220610 345922 220678 345978
rect 220734 345922 220802 345978
rect 220858 345922 220926 345978
rect 220982 345922 221078 345978
rect 206220 334226 206276 334236
rect 210448 328350 210768 328384
rect 210448 328294 210518 328350
rect 210574 328294 210642 328350
rect 210698 328294 210768 328350
rect 210448 328226 210768 328294
rect 210448 328170 210518 328226
rect 210574 328170 210642 328226
rect 210698 328170 210768 328226
rect 210448 328102 210768 328170
rect 210448 328046 210518 328102
rect 210574 328046 210642 328102
rect 210698 328046 210768 328102
rect 210448 327978 210768 328046
rect 210448 327922 210518 327978
rect 210574 327922 210642 327978
rect 210698 327922 210768 327978
rect 210448 327888 210768 327922
rect 220458 328350 221078 345922
rect 220458 328294 220554 328350
rect 220610 328294 220678 328350
rect 220734 328294 220802 328350
rect 220858 328294 220926 328350
rect 220982 328294 221078 328350
rect 220458 328226 221078 328294
rect 220458 328170 220554 328226
rect 220610 328170 220678 328226
rect 220734 328170 220802 328226
rect 220858 328170 220926 328226
rect 220982 328170 221078 328226
rect 220458 328102 221078 328170
rect 220458 328046 220554 328102
rect 220610 328046 220678 328102
rect 220734 328046 220802 328102
rect 220858 328046 220926 328102
rect 220982 328046 221078 328102
rect 220458 327978 221078 328046
rect 220458 327922 220554 327978
rect 220610 327922 220678 327978
rect 220734 327922 220802 327978
rect 220858 327922 220926 327978
rect 220982 327922 221078 327978
rect 206108 325492 206164 325502
rect 205772 313618 205828 313628
rect 200956 312610 201012 312620
rect 220458 310350 221078 327922
rect 220458 310294 220554 310350
rect 220610 310294 220678 310350
rect 220734 310294 220802 310350
rect 220858 310294 220926 310350
rect 220982 310294 221078 310350
rect 220458 310226 221078 310294
rect 220458 310170 220554 310226
rect 220610 310170 220678 310226
rect 220734 310170 220802 310226
rect 220858 310170 220926 310226
rect 220982 310170 221078 310226
rect 220458 310102 221078 310170
rect 220458 310046 220554 310102
rect 220610 310046 220678 310102
rect 220734 310046 220802 310102
rect 220858 310046 220926 310102
rect 220982 310046 221078 310102
rect 220458 309978 221078 310046
rect 220458 309922 220554 309978
rect 220610 309922 220678 309978
rect 220734 309922 220802 309978
rect 220858 309922 220926 309978
rect 220982 309922 221078 309978
rect 202972 295876 203028 295886
rect 201628 271378 201684 271388
rect 201628 271124 201684 271322
rect 201628 271058 201684 271068
rect 202972 264404 203028 295820
rect 203084 294756 203140 294766
rect 203084 267092 203140 294700
rect 204764 293636 204820 293646
rect 203084 267026 203140 267036
rect 204092 283556 204148 283566
rect 202972 264338 203028 264348
rect 204092 263060 204148 283500
rect 204764 279188 204820 293580
rect 206108 293076 206164 293086
rect 204764 279122 204820 279132
rect 204876 291396 204932 291406
rect 204876 266420 204932 291340
rect 205772 284676 205828 284686
rect 205772 267764 205828 284620
rect 205772 267698 205828 267708
rect 204876 266354 204932 266364
rect 206108 265076 206164 293020
rect 220458 292350 221078 309922
rect 220458 292294 220554 292350
rect 220610 292294 220678 292350
rect 220734 292294 220802 292350
rect 220858 292294 220926 292350
rect 220982 292294 221078 292350
rect 220458 292226 221078 292294
rect 220458 292170 220554 292226
rect 220610 292170 220678 292226
rect 220734 292170 220802 292226
rect 220858 292170 220926 292226
rect 220982 292170 221078 292226
rect 220458 292102 221078 292170
rect 220458 292046 220554 292102
rect 220610 292046 220678 292102
rect 220734 292046 220802 292102
rect 220858 292046 220926 292102
rect 220982 292046 221078 292102
rect 220458 291978 221078 292046
rect 220458 291922 220554 291978
rect 220610 291922 220678 291978
rect 220734 291922 220802 291978
rect 220858 291922 220926 291978
rect 220982 291922 221078 291978
rect 210448 274350 210768 274384
rect 210448 274294 210518 274350
rect 210574 274294 210642 274350
rect 210698 274294 210768 274350
rect 210448 274226 210768 274294
rect 210448 274170 210518 274226
rect 210574 274170 210642 274226
rect 210698 274170 210768 274226
rect 210448 274102 210768 274170
rect 210448 274046 210518 274102
rect 210574 274046 210642 274102
rect 210698 274046 210768 274102
rect 210448 273978 210768 274046
rect 210448 273922 210518 273978
rect 210574 273922 210642 273978
rect 210698 273922 210768 273978
rect 210448 273888 210768 273922
rect 220458 274350 221078 291922
rect 220458 274294 220554 274350
rect 220610 274294 220678 274350
rect 220734 274294 220802 274350
rect 220858 274294 220926 274350
rect 220982 274294 221078 274350
rect 220458 274226 221078 274294
rect 220458 274170 220554 274226
rect 220610 274170 220678 274226
rect 220734 274170 220802 274226
rect 220858 274170 220926 274226
rect 220982 274170 221078 274226
rect 220458 274102 221078 274170
rect 220458 274046 220554 274102
rect 220610 274046 220678 274102
rect 220734 274046 220802 274102
rect 220858 274046 220926 274102
rect 220982 274046 221078 274102
rect 220458 273978 221078 274046
rect 220458 273922 220554 273978
rect 220610 273922 220678 273978
rect 220734 273922 220802 273978
rect 220858 273922 220926 273978
rect 220982 273922 221078 273978
rect 206444 267652 206500 267662
rect 206444 267238 206500 267596
rect 206444 267172 206500 267182
rect 206332 266518 206388 266528
rect 206332 266196 206388 266462
rect 206332 266130 206388 266140
rect 206108 265010 206164 265020
rect 204092 262994 204148 263004
rect 206444 261658 206500 261668
rect 206444 261538 206500 261548
rect 210448 256350 210768 256384
rect 210448 256294 210518 256350
rect 210574 256294 210642 256350
rect 210698 256294 210768 256350
rect 210448 256226 210768 256294
rect 210448 256170 210518 256226
rect 210574 256170 210642 256226
rect 210698 256170 210768 256226
rect 210448 256102 210768 256170
rect 210448 256046 210518 256102
rect 210574 256046 210642 256102
rect 210698 256046 210768 256102
rect 210448 255978 210768 256046
rect 210448 255922 210518 255978
rect 210574 255922 210642 255978
rect 210698 255922 210768 255978
rect 210448 255888 210768 255922
rect 220458 256350 221078 273922
rect 220458 256294 220554 256350
rect 220610 256294 220678 256350
rect 220734 256294 220802 256350
rect 220858 256294 220926 256350
rect 220982 256294 221078 256350
rect 220458 256226 221078 256294
rect 220458 256170 220554 256226
rect 220610 256170 220678 256226
rect 220734 256170 220802 256226
rect 220858 256170 220926 256226
rect 220982 256170 221078 256226
rect 220458 256102 221078 256170
rect 220458 256046 220554 256102
rect 220610 256046 220678 256102
rect 220734 256046 220802 256102
rect 220858 256046 220926 256102
rect 220982 256046 221078 256102
rect 220458 255978 221078 256046
rect 220458 255922 220554 255978
rect 220610 255922 220678 255978
rect 220734 255922 220802 255978
rect 220858 255922 220926 255978
rect 220982 255922 221078 255978
rect 220458 238350 221078 255922
rect 220458 238294 220554 238350
rect 220610 238294 220678 238350
rect 220734 238294 220802 238350
rect 220858 238294 220926 238350
rect 220982 238294 221078 238350
rect 220458 238226 221078 238294
rect 220458 238170 220554 238226
rect 220610 238170 220678 238226
rect 220734 238170 220802 238226
rect 220858 238170 220926 238226
rect 220982 238170 221078 238226
rect 220458 238102 221078 238170
rect 220458 238046 220554 238102
rect 220610 238046 220678 238102
rect 220734 238046 220802 238102
rect 220858 238046 220926 238102
rect 220982 238046 221078 238102
rect 220458 237978 221078 238046
rect 220458 237922 220554 237978
rect 220610 237922 220678 237978
rect 220734 237922 220802 237978
rect 220858 237922 220926 237978
rect 220982 237922 221078 237978
rect 203196 236516 203252 236526
rect 203084 234612 203140 234622
rect 202972 205858 203028 205868
rect 201628 199892 201684 199902
rect 201628 199018 201684 199836
rect 201628 198952 201684 198962
rect 202972 195188 203028 205802
rect 202972 195122 203028 195132
rect 203084 187796 203140 234556
rect 203084 187730 203140 187740
rect 203196 187124 203252 236460
rect 204876 236068 204932 236078
rect 204876 189140 204932 236012
rect 220458 220350 221078 237922
rect 220458 220294 220554 220350
rect 220610 220294 220678 220350
rect 220734 220294 220802 220350
rect 220858 220294 220926 220350
rect 220982 220294 221078 220350
rect 220458 220226 221078 220294
rect 220458 220170 220554 220226
rect 220610 220170 220678 220226
rect 220734 220170 220802 220226
rect 220858 220170 220926 220226
rect 220982 220170 221078 220226
rect 220458 220102 221078 220170
rect 220458 220046 220554 220102
rect 220610 220046 220678 220102
rect 220734 220046 220802 220102
rect 220858 220046 220926 220102
rect 220982 220046 221078 220102
rect 220458 219978 221078 220046
rect 220458 219922 220554 219978
rect 220610 219922 220678 219978
rect 220734 219922 220802 219978
rect 220858 219922 220926 219978
rect 220982 219922 221078 219978
rect 206668 214116 206724 214126
rect 206668 211092 206724 214060
rect 206668 211026 206724 211036
rect 210448 202350 210768 202384
rect 210448 202294 210518 202350
rect 210574 202294 210642 202350
rect 210698 202294 210768 202350
rect 210448 202226 210768 202294
rect 210448 202170 210518 202226
rect 210574 202170 210642 202226
rect 210698 202170 210768 202226
rect 210448 202102 210768 202170
rect 210448 202046 210518 202102
rect 210574 202046 210642 202102
rect 210698 202046 210768 202102
rect 210448 201978 210768 202046
rect 210448 201922 210518 201978
rect 210574 201922 210642 201978
rect 210698 201922 210768 201978
rect 210448 201888 210768 201922
rect 220458 202350 221078 219922
rect 220458 202294 220554 202350
rect 220610 202294 220678 202350
rect 220734 202294 220802 202350
rect 220858 202294 220926 202350
rect 220982 202294 221078 202350
rect 220458 202226 221078 202294
rect 220458 202170 220554 202226
rect 220610 202170 220678 202226
rect 220734 202170 220802 202226
rect 220858 202170 220926 202226
rect 220982 202170 221078 202226
rect 220458 202102 221078 202170
rect 220458 202046 220554 202102
rect 220610 202046 220678 202102
rect 220734 202046 220802 202102
rect 220858 202046 220926 202102
rect 220982 202046 221078 202102
rect 220458 201978 221078 202046
rect 220458 201922 220554 201978
rect 220610 201922 220678 201978
rect 220734 201922 220802 201978
rect 220858 201922 220926 201978
rect 220982 201922 221078 201978
rect 205660 198298 205716 198308
rect 204988 195058 205044 195068
rect 204988 192388 205044 195002
rect 204988 192322 205044 192332
rect 205660 191828 205716 198242
rect 205660 191762 205716 191772
rect 204876 189074 204932 189084
rect 203196 187058 203252 187068
rect 210448 184350 210768 184384
rect 210448 184294 210518 184350
rect 210574 184294 210642 184350
rect 210698 184294 210768 184350
rect 210448 184226 210768 184294
rect 210448 184170 210518 184226
rect 210574 184170 210642 184226
rect 210698 184170 210768 184226
rect 210448 184102 210768 184170
rect 210448 184046 210518 184102
rect 210574 184046 210642 184102
rect 210698 184046 210768 184102
rect 210448 183978 210768 184046
rect 210448 183922 210518 183978
rect 210574 183922 210642 183978
rect 210698 183922 210768 183978
rect 210448 183888 210768 183922
rect 220458 184350 221078 201922
rect 220458 184294 220554 184350
rect 220610 184294 220678 184350
rect 220734 184294 220802 184350
rect 220858 184294 220926 184350
rect 220982 184294 221078 184350
rect 220458 184226 221078 184294
rect 220458 184170 220554 184226
rect 220610 184170 220678 184226
rect 220734 184170 220802 184226
rect 220858 184170 220926 184226
rect 220982 184170 221078 184226
rect 220458 184102 221078 184170
rect 220458 184046 220554 184102
rect 220610 184046 220678 184102
rect 220734 184046 220802 184102
rect 220858 184046 220926 184102
rect 220982 184046 221078 184102
rect 220458 183978 221078 184046
rect 220458 183922 220554 183978
rect 220610 183922 220678 183978
rect 220734 183922 220802 183978
rect 220858 183922 220926 183978
rect 220982 183922 221078 183978
rect 206108 174020 206164 174030
rect 204876 172228 204932 172238
rect 203084 147476 203140 147486
rect 201628 128458 201684 128468
rect 201628 127988 201684 128402
rect 201628 127922 201684 127932
rect 203084 123956 203140 147420
rect 203084 123890 203140 123900
rect 203196 145236 203252 145246
rect 203196 119924 203252 145180
rect 203196 119858 203252 119868
rect 204092 144788 204148 144798
rect 204092 119252 204148 144732
rect 204876 125972 204932 172172
rect 204876 125906 204932 125916
rect 205772 140196 205828 140206
rect 205772 123284 205828 140140
rect 206108 125300 206164 173964
rect 220458 166350 221078 183922
rect 220458 166294 220554 166350
rect 220610 166294 220678 166350
rect 220734 166294 220802 166350
rect 220858 166294 220926 166350
rect 220982 166294 221078 166350
rect 220458 166226 221078 166294
rect 220458 166170 220554 166226
rect 220610 166170 220678 166226
rect 220734 166170 220802 166226
rect 220858 166170 220926 166226
rect 220982 166170 221078 166226
rect 220458 166102 221078 166170
rect 220458 166046 220554 166102
rect 220610 166046 220678 166102
rect 220734 166046 220802 166102
rect 220858 166046 220926 166102
rect 220982 166046 221078 166102
rect 220458 165978 221078 166046
rect 220458 165922 220554 165978
rect 220610 165922 220678 165978
rect 220734 165922 220802 165978
rect 220858 165922 220926 165978
rect 220982 165922 221078 165978
rect 220458 148350 221078 165922
rect 220458 148294 220554 148350
rect 220610 148294 220678 148350
rect 220734 148294 220802 148350
rect 220858 148294 220926 148350
rect 220982 148294 221078 148350
rect 220458 148226 221078 148294
rect 220458 148170 220554 148226
rect 220610 148170 220678 148226
rect 220734 148170 220802 148226
rect 220858 148170 220926 148226
rect 220982 148170 221078 148226
rect 220458 148102 221078 148170
rect 220458 148046 220554 148102
rect 220610 148046 220678 148102
rect 220734 148046 220802 148102
rect 220858 148046 220926 148102
rect 220982 148046 221078 148102
rect 220458 147978 221078 148046
rect 220458 147922 220554 147978
rect 220610 147922 220678 147978
rect 220734 147922 220802 147978
rect 220858 147922 220926 147978
rect 220982 147922 221078 147978
rect 206668 142996 206724 143006
rect 206668 138628 206724 142940
rect 206668 138562 206724 138572
rect 210448 130350 210768 130384
rect 210448 130294 210518 130350
rect 210574 130294 210642 130350
rect 210698 130294 210768 130350
rect 210448 130226 210768 130294
rect 210448 130170 210518 130226
rect 210574 130170 210642 130226
rect 210698 130170 210768 130226
rect 210448 130102 210768 130170
rect 210448 130046 210518 130102
rect 210574 130046 210642 130102
rect 210698 130046 210768 130102
rect 210448 129978 210768 130046
rect 210448 129922 210518 129978
rect 210574 129922 210642 129978
rect 210698 129922 210768 129978
rect 210448 129888 210768 129922
rect 220458 130350 221078 147922
rect 220458 130294 220554 130350
rect 220610 130294 220678 130350
rect 220734 130294 220802 130350
rect 220858 130294 220926 130350
rect 220982 130294 221078 130350
rect 220458 130226 221078 130294
rect 220458 130170 220554 130226
rect 220610 130170 220678 130226
rect 220734 130170 220802 130226
rect 220858 130170 220926 130226
rect 220982 130170 221078 130226
rect 220458 130102 221078 130170
rect 220458 130046 220554 130102
rect 220610 130046 220678 130102
rect 220734 130046 220802 130102
rect 220858 130046 220926 130102
rect 220982 130046 221078 130102
rect 220458 129978 221078 130046
rect 220458 129922 220554 129978
rect 220610 129922 220678 129978
rect 220734 129922 220802 129978
rect 220858 129922 220926 129978
rect 220982 129922 221078 129978
rect 206108 125234 206164 125244
rect 205772 123218 205828 123228
rect 204092 119186 204148 119196
rect 210448 112350 210768 112384
rect 210448 112294 210518 112350
rect 210574 112294 210642 112350
rect 210698 112294 210768 112350
rect 210448 112226 210768 112294
rect 210448 112170 210518 112226
rect 210574 112170 210642 112226
rect 210698 112170 210768 112226
rect 210448 112102 210768 112170
rect 210448 112046 210518 112102
rect 210574 112046 210642 112102
rect 210698 112046 210768 112102
rect 210448 111978 210768 112046
rect 210448 111922 210518 111978
rect 210574 111922 210642 111978
rect 210698 111922 210768 111978
rect 210448 111888 210768 111922
rect 220458 112350 221078 129922
rect 220458 112294 220554 112350
rect 220610 112294 220678 112350
rect 220734 112294 220802 112350
rect 220858 112294 220926 112350
rect 220982 112294 221078 112350
rect 220458 112226 221078 112294
rect 220458 112170 220554 112226
rect 220610 112170 220678 112226
rect 220734 112170 220802 112226
rect 220858 112170 220926 112226
rect 220982 112170 221078 112226
rect 220458 112102 221078 112170
rect 220458 112046 220554 112102
rect 220610 112046 220678 112102
rect 220734 112046 220802 112102
rect 220858 112046 220926 112102
rect 220982 112046 221078 112102
rect 220458 111978 221078 112046
rect 220458 111922 220554 111978
rect 220610 111922 220678 111978
rect 220734 111922 220802 111978
rect 220858 111922 220926 111978
rect 220982 111922 221078 111978
rect 200956 98308 201012 98318
rect 200956 50148 201012 98252
rect 220458 94350 221078 111922
rect 220458 94294 220554 94350
rect 220610 94294 220678 94350
rect 220734 94294 220802 94350
rect 220858 94294 220926 94350
rect 220982 94294 221078 94350
rect 220458 94226 221078 94294
rect 220458 94170 220554 94226
rect 220610 94170 220678 94226
rect 220734 94170 220802 94226
rect 220858 94170 220926 94226
rect 220982 94170 221078 94226
rect 220458 94102 221078 94170
rect 220458 94046 220554 94102
rect 220610 94046 220678 94102
rect 220734 94046 220802 94102
rect 220858 94046 220926 94102
rect 220982 94046 221078 94102
rect 220458 93978 221078 94046
rect 220458 93922 220554 93978
rect 220610 93922 220678 93978
rect 220734 93922 220802 93978
rect 220858 93922 220926 93978
rect 220982 93922 221078 93978
rect 202860 90244 202916 90254
rect 202860 54180 202916 90188
rect 204876 88116 204932 88126
rect 203084 78372 203140 78382
rect 202860 54114 202916 54124
rect 202972 69972 203028 69982
rect 202972 52836 203028 69916
rect 203084 53508 203140 78316
rect 203196 73332 203252 73342
rect 203196 65604 203252 73276
rect 203196 65538 203252 65548
rect 203196 56868 203252 56878
rect 203196 56278 203252 56812
rect 203196 56212 203252 56222
rect 204876 56196 204932 88060
rect 204876 56130 204932 56140
rect 205772 86436 205828 86446
rect 203084 53442 203140 53452
rect 202972 52770 203028 52780
rect 200956 50082 201012 50092
rect 205772 46004 205828 86380
rect 220458 76350 221078 93922
rect 220458 76294 220554 76350
rect 220610 76294 220678 76350
rect 220734 76294 220802 76350
rect 220858 76294 220926 76350
rect 220982 76294 221078 76350
rect 220458 76226 221078 76294
rect 220458 76170 220554 76226
rect 220610 76170 220678 76226
rect 220734 76170 220802 76226
rect 220858 76170 220926 76226
rect 220982 76170 221078 76226
rect 220458 76102 221078 76170
rect 220458 76046 220554 76102
rect 220610 76046 220678 76102
rect 220734 76046 220802 76102
rect 220858 76046 220926 76102
rect 220982 76046 221078 76102
rect 220458 75978 221078 76046
rect 220458 75922 220554 75978
rect 220610 75922 220678 75978
rect 220734 75922 220802 75978
rect 220858 75922 220926 75978
rect 220982 75922 221078 75978
rect 210448 58350 210768 58384
rect 210448 58294 210518 58350
rect 210574 58294 210642 58350
rect 210698 58294 210768 58350
rect 210448 58226 210768 58294
rect 210448 58170 210518 58226
rect 210574 58170 210642 58226
rect 210698 58170 210768 58226
rect 210448 58102 210768 58170
rect 210448 58046 210518 58102
rect 210574 58046 210642 58102
rect 210698 58046 210768 58102
rect 210448 57978 210768 58046
rect 210448 57922 210518 57978
rect 210574 57922 210642 57978
rect 210698 57922 210768 57978
rect 210448 57888 210768 57922
rect 220458 58350 221078 75922
rect 220458 58294 220554 58350
rect 220610 58294 220678 58350
rect 220734 58294 220802 58350
rect 220858 58294 220926 58350
rect 220982 58294 221078 58350
rect 220458 58226 221078 58294
rect 220458 58170 220554 58226
rect 220610 58170 220678 58226
rect 220734 58170 220802 58226
rect 220858 58170 220926 58226
rect 220982 58170 221078 58226
rect 220458 58102 221078 58170
rect 220458 58046 220554 58102
rect 220610 58046 220678 58102
rect 220734 58046 220802 58102
rect 220858 58046 220926 58102
rect 220982 58046 221078 58102
rect 220458 57978 221078 58046
rect 220458 57922 220554 57978
rect 220610 57922 220678 57978
rect 220734 57922 220802 57978
rect 220858 57922 220926 57978
rect 220982 57922 221078 57978
rect 206108 56308 206164 56318
rect 206108 56098 206164 56252
rect 206108 56032 206164 56042
rect 205772 45938 205828 45948
rect 210448 40350 210768 40384
rect 210448 40294 210518 40350
rect 210574 40294 210642 40350
rect 210698 40294 210768 40350
rect 210448 40226 210768 40294
rect 210448 40170 210518 40226
rect 210574 40170 210642 40226
rect 210698 40170 210768 40226
rect 210448 40102 210768 40170
rect 210448 40046 210518 40102
rect 210574 40046 210642 40102
rect 210698 40046 210768 40102
rect 210448 39978 210768 40046
rect 210448 39922 210518 39978
rect 210574 39922 210642 39978
rect 210698 39922 210768 39978
rect 210448 39888 210768 39922
rect 220458 40350 221078 57922
rect 220458 40294 220554 40350
rect 220610 40294 220678 40350
rect 220734 40294 220802 40350
rect 220858 40294 220926 40350
rect 220982 40294 221078 40350
rect 220458 40226 221078 40294
rect 220458 40170 220554 40226
rect 220610 40170 220678 40226
rect 220734 40170 220802 40226
rect 220858 40170 220926 40226
rect 220982 40170 221078 40226
rect 220458 40102 221078 40170
rect 220458 40046 220554 40102
rect 220610 40046 220678 40102
rect 220734 40046 220802 40102
rect 220858 40046 220926 40102
rect 220982 40046 221078 40102
rect 220458 39978 221078 40046
rect 220458 39922 220554 39978
rect 220610 39922 220678 39978
rect 220734 39922 220802 39978
rect 220858 39922 220926 39978
rect 220982 39922 221078 39978
rect 200844 8530 200900 8540
rect 220458 22350 221078 39922
rect 220458 22294 220554 22350
rect 220610 22294 220678 22350
rect 220734 22294 220802 22350
rect 220858 22294 220926 22350
rect 220982 22294 221078 22350
rect 220458 22226 221078 22294
rect 220458 22170 220554 22226
rect 220610 22170 220678 22226
rect 220734 22170 220802 22226
rect 220858 22170 220926 22226
rect 220982 22170 221078 22226
rect 220458 22102 221078 22170
rect 220458 22046 220554 22102
rect 220610 22046 220678 22102
rect 220734 22046 220802 22102
rect 220858 22046 220926 22102
rect 220982 22046 221078 22102
rect 220458 21978 221078 22046
rect 220458 21922 220554 21978
rect 220610 21922 220678 21978
rect 220734 21922 220802 21978
rect 220858 21922 220926 21978
rect 220982 21922 221078 21978
rect 193458 -1176 193554 -1120
rect 193610 -1176 193678 -1120
rect 193734 -1176 193802 -1120
rect 193858 -1176 193926 -1120
rect 193982 -1176 194078 -1120
rect 193458 -1244 194078 -1176
rect 193458 -1300 193554 -1244
rect 193610 -1300 193678 -1244
rect 193734 -1300 193802 -1244
rect 193858 -1300 193926 -1244
rect 193982 -1300 194078 -1244
rect 193458 -1368 194078 -1300
rect 193458 -1424 193554 -1368
rect 193610 -1424 193678 -1368
rect 193734 -1424 193802 -1368
rect 193858 -1424 193926 -1368
rect 193982 -1424 194078 -1368
rect 193458 -1492 194078 -1424
rect 193458 -1548 193554 -1492
rect 193610 -1548 193678 -1492
rect 193734 -1548 193802 -1492
rect 193858 -1548 193926 -1492
rect 193982 -1548 194078 -1492
rect 193458 -1644 194078 -1548
rect 220458 4350 221078 21922
rect 220458 4294 220554 4350
rect 220610 4294 220678 4350
rect 220734 4294 220802 4350
rect 220858 4294 220926 4350
rect 220982 4294 221078 4350
rect 220458 4226 221078 4294
rect 220458 4170 220554 4226
rect 220610 4170 220678 4226
rect 220734 4170 220802 4226
rect 220858 4170 220926 4226
rect 220982 4170 221078 4226
rect 220458 4102 221078 4170
rect 220458 4046 220554 4102
rect 220610 4046 220678 4102
rect 220734 4046 220802 4102
rect 220858 4046 220926 4102
rect 220982 4046 221078 4102
rect 220458 3978 221078 4046
rect 220458 3922 220554 3978
rect 220610 3922 220678 3978
rect 220734 3922 220802 3978
rect 220858 3922 220926 3978
rect 220982 3922 221078 3978
rect 220458 -160 221078 3922
rect 220458 -216 220554 -160
rect 220610 -216 220678 -160
rect 220734 -216 220802 -160
rect 220858 -216 220926 -160
rect 220982 -216 221078 -160
rect 220458 -284 221078 -216
rect 220458 -340 220554 -284
rect 220610 -340 220678 -284
rect 220734 -340 220802 -284
rect 220858 -340 220926 -284
rect 220982 -340 221078 -284
rect 220458 -408 221078 -340
rect 220458 -464 220554 -408
rect 220610 -464 220678 -408
rect 220734 -464 220802 -408
rect 220858 -464 220926 -408
rect 220982 -464 221078 -408
rect 220458 -532 221078 -464
rect 220458 -588 220554 -532
rect 220610 -588 220678 -532
rect 220734 -588 220802 -532
rect 220858 -588 220926 -532
rect 220982 -588 221078 -532
rect 220458 -1644 221078 -588
rect 224178 424350 224798 441922
rect 247772 449428 247828 449438
rect 232204 426468 232260 426478
rect 232204 426020 232260 426412
rect 232204 425954 232260 425964
rect 224178 424294 224274 424350
rect 224330 424294 224398 424350
rect 224454 424294 224522 424350
rect 224578 424294 224646 424350
rect 224702 424294 224798 424350
rect 224178 424226 224798 424294
rect 224178 424170 224274 424226
rect 224330 424170 224398 424226
rect 224454 424170 224522 424226
rect 224578 424170 224646 424226
rect 224702 424170 224798 424226
rect 224178 424102 224798 424170
rect 224178 424046 224274 424102
rect 224330 424046 224398 424102
rect 224454 424046 224522 424102
rect 224578 424046 224646 424102
rect 224702 424046 224798 424102
rect 224178 423978 224798 424046
rect 224178 423922 224274 423978
rect 224330 423922 224398 423978
rect 224454 423922 224522 423978
rect 224578 423922 224646 423978
rect 224702 423922 224798 423978
rect 224178 406350 224798 423922
rect 247772 419636 247828 449372
rect 247884 438004 247940 438014
rect 247884 424116 247940 437948
rect 247884 424050 247940 424060
rect 251178 436350 251798 453922
rect 252812 477316 252868 477326
rect 252812 439796 252868 477260
rect 254898 460350 255518 477922
rect 256172 530068 256228 530078
rect 256172 477876 256228 530012
rect 256284 524916 256340 544460
rect 256284 524850 256340 524860
rect 256508 521780 256564 521790
rect 256172 477810 256228 477820
rect 256284 521668 256340 521678
rect 256284 475076 256340 521612
rect 256508 485156 256564 521724
rect 257852 500276 257908 548492
rect 259980 545188 260036 545198
rect 259532 530180 259588 530190
rect 257852 500210 257908 500220
rect 257964 514948 258020 514958
rect 257964 486276 258020 514892
rect 257964 486210 258020 486220
rect 256508 485090 256564 485100
rect 259532 479556 259588 530124
rect 259980 526596 260036 545132
rect 259980 526530 260036 526540
rect 261212 543844 261268 543854
rect 261212 499156 261268 543788
rect 261324 528836 261380 552524
rect 261324 528770 261380 528780
rect 262892 551236 262948 551246
rect 261548 528276 261604 528286
rect 261548 507556 261604 528220
rect 261548 507490 261604 507500
rect 262892 500164 262948 551180
rect 287808 550350 288128 550384
rect 287808 550294 287878 550350
rect 287934 550294 288002 550350
rect 288058 550294 288128 550350
rect 287808 550226 288128 550294
rect 287808 550170 287878 550226
rect 287934 550170 288002 550226
rect 288058 550170 288128 550226
rect 287808 550102 288128 550170
rect 287808 550046 287878 550102
rect 287934 550046 288002 550102
rect 288058 550046 288128 550102
rect 287808 549978 288128 550046
rect 287808 549922 287878 549978
rect 287934 549922 288002 549978
rect 288058 549922 288128 549978
rect 287808 549888 288128 549922
rect 318528 550350 318848 550384
rect 318528 550294 318598 550350
rect 318654 550294 318722 550350
rect 318778 550294 318848 550350
rect 318528 550226 318848 550294
rect 318528 550170 318598 550226
rect 318654 550170 318722 550226
rect 318778 550170 318848 550226
rect 318528 550102 318848 550170
rect 318528 550046 318598 550102
rect 318654 550046 318722 550102
rect 318778 550046 318848 550102
rect 318528 549978 318848 550046
rect 318528 549922 318598 549978
rect 318654 549922 318722 549978
rect 318778 549922 318848 549978
rect 318528 549888 318848 549922
rect 264572 547876 264628 547886
rect 263788 533458 263844 533468
rect 263788 531076 263844 533402
rect 263788 531010 263844 531020
rect 263900 533428 263956 533438
rect 263900 529396 263956 533372
rect 263900 529330 263956 529340
rect 263788 519988 263844 519998
rect 262892 500098 262948 500108
rect 263116 518308 263172 518318
rect 261212 499090 261268 499100
rect 259532 479490 259588 479500
rect 259644 482692 259700 482702
rect 256284 475010 256340 475020
rect 259532 476644 259588 476654
rect 254898 460294 254994 460350
rect 255050 460294 255118 460350
rect 255174 460294 255242 460350
rect 255298 460294 255366 460350
rect 255422 460294 255518 460350
rect 254898 460226 255518 460294
rect 254898 460170 254994 460226
rect 255050 460170 255118 460226
rect 255174 460170 255242 460226
rect 255298 460170 255366 460226
rect 255422 460170 255518 460226
rect 254898 460102 255518 460170
rect 254898 460046 254994 460102
rect 255050 460046 255118 460102
rect 255174 460046 255242 460102
rect 255298 460046 255366 460102
rect 255422 460046 255518 460102
rect 254898 459978 255518 460046
rect 254898 459922 254994 459978
rect 255050 459922 255118 459978
rect 255174 459922 255242 459978
rect 255298 459922 255366 459978
rect 255422 459922 255518 459978
rect 252812 439730 252868 439740
rect 253148 444500 253204 444510
rect 251178 436294 251274 436350
rect 251330 436294 251398 436350
rect 251454 436294 251522 436350
rect 251578 436294 251646 436350
rect 251702 436294 251798 436350
rect 251178 436226 251798 436294
rect 251178 436170 251274 436226
rect 251330 436170 251398 436226
rect 251454 436170 251522 436226
rect 251578 436170 251646 436226
rect 251702 436170 251798 436226
rect 251178 436102 251798 436170
rect 251178 436046 251274 436102
rect 251330 436046 251398 436102
rect 251454 436046 251522 436102
rect 251578 436046 251646 436102
rect 251702 436046 251798 436102
rect 251178 435978 251798 436046
rect 251178 435922 251274 435978
rect 251330 435922 251398 435978
rect 251454 435922 251522 435978
rect 251578 435922 251646 435978
rect 251702 435922 251798 435978
rect 247772 419570 247828 419580
rect 241168 418350 241488 418384
rect 241168 418294 241238 418350
rect 241294 418294 241362 418350
rect 241418 418294 241488 418350
rect 241168 418226 241488 418294
rect 241168 418170 241238 418226
rect 241294 418170 241362 418226
rect 241418 418170 241488 418226
rect 241168 418102 241488 418170
rect 241168 418046 241238 418102
rect 241294 418046 241362 418102
rect 241418 418046 241488 418102
rect 241168 417978 241488 418046
rect 241168 417922 241238 417978
rect 241294 417922 241362 417978
rect 241418 417922 241488 417978
rect 241168 417888 241488 417922
rect 251178 418350 251798 435922
rect 253148 429156 253204 444444
rect 253148 429090 253204 429100
rect 254898 442350 255518 459922
rect 254898 442294 254994 442350
rect 255050 442294 255118 442350
rect 255174 442294 255242 442350
rect 255298 442294 255366 442350
rect 255422 442294 255518 442350
rect 254898 442226 255518 442294
rect 254898 442170 254994 442226
rect 255050 442170 255118 442226
rect 255174 442170 255242 442226
rect 255298 442170 255366 442226
rect 255422 442170 255518 442226
rect 254898 442102 255518 442170
rect 254898 442046 254994 442102
rect 255050 442046 255118 442102
rect 255174 442046 255242 442102
rect 255298 442046 255366 442102
rect 255422 442046 255518 442102
rect 254898 441978 255518 442046
rect 254898 441922 254994 441978
rect 255050 441922 255118 441978
rect 255174 441922 255242 441978
rect 255298 441922 255366 441978
rect 255422 441922 255518 441978
rect 251178 418294 251274 418350
rect 251330 418294 251398 418350
rect 251454 418294 251522 418350
rect 251578 418294 251646 418350
rect 251702 418294 251798 418350
rect 251178 418226 251798 418294
rect 251178 418170 251274 418226
rect 251330 418170 251398 418226
rect 251454 418170 251522 418226
rect 251578 418170 251646 418226
rect 251702 418170 251798 418226
rect 251178 418102 251798 418170
rect 251178 418046 251274 418102
rect 251330 418046 251398 418102
rect 251454 418046 251522 418102
rect 251578 418046 251646 418102
rect 251702 418046 251798 418102
rect 251178 417978 251798 418046
rect 251178 417922 251274 417978
rect 251330 417922 251398 417978
rect 251454 417922 251522 417978
rect 251578 417922 251646 417978
rect 251702 417922 251798 417978
rect 249452 409078 249508 409088
rect 224178 406294 224274 406350
rect 224330 406294 224398 406350
rect 224454 406294 224522 406350
rect 224578 406294 224646 406350
rect 224702 406294 224798 406350
rect 224178 406226 224798 406294
rect 224178 406170 224274 406226
rect 224330 406170 224398 406226
rect 224454 406170 224522 406226
rect 224578 406170 224646 406226
rect 224702 406170 224798 406226
rect 224178 406102 224798 406170
rect 224178 406046 224274 406102
rect 224330 406046 224398 406102
rect 224454 406046 224522 406102
rect 224578 406046 224646 406102
rect 224702 406046 224798 406102
rect 224178 405978 224798 406046
rect 224178 405922 224274 405978
rect 224330 405922 224398 405978
rect 224454 405922 224522 405978
rect 224578 405922 224646 405978
rect 224702 405922 224798 405978
rect 224178 388350 224798 405922
rect 225808 406350 226128 406384
rect 225808 406294 225878 406350
rect 225934 406294 226002 406350
rect 226058 406294 226128 406350
rect 225808 406226 226128 406294
rect 225808 406170 225878 406226
rect 225934 406170 226002 406226
rect 226058 406170 226128 406226
rect 225808 406102 226128 406170
rect 225808 406046 225878 406102
rect 225934 406046 226002 406102
rect 226058 406046 226128 406102
rect 225808 405978 226128 406046
rect 225808 405922 225878 405978
rect 225934 405922 226002 405978
rect 226058 405922 226128 405978
rect 225808 405888 226128 405922
rect 241168 400350 241488 400384
rect 241168 400294 241238 400350
rect 241294 400294 241362 400350
rect 241418 400294 241488 400350
rect 241168 400226 241488 400294
rect 241168 400170 241238 400226
rect 241294 400170 241362 400226
rect 241418 400170 241488 400226
rect 241168 400102 241488 400170
rect 241168 400046 241238 400102
rect 241294 400046 241362 400102
rect 241418 400046 241488 400102
rect 241168 399978 241488 400046
rect 241168 399922 241238 399978
rect 241294 399922 241362 399978
rect 241418 399922 241488 399978
rect 241168 399888 241488 399922
rect 249452 396676 249508 409022
rect 249452 396610 249508 396620
rect 251178 400350 251798 417922
rect 254898 424350 255518 441922
rect 256508 474852 256564 474862
rect 256172 441140 256228 441150
rect 255612 432628 255668 432638
rect 255612 428596 255668 432572
rect 255612 428530 255668 428540
rect 254898 424294 254994 424350
rect 255050 424294 255118 424350
rect 255174 424294 255242 424350
rect 255298 424294 255366 424350
rect 255422 424294 255518 424350
rect 254898 424226 255518 424294
rect 254898 424170 254994 424226
rect 255050 424170 255118 424226
rect 255174 424170 255242 424226
rect 255298 424170 255366 424226
rect 255422 424170 255518 424226
rect 254898 424102 255518 424170
rect 254898 424046 254994 424102
rect 255050 424046 255118 424102
rect 255174 424046 255242 424102
rect 255298 424046 255366 424102
rect 255422 424046 255518 424102
rect 254898 423978 255518 424046
rect 254898 423922 254994 423978
rect 255050 423922 255118 423978
rect 255174 423922 255242 423978
rect 255298 423922 255366 423978
rect 255422 423922 255518 423978
rect 252812 409978 252868 409988
rect 252812 403508 252868 409922
rect 254898 406350 255518 423922
rect 256172 419076 256228 441084
rect 256508 440916 256564 474796
rect 256508 440850 256564 440860
rect 257852 473284 257908 473294
rect 257852 439236 257908 473228
rect 259532 466116 259588 476588
rect 259532 466050 259588 466060
rect 257852 439170 257908 439180
rect 258188 452900 258244 452910
rect 258188 425236 258244 452844
rect 258188 425170 258244 425180
rect 259532 441028 259588 441038
rect 259532 420756 259588 440972
rect 259644 438116 259700 482636
rect 262892 482020 262948 482030
rect 261324 480676 261380 480686
rect 261212 475972 261268 475982
rect 261212 441924 261268 475916
rect 261324 467796 261380 480620
rect 262108 473956 262164 473966
rect 262108 470036 262164 473900
rect 262108 469970 262164 469980
rect 261324 467730 261380 467740
rect 261212 441858 261268 441868
rect 261324 446068 261380 446078
rect 259644 438050 259700 438060
rect 259532 420690 259588 420700
rect 261212 437668 261268 437678
rect 261212 420196 261268 437612
rect 261324 423556 261380 446012
rect 262892 437556 262948 481964
rect 263116 481796 263172 518252
rect 263788 514276 263844 519932
rect 263788 514210 263844 514220
rect 263788 509908 263844 509918
rect 263788 508116 263844 509852
rect 263788 508050 263844 508060
rect 263900 500164 263956 500174
rect 263900 498036 263956 500108
rect 264572 499716 264628 547820
rect 272448 544350 272768 544384
rect 272448 544294 272518 544350
rect 272574 544294 272642 544350
rect 272698 544294 272768 544350
rect 272448 544226 272768 544294
rect 272448 544170 272518 544226
rect 272574 544170 272642 544226
rect 272698 544170 272768 544226
rect 272448 544102 272768 544170
rect 272448 544046 272518 544102
rect 272574 544046 272642 544102
rect 272698 544046 272768 544102
rect 272448 543978 272768 544046
rect 272448 543922 272518 543978
rect 272574 543922 272642 543978
rect 272698 543922 272768 543978
rect 272448 543888 272768 543922
rect 303168 544350 303488 544384
rect 303168 544294 303238 544350
rect 303294 544294 303362 544350
rect 303418 544294 303488 544350
rect 303168 544226 303488 544294
rect 303168 544170 303238 544226
rect 303294 544170 303362 544226
rect 303418 544170 303488 544226
rect 303168 544102 303488 544170
rect 303168 544046 303238 544102
rect 303294 544046 303362 544102
rect 303418 544046 303488 544102
rect 303168 543978 303488 544046
rect 303168 543922 303238 543978
rect 303294 543922 303362 543978
rect 303418 543922 303488 543978
rect 303168 543888 303488 543922
rect 287808 532350 288128 532384
rect 287808 532294 287878 532350
rect 287934 532294 288002 532350
rect 288058 532294 288128 532350
rect 287808 532226 288128 532294
rect 287808 532170 287878 532226
rect 287934 532170 288002 532226
rect 288058 532170 288128 532226
rect 287808 532102 288128 532170
rect 287808 532046 287878 532102
rect 287934 532046 288002 532102
rect 288058 532046 288128 532102
rect 287808 531978 288128 532046
rect 287808 531922 287878 531978
rect 287934 531922 288002 531978
rect 288058 531922 288128 531978
rect 287808 531888 288128 531922
rect 318528 532350 318848 532384
rect 318528 532294 318598 532350
rect 318654 532294 318722 532350
rect 318778 532294 318848 532350
rect 318528 532226 318848 532294
rect 318528 532170 318598 532226
rect 318654 532170 318722 532226
rect 318778 532170 318848 532226
rect 318528 532102 318848 532170
rect 318528 532046 318598 532102
rect 318654 532046 318722 532102
rect 318778 532046 318848 532102
rect 318528 531978 318848 532046
rect 318528 531922 318598 531978
rect 318654 531922 318722 531978
rect 318778 531922 318848 531978
rect 318528 531888 318848 531922
rect 332668 528388 332724 528398
rect 332668 527828 332724 528332
rect 332668 527762 332724 527772
rect 272448 526350 272768 526384
rect 272448 526294 272518 526350
rect 272574 526294 272642 526350
rect 272698 526294 272768 526350
rect 272448 526226 272768 526294
rect 272448 526170 272518 526226
rect 272574 526170 272642 526226
rect 272698 526170 272768 526226
rect 272448 526102 272768 526170
rect 272448 526046 272518 526102
rect 272574 526046 272642 526102
rect 272698 526046 272768 526102
rect 272448 525978 272768 526046
rect 272448 525922 272518 525978
rect 272574 525922 272642 525978
rect 272698 525922 272768 525978
rect 272448 525888 272768 525922
rect 303168 526350 303488 526384
rect 303168 526294 303238 526350
rect 303294 526294 303362 526350
rect 303418 526294 303488 526350
rect 303168 526226 303488 526294
rect 303168 526170 303238 526226
rect 303294 526170 303362 526226
rect 303418 526170 303488 526226
rect 303168 526102 303488 526170
rect 303168 526046 303238 526102
rect 303294 526046 303362 526102
rect 303418 526046 303488 526102
rect 303168 525978 303488 526046
rect 303168 525922 303238 525978
rect 303294 525922 303362 525978
rect 303418 525922 303488 525978
rect 303168 525888 303488 525922
rect 264908 518420 264964 518430
rect 264908 512596 264964 518364
rect 287808 514350 288128 514384
rect 287808 514294 287878 514350
rect 287934 514294 288002 514350
rect 288058 514294 288128 514350
rect 287808 514226 288128 514294
rect 287808 514170 287878 514226
rect 287934 514170 288002 514226
rect 288058 514170 288128 514226
rect 287808 514102 288128 514170
rect 287808 514046 287878 514102
rect 287934 514046 288002 514102
rect 288058 514046 288128 514102
rect 287808 513978 288128 514046
rect 287808 513922 287878 513978
rect 287934 513922 288002 513978
rect 288058 513922 288128 513978
rect 287808 513888 288128 513922
rect 318528 514350 318848 514384
rect 318528 514294 318598 514350
rect 318654 514294 318722 514350
rect 318778 514294 318848 514350
rect 318528 514226 318848 514294
rect 318528 514170 318598 514226
rect 318654 514170 318722 514226
rect 318778 514170 318848 514226
rect 318528 514102 318848 514170
rect 318528 514046 318598 514102
rect 318654 514046 318722 514102
rect 318778 514046 318848 514102
rect 318528 513978 318848 514046
rect 318528 513922 318598 513978
rect 318654 513922 318722 513978
rect 318778 513922 318848 513978
rect 318528 513888 318848 513922
rect 264908 512530 264964 512540
rect 272448 508350 272768 508384
rect 272448 508294 272518 508350
rect 272574 508294 272642 508350
rect 272698 508294 272768 508350
rect 272448 508226 272768 508294
rect 272448 508170 272518 508226
rect 272574 508170 272642 508226
rect 272698 508170 272768 508226
rect 272448 508102 272768 508170
rect 272448 508046 272518 508102
rect 272574 508046 272642 508102
rect 272698 508046 272768 508102
rect 272448 507978 272768 508046
rect 272448 507922 272518 507978
rect 272574 507922 272642 507978
rect 272698 507922 272768 507978
rect 272448 507888 272768 507922
rect 303168 508350 303488 508384
rect 303168 508294 303238 508350
rect 303294 508294 303362 508350
rect 303418 508294 303488 508350
rect 303168 508226 303488 508294
rect 303168 508170 303238 508226
rect 303294 508170 303362 508226
rect 303418 508170 303488 508226
rect 303168 508102 303488 508170
rect 303168 508046 303238 508102
rect 303294 508046 303362 508102
rect 303418 508046 303488 508102
rect 303168 507978 303488 508046
rect 303168 507922 303238 507978
rect 303294 507922 303362 507978
rect 303418 507922 303488 507978
rect 303168 507888 303488 507922
rect 264572 499650 264628 499660
rect 264684 504868 264740 504878
rect 263900 497970 263956 497980
rect 263116 481730 263172 481740
rect 264684 478996 264740 504812
rect 287808 496350 288128 496384
rect 287808 496294 287878 496350
rect 287934 496294 288002 496350
rect 288058 496294 288128 496350
rect 287808 496226 288128 496294
rect 287808 496170 287878 496226
rect 287934 496170 288002 496226
rect 288058 496170 288128 496226
rect 287808 496102 288128 496170
rect 287808 496046 287878 496102
rect 287934 496046 288002 496102
rect 288058 496046 288128 496102
rect 287808 495978 288128 496046
rect 287808 495922 287878 495978
rect 287934 495922 288002 495978
rect 288058 495922 288128 495978
rect 287808 495888 288128 495922
rect 318528 496350 318848 496384
rect 318528 496294 318598 496350
rect 318654 496294 318722 496350
rect 318778 496294 318848 496350
rect 318528 496226 318848 496294
rect 318528 496170 318598 496226
rect 318654 496170 318722 496226
rect 318778 496170 318848 496226
rect 318528 496102 318848 496170
rect 318528 496046 318598 496102
rect 318654 496046 318722 496102
rect 318778 496046 318848 496102
rect 318528 495978 318848 496046
rect 318528 495922 318598 495978
rect 318654 495922 318722 495978
rect 318778 495922 318848 495978
rect 318528 495888 318848 495922
rect 272448 490350 272768 490384
rect 272448 490294 272518 490350
rect 272574 490294 272642 490350
rect 272698 490294 272768 490350
rect 272448 490226 272768 490294
rect 272448 490170 272518 490226
rect 272574 490170 272642 490226
rect 272698 490170 272768 490226
rect 272448 490102 272768 490170
rect 272448 490046 272518 490102
rect 272574 490046 272642 490102
rect 272698 490046 272768 490102
rect 272448 489978 272768 490046
rect 272448 489922 272518 489978
rect 272574 489922 272642 489978
rect 272698 489922 272768 489978
rect 272448 489888 272768 489922
rect 303168 490350 303488 490384
rect 303168 490294 303238 490350
rect 303294 490294 303362 490350
rect 303418 490294 303488 490350
rect 303168 490226 303488 490294
rect 303168 490170 303238 490226
rect 303294 490170 303362 490226
rect 303418 490170 303488 490226
rect 303168 490102 303488 490170
rect 303168 490046 303238 490102
rect 303294 490046 303362 490102
rect 303418 490046 303488 490102
rect 303168 489978 303488 490046
rect 303168 489922 303238 489978
rect 303294 489922 303362 489978
rect 303418 489922 303488 489978
rect 303168 489888 303488 489922
rect 264684 478930 264740 478940
rect 287808 478350 288128 478384
rect 287808 478294 287878 478350
rect 287934 478294 288002 478350
rect 288058 478294 288128 478350
rect 287808 478226 288128 478294
rect 287808 478170 287878 478226
rect 287934 478170 288002 478226
rect 288058 478170 288128 478226
rect 287808 478102 288128 478170
rect 287808 478046 287878 478102
rect 287934 478046 288002 478102
rect 288058 478046 288128 478102
rect 287808 477978 288128 478046
rect 287808 477922 287878 477978
rect 287934 477922 288002 477978
rect 288058 477922 288128 477978
rect 287808 477888 288128 477922
rect 318528 478350 318848 478384
rect 318528 478294 318598 478350
rect 318654 478294 318722 478350
rect 318778 478294 318848 478350
rect 318528 478226 318848 478294
rect 318528 478170 318598 478226
rect 318654 478170 318722 478226
rect 318778 478170 318848 478226
rect 318528 478102 318848 478170
rect 318528 478046 318598 478102
rect 318654 478046 318722 478102
rect 318778 478046 318848 478102
rect 318528 477978 318848 478046
rect 318528 477922 318598 477978
rect 318654 477922 318722 477978
rect 318778 477922 318848 477978
rect 318528 477888 318848 477922
rect 264572 476308 264628 476318
rect 263788 473698 263844 473708
rect 263788 473396 263844 473642
rect 263788 473330 263844 473340
rect 264124 469558 264180 469568
rect 264012 467938 264068 467948
rect 263900 466228 263956 466238
rect 263788 465238 263844 465248
rect 263788 464996 263844 465182
rect 263788 464930 263844 464940
rect 263788 463618 263844 463628
rect 263788 462756 263844 463562
rect 263900 463316 263956 466172
rect 263900 463250 263956 463260
rect 263788 462690 263844 462700
rect 264012 461636 264068 467882
rect 264012 461570 264068 461580
rect 264124 460516 264180 469502
rect 264124 460450 264180 460460
rect 263900 457940 263956 457950
rect 263788 456148 263844 456158
rect 263788 452676 263844 456092
rect 263900 453796 263956 457884
rect 263900 453730 263956 453740
rect 263788 452610 263844 452620
rect 262892 437490 262948 437500
rect 264572 436436 264628 476252
rect 264684 474598 264740 474608
rect 264684 463876 264740 474542
rect 272448 472350 272768 472384
rect 272448 472294 272518 472350
rect 272574 472294 272642 472350
rect 272698 472294 272768 472350
rect 272448 472226 272768 472294
rect 272448 472170 272518 472226
rect 272574 472170 272642 472226
rect 272698 472170 272768 472226
rect 272448 472102 272768 472170
rect 272448 472046 272518 472102
rect 272574 472046 272642 472102
rect 272698 472046 272768 472102
rect 272448 471978 272768 472046
rect 272448 471922 272518 471978
rect 272574 471922 272642 471978
rect 272698 471922 272768 471978
rect 272448 471888 272768 471922
rect 303168 472350 303488 472384
rect 303168 472294 303238 472350
rect 303294 472294 303362 472350
rect 303418 472294 303488 472350
rect 303168 472226 303488 472294
rect 303168 472170 303238 472226
rect 303294 472170 303362 472226
rect 303418 472170 303488 472226
rect 303168 472102 303488 472170
rect 303168 472046 303238 472102
rect 303294 472046 303362 472102
rect 303418 472046 303488 472102
rect 303168 471978 303488 472046
rect 303168 471922 303238 471978
rect 303294 471922 303362 471978
rect 303418 471922 303488 471978
rect 303168 471888 303488 471922
rect 264684 463810 264740 463820
rect 287808 460350 288128 460384
rect 287808 460294 287878 460350
rect 287934 460294 288002 460350
rect 288058 460294 288128 460350
rect 287808 460226 288128 460294
rect 287808 460170 287878 460226
rect 287934 460170 288002 460226
rect 288058 460170 288128 460226
rect 287808 460102 288128 460170
rect 287808 460046 287878 460102
rect 287934 460046 288002 460102
rect 288058 460046 288128 460102
rect 287808 459978 288128 460046
rect 287808 459922 287878 459978
rect 287934 459922 288002 459978
rect 288058 459922 288128 459978
rect 287808 459888 288128 459922
rect 318528 460350 318848 460384
rect 318528 460294 318598 460350
rect 318654 460294 318722 460350
rect 318778 460294 318848 460350
rect 318528 460226 318848 460294
rect 318528 460170 318598 460226
rect 318654 460170 318722 460226
rect 318778 460170 318848 460226
rect 318528 460102 318848 460170
rect 318528 460046 318598 460102
rect 318654 460046 318722 460102
rect 318778 460046 318848 460102
rect 318528 459978 318848 460046
rect 318528 459922 318598 459978
rect 318654 459922 318722 459978
rect 318778 459922 318848 459978
rect 318528 459888 318848 459922
rect 264684 457828 264740 457838
rect 264684 442596 264740 457772
rect 272448 454350 272768 454384
rect 272448 454294 272518 454350
rect 272574 454294 272642 454350
rect 272698 454294 272768 454350
rect 272448 454226 272768 454294
rect 272448 454170 272518 454226
rect 272574 454170 272642 454226
rect 272698 454170 272768 454226
rect 272448 454102 272768 454170
rect 272448 454046 272518 454102
rect 272574 454046 272642 454102
rect 272698 454046 272768 454102
rect 272448 453978 272768 454046
rect 272448 453922 272518 453978
rect 272574 453922 272642 453978
rect 272698 453922 272768 453978
rect 272448 453888 272768 453922
rect 303168 454350 303488 454384
rect 303168 454294 303238 454350
rect 303294 454294 303362 454350
rect 303418 454294 303488 454350
rect 303168 454226 303488 454294
rect 303168 454170 303238 454226
rect 303294 454170 303362 454226
rect 303418 454170 303488 454226
rect 303168 454102 303488 454170
rect 303168 454046 303238 454102
rect 303294 454046 303362 454102
rect 303418 454046 303488 454102
rect 303168 453978 303488 454046
rect 303168 453922 303238 453978
rect 303294 453922 303362 453978
rect 303418 453922 303488 453978
rect 303168 453888 303488 453922
rect 264908 451108 264964 451118
rect 264908 443156 264964 451052
rect 264908 443090 264964 443100
rect 264684 442530 264740 442540
rect 287808 442350 288128 442384
rect 287808 442294 287878 442350
rect 287934 442294 288002 442350
rect 288058 442294 288128 442350
rect 287808 442226 288128 442294
rect 287808 442170 287878 442226
rect 287934 442170 288002 442226
rect 288058 442170 288128 442226
rect 287808 442102 288128 442170
rect 287808 442046 287878 442102
rect 287934 442046 288002 442102
rect 288058 442046 288128 442102
rect 287808 441978 288128 442046
rect 287808 441922 287878 441978
rect 287934 441922 288002 441978
rect 288058 441922 288128 441978
rect 287808 441888 288128 441922
rect 318528 442350 318848 442384
rect 318528 442294 318598 442350
rect 318654 442294 318722 442350
rect 318778 442294 318848 442350
rect 318528 442226 318848 442294
rect 318528 442170 318598 442226
rect 318654 442170 318722 442226
rect 318778 442170 318848 442226
rect 318528 442102 318848 442170
rect 318528 442046 318598 442102
rect 318654 442046 318722 442102
rect 318778 442046 318848 442102
rect 318528 441978 318848 442046
rect 318528 441922 318598 441978
rect 318654 441922 318722 441978
rect 318778 441922 318848 441978
rect 318528 441888 318848 441922
rect 264572 436370 264628 436380
rect 264684 439572 264740 439582
rect 263340 434420 263396 434430
rect 263340 425796 263396 434364
rect 263340 425730 263396 425740
rect 264572 434308 264628 434318
rect 261324 423490 261380 423500
rect 261212 420130 261268 420140
rect 256172 419010 256228 419020
rect 264572 418516 264628 434252
rect 264572 418450 264628 418460
rect 264684 416276 264740 439516
rect 272448 436350 272768 436384
rect 272448 436294 272518 436350
rect 272574 436294 272642 436350
rect 272698 436294 272768 436350
rect 272448 436226 272768 436294
rect 272448 436170 272518 436226
rect 272574 436170 272642 436226
rect 272698 436170 272768 436226
rect 272448 436102 272768 436170
rect 272448 436046 272518 436102
rect 272574 436046 272642 436102
rect 272698 436046 272768 436102
rect 272448 435978 272768 436046
rect 272448 435922 272518 435978
rect 272574 435922 272642 435978
rect 272698 435922 272768 435978
rect 272448 435888 272768 435922
rect 303168 436350 303488 436384
rect 303168 436294 303238 436350
rect 303294 436294 303362 436350
rect 303418 436294 303488 436350
rect 303168 436226 303488 436294
rect 303168 436170 303238 436226
rect 303294 436170 303362 436226
rect 303418 436170 303488 436226
rect 303168 436102 303488 436170
rect 303168 436046 303238 436102
rect 303294 436046 303362 436102
rect 303418 436046 303488 436102
rect 303168 435978 303488 436046
rect 303168 435922 303238 435978
rect 303294 435922 303362 435978
rect 303418 435922 303488 435978
rect 303168 435888 303488 435922
rect 287808 424350 288128 424384
rect 287808 424294 287878 424350
rect 287934 424294 288002 424350
rect 288058 424294 288128 424350
rect 287808 424226 288128 424294
rect 287808 424170 287878 424226
rect 287934 424170 288002 424226
rect 288058 424170 288128 424226
rect 287808 424102 288128 424170
rect 287808 424046 287878 424102
rect 287934 424046 288002 424102
rect 288058 424046 288128 424102
rect 287808 423978 288128 424046
rect 287808 423922 287878 423978
rect 287934 423922 288002 423978
rect 288058 423922 288128 423978
rect 287808 423888 288128 423922
rect 318528 424350 318848 424384
rect 318528 424294 318598 424350
rect 318654 424294 318722 424350
rect 318778 424294 318848 424350
rect 318528 424226 318848 424294
rect 318528 424170 318598 424226
rect 318654 424170 318722 424226
rect 318778 424170 318848 424226
rect 318528 424102 318848 424170
rect 318528 424046 318598 424102
rect 318654 424046 318722 424102
rect 318778 424046 318848 424102
rect 318528 423978 318848 424046
rect 318528 423922 318598 423978
rect 318654 423922 318722 423978
rect 318778 423922 318848 423978
rect 318528 423888 318848 423922
rect 272448 418350 272768 418384
rect 272448 418294 272518 418350
rect 272574 418294 272642 418350
rect 272698 418294 272768 418350
rect 272448 418226 272768 418294
rect 272448 418170 272518 418226
rect 272574 418170 272642 418226
rect 272698 418170 272768 418226
rect 272448 418102 272768 418170
rect 272448 418046 272518 418102
rect 272574 418046 272642 418102
rect 272698 418046 272768 418102
rect 272448 417978 272768 418046
rect 272448 417922 272518 417978
rect 272574 417922 272642 417978
rect 272698 417922 272768 417978
rect 272448 417888 272768 417922
rect 303168 418350 303488 418384
rect 303168 418294 303238 418350
rect 303294 418294 303362 418350
rect 303418 418294 303488 418350
rect 303168 418226 303488 418294
rect 303168 418170 303238 418226
rect 303294 418170 303362 418226
rect 303418 418170 303488 418226
rect 303168 418102 303488 418170
rect 303168 418046 303238 418102
rect 303294 418046 303362 418102
rect 303418 418046 303488 418102
rect 303168 417978 303488 418046
rect 303168 417922 303238 417978
rect 303294 417922 303362 417978
rect 303418 417922 303488 417978
rect 303168 417888 303488 417922
rect 264684 416210 264740 416220
rect 263900 415156 263956 415166
rect 260316 415018 260372 415028
rect 260316 408996 260372 414962
rect 262892 414036 262948 414046
rect 262108 412132 262164 412142
rect 262108 410676 262164 412076
rect 262108 410610 262164 410620
rect 260316 408930 260372 408940
rect 254898 406294 254994 406350
rect 255050 406294 255118 406350
rect 255174 406294 255242 406350
rect 255298 406294 255366 406350
rect 255422 406294 255518 406350
rect 254898 406226 255518 406294
rect 254898 406170 254994 406226
rect 255050 406170 255118 406226
rect 255174 406170 255242 406226
rect 255298 406170 255366 406226
rect 255422 406170 255518 406226
rect 254898 406102 255518 406170
rect 252812 403442 252868 403452
rect 253148 406084 253204 406094
rect 251178 400294 251274 400350
rect 251330 400294 251398 400350
rect 251454 400294 251522 400350
rect 251578 400294 251646 400350
rect 251702 400294 251798 400350
rect 251178 400226 251798 400294
rect 251178 400170 251274 400226
rect 251330 400170 251398 400226
rect 251454 400170 251522 400226
rect 251578 400170 251646 400226
rect 251702 400170 251798 400226
rect 251178 400102 251798 400170
rect 251178 400046 251274 400102
rect 251330 400046 251398 400102
rect 251454 400046 251522 400102
rect 251578 400046 251646 400102
rect 251702 400046 251798 400102
rect 251178 399978 251798 400046
rect 251178 399922 251274 399978
rect 251330 399922 251398 399978
rect 251454 399922 251522 399978
rect 251578 399922 251646 399978
rect 251702 399922 251798 399978
rect 224178 388294 224274 388350
rect 224330 388294 224398 388350
rect 224454 388294 224522 388350
rect 224578 388294 224646 388350
rect 224702 388294 224798 388350
rect 224178 388226 224798 388294
rect 225808 388389 226128 388446
rect 225808 388333 225836 388389
rect 225892 388333 225940 388389
rect 225996 388333 226044 388389
rect 226100 388333 226128 388389
rect 225808 388276 226128 388333
rect 224178 388170 224274 388226
rect 224330 388170 224398 388226
rect 224454 388170 224522 388226
rect 224578 388170 224646 388226
rect 224702 388170 224798 388226
rect 224178 388102 224798 388170
rect 224178 388046 224274 388102
rect 224330 388046 224398 388102
rect 224454 388046 224522 388102
rect 224578 388046 224646 388102
rect 224702 388046 224798 388102
rect 224178 387978 224798 388046
rect 224178 387922 224274 387978
rect 224330 387922 224398 387978
rect 224454 387922 224522 387978
rect 224578 387922 224646 387978
rect 224702 387922 224798 387978
rect 224178 370350 224798 387922
rect 224178 370294 224274 370350
rect 224330 370294 224398 370350
rect 224454 370294 224522 370350
rect 224578 370294 224646 370350
rect 224702 370294 224798 370350
rect 224178 370226 224798 370294
rect 224178 370170 224274 370226
rect 224330 370170 224398 370226
rect 224454 370170 224522 370226
rect 224578 370170 224646 370226
rect 224702 370170 224798 370226
rect 224178 370102 224798 370170
rect 224178 370046 224274 370102
rect 224330 370046 224398 370102
rect 224454 370046 224522 370102
rect 224578 370046 224646 370102
rect 224702 370046 224798 370102
rect 224178 369978 224798 370046
rect 224178 369922 224274 369978
rect 224330 369922 224398 369978
rect 224454 369922 224522 369978
rect 224578 369922 224646 369978
rect 224702 369922 224798 369978
rect 224178 352350 224798 369922
rect 251178 382350 251798 399922
rect 253148 388948 253204 406028
rect 253148 388882 253204 388892
rect 254898 406046 254994 406102
rect 255050 406046 255118 406102
rect 255174 406046 255242 406102
rect 255298 406046 255366 406102
rect 255422 406046 255518 406102
rect 254898 405978 255518 406046
rect 254898 405922 254994 405978
rect 255050 405922 255118 405978
rect 255174 405922 255242 405978
rect 255298 405922 255366 405978
rect 255422 405922 255518 405978
rect 251178 382294 251274 382350
rect 251330 382294 251398 382350
rect 251454 382294 251522 382350
rect 251578 382294 251646 382350
rect 251702 382294 251798 382350
rect 251178 382226 251798 382294
rect 251178 382170 251274 382226
rect 251330 382170 251398 382226
rect 251454 382170 251522 382226
rect 251578 382170 251646 382226
rect 251702 382170 251798 382226
rect 251178 382102 251798 382170
rect 251178 382046 251274 382102
rect 251330 382046 251398 382102
rect 251454 382046 251522 382102
rect 251578 382046 251646 382102
rect 251702 382046 251798 382102
rect 251178 381978 251798 382046
rect 251178 381922 251274 381978
rect 251330 381922 251398 381978
rect 251454 381922 251522 381978
rect 251578 381922 251646 381978
rect 251702 381922 251798 381978
rect 251178 364350 251798 381922
rect 251178 364294 251274 364350
rect 251330 364294 251398 364350
rect 251454 364294 251522 364350
rect 251578 364294 251646 364350
rect 251702 364294 251798 364350
rect 251178 364226 251798 364294
rect 251178 364170 251274 364226
rect 251330 364170 251398 364226
rect 251454 364170 251522 364226
rect 251578 364170 251646 364226
rect 251702 364170 251798 364226
rect 251178 364102 251798 364170
rect 251178 364046 251274 364102
rect 251330 364046 251398 364102
rect 251454 364046 251522 364102
rect 251578 364046 251646 364102
rect 251702 364046 251798 364102
rect 251178 363978 251798 364046
rect 251178 363922 251274 363978
rect 251330 363922 251398 363978
rect 251454 363922 251522 363978
rect 251578 363922 251646 363978
rect 251702 363922 251798 363978
rect 224178 352294 224274 352350
rect 224330 352294 224398 352350
rect 224454 352294 224522 352350
rect 224578 352294 224646 352350
rect 224702 352294 224798 352350
rect 224178 352226 224798 352294
rect 224178 352170 224274 352226
rect 224330 352170 224398 352226
rect 224454 352170 224522 352226
rect 224578 352170 224646 352226
rect 224702 352170 224798 352226
rect 224178 352102 224798 352170
rect 224178 352046 224274 352102
rect 224330 352046 224398 352102
rect 224454 352046 224522 352102
rect 224578 352046 224646 352102
rect 224702 352046 224798 352102
rect 224178 351978 224798 352046
rect 224178 351922 224274 351978
rect 224330 351922 224398 351978
rect 224454 351922 224522 351978
rect 224578 351922 224646 351978
rect 224702 351922 224798 351978
rect 224178 334350 224798 351922
rect 225808 352350 226128 352384
rect 225808 352294 225878 352350
rect 225934 352294 226002 352350
rect 226058 352294 226128 352350
rect 225808 352226 226128 352294
rect 225808 352170 225878 352226
rect 225934 352170 226002 352226
rect 226058 352170 226128 352226
rect 225808 352102 226128 352170
rect 225808 352046 225878 352102
rect 225934 352046 226002 352102
rect 226058 352046 226128 352102
rect 225808 351978 226128 352046
rect 225808 351922 225878 351978
rect 225934 351922 226002 351978
rect 226058 351922 226128 351978
rect 225808 351888 226128 351922
rect 241168 346350 241488 346384
rect 241168 346294 241238 346350
rect 241294 346294 241362 346350
rect 241418 346294 241488 346350
rect 241168 346226 241488 346294
rect 241168 346170 241238 346226
rect 241294 346170 241362 346226
rect 241418 346170 241488 346226
rect 241168 346102 241488 346170
rect 241168 346046 241238 346102
rect 241294 346046 241362 346102
rect 241418 346046 241488 346102
rect 241168 345978 241488 346046
rect 241168 345922 241238 345978
rect 241294 345922 241362 345978
rect 241418 345922 241488 345978
rect 241168 345888 241488 345922
rect 251178 346350 251798 363922
rect 251178 346294 251274 346350
rect 251330 346294 251398 346350
rect 251454 346294 251522 346350
rect 251578 346294 251646 346350
rect 251702 346294 251798 346350
rect 251178 346226 251798 346294
rect 251178 346170 251274 346226
rect 251330 346170 251398 346226
rect 251454 346170 251522 346226
rect 251578 346170 251646 346226
rect 251702 346170 251798 346226
rect 251178 346102 251798 346170
rect 251178 346046 251274 346102
rect 251330 346046 251398 346102
rect 251454 346046 251522 346102
rect 251578 346046 251646 346102
rect 251702 346046 251798 346102
rect 251178 345978 251798 346046
rect 251178 345922 251274 345978
rect 251330 345922 251398 345978
rect 251454 345922 251522 345978
rect 251578 345922 251646 345978
rect 251702 345922 251798 345978
rect 224178 334294 224274 334350
rect 224330 334294 224398 334350
rect 224454 334294 224522 334350
rect 224578 334294 224646 334350
rect 224702 334294 224798 334350
rect 224178 334226 224798 334294
rect 224178 334170 224274 334226
rect 224330 334170 224398 334226
rect 224454 334170 224522 334226
rect 224578 334170 224646 334226
rect 224702 334170 224798 334226
rect 224178 334102 224798 334170
rect 224178 334046 224274 334102
rect 224330 334046 224398 334102
rect 224454 334046 224522 334102
rect 224578 334046 224646 334102
rect 224702 334046 224798 334102
rect 224178 333978 224798 334046
rect 224178 333922 224274 333978
rect 224330 333922 224398 333978
rect 224454 333922 224522 333978
rect 224578 333922 224646 333978
rect 224702 333922 224798 333978
rect 224178 316350 224798 333922
rect 225808 334350 226128 334384
rect 225808 334294 225878 334350
rect 225934 334294 226002 334350
rect 226058 334294 226128 334350
rect 225808 334226 226128 334294
rect 225808 334170 225878 334226
rect 225934 334170 226002 334226
rect 226058 334170 226128 334226
rect 225808 334102 226128 334170
rect 225808 334046 225878 334102
rect 225934 334046 226002 334102
rect 226058 334046 226128 334102
rect 225808 333978 226128 334046
rect 225808 333922 225878 333978
rect 225934 333922 226002 333978
rect 226058 333922 226128 333978
rect 225808 333888 226128 333922
rect 251020 334292 251076 334302
rect 241168 328350 241488 328384
rect 241168 328294 241238 328350
rect 241294 328294 241362 328350
rect 241418 328294 241488 328350
rect 241168 328226 241488 328294
rect 241168 328170 241238 328226
rect 241294 328170 241362 328226
rect 241418 328170 241488 328226
rect 241168 328102 241488 328170
rect 241168 328046 241238 328102
rect 241294 328046 241362 328102
rect 241418 328046 241488 328102
rect 241168 327978 241488 328046
rect 241168 327922 241238 327978
rect 241294 327922 241362 327978
rect 241418 327922 241488 327978
rect 241168 327888 241488 327922
rect 251020 324996 251076 334236
rect 251020 324930 251076 324940
rect 251178 328350 251798 345922
rect 254898 388350 255518 405922
rect 254898 388294 254994 388350
rect 255050 388294 255118 388350
rect 255174 388294 255242 388350
rect 255298 388294 255366 388350
rect 255422 388294 255518 388350
rect 254898 388226 255518 388294
rect 254898 388170 254994 388226
rect 255050 388170 255118 388226
rect 255174 388170 255242 388226
rect 255298 388170 255366 388226
rect 255422 388170 255518 388226
rect 254898 388102 255518 388170
rect 254898 388046 254994 388102
rect 255050 388046 255118 388102
rect 255174 388046 255242 388102
rect 255298 388046 255366 388102
rect 255422 388046 255518 388102
rect 254898 387978 255518 388046
rect 254898 387922 254994 387978
rect 255050 387922 255118 387978
rect 255174 387922 255242 387978
rect 255298 387922 255366 387978
rect 255422 387922 255518 387978
rect 254898 370350 255518 387922
rect 256172 407428 256228 407438
rect 256172 378756 256228 407372
rect 259532 406756 259588 406766
rect 259532 386372 259588 406700
rect 260316 406756 260372 406766
rect 260316 404578 260372 406700
rect 262220 406738 262276 406748
rect 262108 406196 262164 406206
rect 262108 404758 262164 406140
rect 262108 404692 262164 404702
rect 260316 404512 260372 404522
rect 259532 386306 259588 386316
rect 259644 402724 259700 402734
rect 259644 383236 259700 402668
rect 262108 400596 262164 400606
rect 262108 399538 262164 400540
rect 262220 400036 262276 406682
rect 262892 403396 262948 413980
rect 263340 413476 263396 413486
rect 263340 408100 263396 413420
rect 263788 412916 263844 412926
rect 263788 411778 263844 412860
rect 263788 411712 263844 411722
rect 263900 410228 263956 415100
rect 263900 410162 263956 410172
rect 263340 408034 263396 408044
rect 263452 408358 263508 408368
rect 263452 403956 263508 408302
rect 263788 407316 263844 407326
rect 263788 406918 263844 407260
rect 263788 406852 263844 406862
rect 263900 407098 263956 407108
rect 263900 405076 263956 407042
rect 287808 406350 288128 406384
rect 287808 406294 287878 406350
rect 287934 406294 288002 406350
rect 288058 406294 288128 406350
rect 287808 406226 288128 406294
rect 287808 406170 287878 406226
rect 287934 406170 288002 406226
rect 288058 406170 288128 406226
rect 287808 406102 288128 406170
rect 287808 406046 287878 406102
rect 287934 406046 288002 406102
rect 288058 406046 288128 406102
rect 287808 405978 288128 406046
rect 287808 405922 287878 405978
rect 287934 405922 288002 405978
rect 288058 405922 288128 405978
rect 287808 405888 288128 405922
rect 318528 406350 318848 406384
rect 318528 406294 318598 406350
rect 318654 406294 318722 406350
rect 318778 406294 318848 406350
rect 318528 406226 318848 406294
rect 318528 406170 318598 406226
rect 318654 406170 318722 406226
rect 318778 406170 318848 406226
rect 318528 406102 318848 406170
rect 318528 406046 318598 406102
rect 318654 406046 318722 406102
rect 318778 406046 318848 406102
rect 318528 405978 318848 406046
rect 318528 405922 318598 405978
rect 318654 405922 318722 405978
rect 318778 405922 318848 405978
rect 318528 405888 318848 405922
rect 263900 405010 263956 405020
rect 263788 404516 263844 404526
rect 263788 404038 263844 404460
rect 263788 403972 263844 403982
rect 263452 403890 263508 403900
rect 262892 403330 262948 403340
rect 263788 403138 263844 403148
rect 263788 402836 263844 403082
rect 263788 402770 263844 402780
rect 263900 402958 263956 402968
rect 263900 401716 263956 402902
rect 263900 401650 263956 401660
rect 262220 399970 262276 399980
rect 272448 400350 272768 400384
rect 272448 400294 272518 400350
rect 272574 400294 272642 400350
rect 272698 400294 272768 400350
rect 272448 400226 272768 400294
rect 272448 400170 272518 400226
rect 272574 400170 272642 400226
rect 272698 400170 272768 400226
rect 272448 400102 272768 400170
rect 272448 400046 272518 400102
rect 272574 400046 272642 400102
rect 272698 400046 272768 400102
rect 272448 399978 272768 400046
rect 272448 399922 272518 399978
rect 272574 399922 272642 399978
rect 272698 399922 272768 399978
rect 272448 399888 272768 399922
rect 303168 400350 303488 400384
rect 303168 400294 303238 400350
rect 303294 400294 303362 400350
rect 303418 400294 303488 400350
rect 303168 400226 303488 400294
rect 303168 400170 303238 400226
rect 303294 400170 303362 400226
rect 303418 400170 303488 400226
rect 303168 400102 303488 400170
rect 303168 400046 303238 400102
rect 303294 400046 303362 400102
rect 303418 400046 303488 400102
rect 303168 399978 303488 400046
rect 303168 399922 303238 399978
rect 303294 399922 303362 399978
rect 303418 399922 303488 399978
rect 303168 399888 303488 399922
rect 262108 399472 262164 399482
rect 263788 399718 263844 399728
rect 263788 398356 263844 399662
rect 263788 398290 263844 398300
rect 263788 398098 263844 398108
rect 263788 397796 263844 398042
rect 263788 397730 263844 397740
rect 263788 396478 263844 396488
rect 263788 395556 263844 396422
rect 263788 395490 263844 395500
rect 263900 396298 263956 396308
rect 263900 394996 263956 396242
rect 263900 394930 263956 394940
rect 263788 393058 263844 393068
rect 263788 392756 263844 393002
rect 263788 392690 263844 392700
rect 263788 391438 263844 391448
rect 263788 391076 263844 391382
rect 263788 391010 263844 391020
rect 263900 390516 263956 390526
rect 263788 389956 263844 389966
rect 263788 387940 263844 389900
rect 263900 388052 263956 390460
rect 263900 387986 263956 387996
rect 265020 388948 265076 388958
rect 263788 387874 263844 387884
rect 259644 383170 259700 383180
rect 263788 386372 263844 386382
rect 263788 382676 263844 386316
rect 263788 382610 263844 382620
rect 265020 382116 265076 388892
rect 287808 388350 288128 388384
rect 287808 388294 287878 388350
rect 287934 388294 288002 388350
rect 288058 388294 288128 388350
rect 287808 388226 288128 388294
rect 287808 388170 287878 388226
rect 287934 388170 288002 388226
rect 288058 388170 288128 388226
rect 287808 388102 288128 388170
rect 287808 388046 287878 388102
rect 287934 388046 288002 388102
rect 288058 388046 288128 388102
rect 287808 387978 288128 388046
rect 287808 387922 287878 387978
rect 287934 387922 288002 387978
rect 288058 387922 288128 387978
rect 287808 387888 288128 387922
rect 318528 388350 318848 388384
rect 318528 388294 318598 388350
rect 318654 388294 318722 388350
rect 318778 388294 318848 388350
rect 318528 388226 318848 388294
rect 318528 388170 318598 388226
rect 318654 388170 318722 388226
rect 318778 388170 318848 388226
rect 318528 388102 318848 388170
rect 318528 388046 318598 388102
rect 318654 388046 318722 388102
rect 318778 388046 318848 388102
rect 318528 387978 318848 388046
rect 318528 387922 318598 387978
rect 318654 387922 318722 387978
rect 318778 387922 318848 387978
rect 318528 387888 318848 387922
rect 265020 382050 265076 382060
rect 272448 382350 272768 382384
rect 272448 382294 272518 382350
rect 272574 382294 272642 382350
rect 272698 382294 272768 382350
rect 272448 382226 272768 382294
rect 272448 382170 272518 382226
rect 272574 382170 272642 382226
rect 272698 382170 272768 382226
rect 272448 382102 272768 382170
rect 272448 382046 272518 382102
rect 272574 382046 272642 382102
rect 272698 382046 272768 382102
rect 272448 381978 272768 382046
rect 272448 381922 272518 381978
rect 272574 381922 272642 381978
rect 272698 381922 272768 381978
rect 272448 381888 272768 381922
rect 303168 382350 303488 382384
rect 303168 382294 303238 382350
rect 303294 382294 303362 382350
rect 303418 382294 303488 382350
rect 303168 382226 303488 382294
rect 303168 382170 303238 382226
rect 303294 382170 303362 382226
rect 303418 382170 303488 382226
rect 303168 382102 303488 382170
rect 303168 382046 303238 382102
rect 303294 382046 303362 382102
rect 303418 382046 303488 382102
rect 303168 381978 303488 382046
rect 303168 381922 303238 381978
rect 303294 381922 303362 381978
rect 303418 381922 303488 381978
rect 303168 381888 303488 381922
rect 264908 380772 264964 380782
rect 264796 379092 264852 379102
rect 256172 378690 256228 378700
rect 257852 378980 257908 378990
rect 254898 370294 254994 370350
rect 255050 370294 255118 370350
rect 255174 370294 255242 370350
rect 255298 370294 255366 370350
rect 255422 370294 255518 370350
rect 254898 370226 255518 370294
rect 254898 370170 254994 370226
rect 255050 370170 255118 370226
rect 255174 370170 255242 370226
rect 255298 370170 255366 370226
rect 255422 370170 255518 370226
rect 254898 370102 255518 370170
rect 254898 370046 254994 370102
rect 255050 370046 255118 370102
rect 255174 370046 255242 370102
rect 255298 370046 255366 370102
rect 255422 370046 255518 370102
rect 254898 369978 255518 370046
rect 254898 369922 254994 369978
rect 255050 369922 255118 369978
rect 255174 369922 255242 369978
rect 255298 369922 255366 369978
rect 255422 369922 255518 369978
rect 254898 352350 255518 369922
rect 257852 363636 257908 378924
rect 264572 378868 264628 378878
rect 257852 363570 257908 363580
rect 263788 372148 263844 372158
rect 263788 363076 263844 372092
rect 263788 363010 263844 363020
rect 264572 357476 264628 378812
rect 264684 377188 264740 377198
rect 264684 361396 264740 377132
rect 264684 361330 264740 361340
rect 264796 358596 264852 379036
rect 264908 370356 264964 380716
rect 264908 370290 264964 370300
rect 287808 370350 288128 370384
rect 287808 370294 287878 370350
rect 287934 370294 288002 370350
rect 288058 370294 288128 370350
rect 287808 370226 288128 370294
rect 287808 370170 287878 370226
rect 287934 370170 288002 370226
rect 288058 370170 288128 370226
rect 287808 370102 288128 370170
rect 287808 370046 287878 370102
rect 287934 370046 288002 370102
rect 288058 370046 288128 370102
rect 287808 369978 288128 370046
rect 287808 369922 287878 369978
rect 287934 369922 288002 369978
rect 288058 369922 288128 369978
rect 287808 369888 288128 369922
rect 318528 370350 318848 370384
rect 318528 370294 318598 370350
rect 318654 370294 318722 370350
rect 318778 370294 318848 370350
rect 318528 370226 318848 370294
rect 318528 370170 318598 370226
rect 318654 370170 318722 370226
rect 318778 370170 318848 370226
rect 318528 370102 318848 370170
rect 318528 370046 318598 370102
rect 318654 370046 318722 370102
rect 318778 370046 318848 370102
rect 318528 369978 318848 370046
rect 318528 369922 318598 369978
rect 318654 369922 318722 369978
rect 318778 369922 318848 369978
rect 318528 369888 318848 369922
rect 272448 364350 272768 364384
rect 272448 364294 272518 364350
rect 272574 364294 272642 364350
rect 272698 364294 272768 364350
rect 272448 364226 272768 364294
rect 272448 364170 272518 364226
rect 272574 364170 272642 364226
rect 272698 364170 272768 364226
rect 272448 364102 272768 364170
rect 272448 364046 272518 364102
rect 272574 364046 272642 364102
rect 272698 364046 272768 364102
rect 272448 363978 272768 364046
rect 272448 363922 272518 363978
rect 272574 363922 272642 363978
rect 272698 363922 272768 363978
rect 272448 363888 272768 363922
rect 303168 364350 303488 364384
rect 303168 364294 303238 364350
rect 303294 364294 303362 364350
rect 303418 364294 303488 364350
rect 303168 364226 303488 364294
rect 303168 364170 303238 364226
rect 303294 364170 303362 364226
rect 303418 364170 303488 364226
rect 303168 364102 303488 364170
rect 303168 364046 303238 364102
rect 303294 364046 303362 364102
rect 303418 364046 303488 364102
rect 303168 363978 303488 364046
rect 303168 363922 303238 363978
rect 303294 363922 303362 363978
rect 303418 363922 303488 363978
rect 303168 363888 303488 363922
rect 264796 358530 264852 358540
rect 264572 357410 264628 357420
rect 264796 355236 264852 355246
rect 254898 352294 254994 352350
rect 255050 352294 255118 352350
rect 255174 352294 255242 352350
rect 255298 352294 255366 352350
rect 255422 352294 255518 352350
rect 254898 352226 255518 352294
rect 254898 352170 254994 352226
rect 255050 352170 255118 352226
rect 255174 352170 255242 352226
rect 255298 352170 255366 352226
rect 255422 352170 255518 352226
rect 254898 352102 255518 352170
rect 254898 352046 254994 352102
rect 255050 352046 255118 352102
rect 255174 352046 255242 352102
rect 255298 352046 255366 352102
rect 255422 352046 255518 352102
rect 254898 351978 255518 352046
rect 254898 351922 254994 351978
rect 255050 351922 255118 351978
rect 255174 351922 255242 351978
rect 255298 351922 255366 351978
rect 255422 351922 255518 351978
rect 254898 334350 255518 351922
rect 264572 352436 264628 352446
rect 263340 351876 263396 351886
rect 263340 348598 263396 351820
rect 263788 350196 263844 350206
rect 263788 349498 263844 350140
rect 263788 349432 263844 349442
rect 263340 348532 263396 348542
rect 263788 347956 263844 347966
rect 263788 347878 263844 347900
rect 263788 347812 263844 347822
rect 260092 347396 260148 347406
rect 260092 338518 260148 347340
rect 262108 346276 262164 346286
rect 262108 343558 262164 346220
rect 263788 345716 263844 345726
rect 263788 344638 263844 345660
rect 263788 344572 263844 344582
rect 263900 345156 263956 345166
rect 263900 344458 263956 345100
rect 263900 344392 263956 344402
rect 262108 343492 262164 343502
rect 263788 344036 263844 344046
rect 263788 343018 263844 343980
rect 263788 342952 263844 342962
rect 263788 342356 263844 342366
rect 263788 341758 263844 342300
rect 263788 341692 263844 341702
rect 263900 341578 263956 341588
rect 263788 341398 263844 341408
rect 263788 341236 263844 341342
rect 263788 341170 263844 341180
rect 263900 340676 263956 341522
rect 263900 340610 263956 340620
rect 263788 340498 263844 340508
rect 260092 338452 260148 338462
rect 260316 340318 260372 340328
rect 260316 335076 260372 340262
rect 263788 339556 263844 340442
rect 264572 340340 264628 352380
rect 264572 340274 264628 340284
rect 264684 342838 264740 342848
rect 263788 339490 263844 339500
rect 260316 335010 260372 335020
rect 261212 337652 261268 337662
rect 254898 334294 254994 334350
rect 255050 334294 255118 334350
rect 255174 334294 255242 334350
rect 255298 334294 255366 334350
rect 255422 334294 255518 334350
rect 254898 334226 255518 334294
rect 254898 334170 254994 334226
rect 255050 334170 255118 334226
rect 255174 334170 255242 334226
rect 255298 334170 255366 334226
rect 255422 334170 255518 334226
rect 254898 334102 255518 334170
rect 254898 334046 254994 334102
rect 255050 334046 255118 334102
rect 255174 334046 255242 334102
rect 255298 334046 255366 334102
rect 255422 334046 255518 334102
rect 254898 333978 255518 334046
rect 254898 333922 254994 333978
rect 255050 333922 255118 333978
rect 255174 333922 255242 333978
rect 255298 333922 255366 333978
rect 255422 333922 255518 333978
rect 251178 328294 251274 328350
rect 251330 328294 251398 328350
rect 251454 328294 251522 328350
rect 251578 328294 251646 328350
rect 251702 328294 251798 328350
rect 251178 328226 251798 328294
rect 251178 328170 251274 328226
rect 251330 328170 251398 328226
rect 251454 328170 251522 328226
rect 251578 328170 251646 328226
rect 251702 328170 251798 328226
rect 251178 328102 251798 328170
rect 251178 328046 251274 328102
rect 251330 328046 251398 328102
rect 251454 328046 251522 328102
rect 251578 328046 251646 328102
rect 251702 328046 251798 328102
rect 251178 327978 251798 328046
rect 251178 327922 251274 327978
rect 251330 327922 251398 327978
rect 251454 327922 251522 327978
rect 251578 327922 251646 327978
rect 251702 327922 251798 327978
rect 224178 316294 224274 316350
rect 224330 316294 224398 316350
rect 224454 316294 224522 316350
rect 224578 316294 224646 316350
rect 224702 316294 224798 316350
rect 224178 316226 224798 316294
rect 224178 316170 224274 316226
rect 224330 316170 224398 316226
rect 224454 316170 224522 316226
rect 224578 316170 224646 316226
rect 224702 316170 224798 316226
rect 224178 316102 224798 316170
rect 224178 316046 224274 316102
rect 224330 316046 224398 316102
rect 224454 316046 224522 316102
rect 224578 316046 224646 316102
rect 224702 316046 224798 316102
rect 224178 315978 224798 316046
rect 224178 315922 224274 315978
rect 224330 315922 224398 315978
rect 224454 315922 224522 315978
rect 224578 315922 224646 315978
rect 224702 315922 224798 315978
rect 224178 298350 224798 315922
rect 224178 298294 224274 298350
rect 224330 298294 224398 298350
rect 224454 298294 224522 298350
rect 224578 298294 224646 298350
rect 224702 298294 224798 298350
rect 224178 298226 224798 298294
rect 224178 298170 224274 298226
rect 224330 298170 224398 298226
rect 224454 298170 224522 298226
rect 224578 298170 224646 298226
rect 224702 298170 224798 298226
rect 224178 298102 224798 298170
rect 224178 298046 224274 298102
rect 224330 298046 224398 298102
rect 224454 298046 224522 298102
rect 224578 298046 224646 298102
rect 224702 298046 224798 298102
rect 224178 297978 224798 298046
rect 224178 297922 224274 297978
rect 224330 297922 224398 297978
rect 224454 297922 224522 297978
rect 224578 297922 224646 297978
rect 224702 297922 224798 297978
rect 224178 280350 224798 297922
rect 251178 310350 251798 327922
rect 251916 330260 251972 330270
rect 251916 321636 251972 330204
rect 251916 321570 251972 321580
rect 251178 310294 251274 310350
rect 251330 310294 251398 310350
rect 251454 310294 251522 310350
rect 251578 310294 251646 310350
rect 251702 310294 251798 310350
rect 251178 310226 251798 310294
rect 251178 310170 251274 310226
rect 251330 310170 251398 310226
rect 251454 310170 251522 310226
rect 251578 310170 251646 310226
rect 251702 310170 251798 310226
rect 251178 310102 251798 310170
rect 251178 310046 251274 310102
rect 251330 310046 251398 310102
rect 251454 310046 251522 310102
rect 251578 310046 251646 310102
rect 251702 310046 251798 310102
rect 251178 309978 251798 310046
rect 251178 309922 251274 309978
rect 251330 309922 251398 309978
rect 251454 309922 251522 309978
rect 251578 309922 251646 309978
rect 251702 309922 251798 309978
rect 251178 292350 251798 309922
rect 254898 316350 255518 333922
rect 259532 329588 259588 329598
rect 259532 322756 259588 329532
rect 259532 322690 259588 322700
rect 261212 322196 261268 337596
rect 264572 336756 264628 336766
rect 264012 335636 264068 335646
rect 263788 332836 263844 332846
rect 261212 322130 261268 322140
rect 261324 332276 261380 332286
rect 261324 320516 261380 332220
rect 263788 331498 263844 332780
rect 263788 331432 263844 331442
rect 263900 331716 263956 331726
rect 263788 331156 263844 331166
rect 263788 330958 263844 331100
rect 263900 331138 263956 331660
rect 263900 331072 263956 331082
rect 263788 330892 263844 330902
rect 264012 330778 264068 335580
rect 264012 330712 264068 330722
rect 263788 330598 263844 330634
rect 263788 330530 263844 330540
rect 263900 328916 263956 328926
rect 263788 327796 263844 327806
rect 263788 327538 263844 327740
rect 263788 327472 263844 327482
rect 263900 327358 263956 328860
rect 263900 327292 263956 327302
rect 264572 325738 264628 336700
rect 264684 333396 264740 342782
rect 264796 336308 264852 355180
rect 265132 352996 265188 353006
rect 265132 336980 265188 352940
rect 287808 352350 288128 352384
rect 287808 352294 287878 352350
rect 287934 352294 288002 352350
rect 288058 352294 288128 352350
rect 287808 352226 288128 352294
rect 287808 352170 287878 352226
rect 287934 352170 288002 352226
rect 288058 352170 288128 352226
rect 287808 352102 288128 352170
rect 287808 352046 287878 352102
rect 287934 352046 288002 352102
rect 288058 352046 288128 352102
rect 287808 351978 288128 352046
rect 287808 351922 287878 351978
rect 287934 351922 288002 351978
rect 288058 351922 288128 351978
rect 287808 351888 288128 351922
rect 318528 352350 318848 352384
rect 318528 352294 318598 352350
rect 318654 352294 318722 352350
rect 318778 352294 318848 352350
rect 318528 352226 318848 352294
rect 318528 352170 318598 352226
rect 318654 352170 318722 352226
rect 318778 352170 318848 352226
rect 318528 352102 318848 352170
rect 318528 352046 318598 352102
rect 318654 352046 318722 352102
rect 318778 352046 318848 352102
rect 318528 351978 318848 352046
rect 318528 351922 318598 351978
rect 318654 351922 318722 351978
rect 318778 351922 318848 351978
rect 318528 351888 318848 351922
rect 272448 346350 272768 346384
rect 272448 346294 272518 346350
rect 272574 346294 272642 346350
rect 272698 346294 272768 346350
rect 272448 346226 272768 346294
rect 272448 346170 272518 346226
rect 272574 346170 272642 346226
rect 272698 346170 272768 346226
rect 272448 346102 272768 346170
rect 272448 346046 272518 346102
rect 272574 346046 272642 346102
rect 272698 346046 272768 346102
rect 272448 345978 272768 346046
rect 272448 345922 272518 345978
rect 272574 345922 272642 345978
rect 272698 345922 272768 345978
rect 272448 345888 272768 345922
rect 303168 346350 303488 346384
rect 303168 346294 303238 346350
rect 303294 346294 303362 346350
rect 303418 346294 303488 346350
rect 303168 346226 303488 346294
rect 303168 346170 303238 346226
rect 303294 346170 303362 346226
rect 303418 346170 303488 346226
rect 303168 346102 303488 346170
rect 303168 346046 303238 346102
rect 303294 346046 303362 346102
rect 303418 346046 303488 346102
rect 303168 345978 303488 346046
rect 303168 345922 303238 345978
rect 303294 345922 303362 345978
rect 303418 345922 303488 345978
rect 303168 345888 303488 345922
rect 265132 336914 265188 336924
rect 264796 336242 264852 336252
rect 287808 334350 288128 334384
rect 287808 334294 287878 334350
rect 287934 334294 288002 334350
rect 288058 334294 288128 334350
rect 287808 334226 288128 334294
rect 287808 334170 287878 334226
rect 287934 334170 288002 334226
rect 288058 334170 288128 334226
rect 287808 334102 288128 334170
rect 287808 334046 287878 334102
rect 287934 334046 288002 334102
rect 288058 334046 288128 334102
rect 287808 333978 288128 334046
rect 264684 333330 264740 333340
rect 264908 333956 264964 333966
rect 264908 325918 264964 333900
rect 287808 333922 287878 333978
rect 287934 333922 288002 333978
rect 288058 333922 288128 333978
rect 287808 333888 288128 333922
rect 318528 334350 318848 334384
rect 318528 334294 318598 334350
rect 318654 334294 318722 334350
rect 318778 334294 318848 334350
rect 318528 334226 318848 334294
rect 318528 334170 318598 334226
rect 318654 334170 318722 334226
rect 318778 334170 318848 334226
rect 318528 334102 318848 334170
rect 318528 334046 318598 334102
rect 318654 334046 318722 334102
rect 318778 334046 318848 334102
rect 318528 333978 318848 334046
rect 318528 333922 318598 333978
rect 318654 333922 318722 333978
rect 318778 333922 318848 333978
rect 318528 333888 318848 333922
rect 272448 328350 272768 328384
rect 272448 328294 272518 328350
rect 272574 328294 272642 328350
rect 272698 328294 272768 328350
rect 272448 328226 272768 328294
rect 272448 328170 272518 328226
rect 272574 328170 272642 328226
rect 272698 328170 272768 328226
rect 272448 328102 272768 328170
rect 272448 328046 272518 328102
rect 272574 328046 272642 328102
rect 272698 328046 272768 328102
rect 272448 327978 272768 328046
rect 272448 327922 272518 327978
rect 272574 327922 272642 327978
rect 272698 327922 272768 327978
rect 272448 327888 272768 327922
rect 303168 328350 303488 328384
rect 303168 328294 303238 328350
rect 303294 328294 303362 328350
rect 303418 328294 303488 328350
rect 303168 328226 303488 328294
rect 303168 328170 303238 328226
rect 303294 328170 303362 328226
rect 303418 328170 303488 328226
rect 303168 328102 303488 328170
rect 303168 328046 303238 328102
rect 303294 328046 303362 328102
rect 303418 328046 303488 328102
rect 303168 327978 303488 328046
rect 303168 327922 303238 327978
rect 303294 327922 303362 327978
rect 303418 327922 303488 327978
rect 303168 327888 303488 327922
rect 264908 325852 264964 325862
rect 264572 325672 264628 325682
rect 263788 325558 263844 325594
rect 263788 325490 263844 325500
rect 263788 324118 263844 324128
rect 263788 323876 263844 324062
rect 263788 323810 263844 323820
rect 261324 320450 261380 320460
rect 254898 316294 254994 316350
rect 255050 316294 255118 316350
rect 255174 316294 255242 316350
rect 255298 316294 255366 316350
rect 255422 316294 255518 316350
rect 254898 316226 255518 316294
rect 254898 316170 254994 316226
rect 255050 316170 255118 316226
rect 255174 316170 255242 316226
rect 255298 316170 255366 316226
rect 255422 316170 255518 316226
rect 254898 316102 255518 316170
rect 254898 316046 254994 316102
rect 255050 316046 255118 316102
rect 255174 316046 255242 316102
rect 255298 316046 255366 316102
rect 255422 316046 255518 316102
rect 254898 315978 255518 316046
rect 254898 315922 254994 315978
rect 255050 315922 255118 315978
rect 255174 315922 255242 315978
rect 255298 315922 255366 315978
rect 255422 315922 255518 315978
rect 254898 298350 255518 315922
rect 287808 316350 288128 316384
rect 287808 316294 287878 316350
rect 287934 316294 288002 316350
rect 288058 316294 288128 316350
rect 287808 316226 288128 316294
rect 287808 316170 287878 316226
rect 287934 316170 288002 316226
rect 288058 316170 288128 316226
rect 287808 316102 288128 316170
rect 287808 316046 287878 316102
rect 287934 316046 288002 316102
rect 288058 316046 288128 316102
rect 287808 315978 288128 316046
rect 287808 315922 287878 315978
rect 287934 315922 288002 315978
rect 288058 315922 288128 315978
rect 287808 315888 288128 315922
rect 318528 316350 318848 316384
rect 318528 316294 318598 316350
rect 318654 316294 318722 316350
rect 318778 316294 318848 316350
rect 318528 316226 318848 316294
rect 318528 316170 318598 316226
rect 318654 316170 318722 316226
rect 318778 316170 318848 316226
rect 318528 316102 318848 316170
rect 318528 316046 318598 316102
rect 318654 316046 318722 316102
rect 318778 316046 318848 316102
rect 318528 315978 318848 316046
rect 318528 315922 318598 315978
rect 318654 315922 318722 315978
rect 318778 315922 318848 315978
rect 318528 315888 318848 315922
rect 261436 314580 261492 314590
rect 261436 314356 261492 314524
rect 261436 314290 261492 314300
rect 272448 310350 272768 310384
rect 272448 310294 272518 310350
rect 272574 310294 272642 310350
rect 272698 310294 272768 310350
rect 272448 310226 272768 310294
rect 272448 310170 272518 310226
rect 272574 310170 272642 310226
rect 272698 310170 272768 310226
rect 272448 310102 272768 310170
rect 272448 310046 272518 310102
rect 272574 310046 272642 310102
rect 272698 310046 272768 310102
rect 272448 309978 272768 310046
rect 272448 309922 272518 309978
rect 272574 309922 272642 309978
rect 272698 309922 272768 309978
rect 272448 309888 272768 309922
rect 303168 310350 303488 310384
rect 303168 310294 303238 310350
rect 303294 310294 303362 310350
rect 303418 310294 303488 310350
rect 303168 310226 303488 310294
rect 303168 310170 303238 310226
rect 303294 310170 303362 310226
rect 303418 310170 303488 310226
rect 303168 310102 303488 310170
rect 303168 310046 303238 310102
rect 303294 310046 303362 310102
rect 303418 310046 303488 310102
rect 303168 309978 303488 310046
rect 303168 309922 303238 309978
rect 303294 309922 303362 309978
rect 303418 309922 303488 309978
rect 303168 309888 303488 309922
rect 263788 308308 263844 308318
rect 263788 304276 263844 308252
rect 263788 304210 263844 304220
rect 254898 298294 254994 298350
rect 255050 298294 255118 298350
rect 255174 298294 255242 298350
rect 255298 298294 255366 298350
rect 255422 298294 255518 298350
rect 254898 298226 255518 298294
rect 254898 298170 254994 298226
rect 255050 298170 255118 298226
rect 255174 298170 255242 298226
rect 255298 298170 255366 298226
rect 255422 298170 255518 298226
rect 254898 298102 255518 298170
rect 254898 298046 254994 298102
rect 255050 298046 255118 298102
rect 255174 298046 255242 298102
rect 255298 298046 255366 298102
rect 255422 298046 255518 298102
rect 254898 297978 255518 298046
rect 254898 297922 254994 297978
rect 255050 297922 255118 297978
rect 255174 297922 255242 297978
rect 255298 297922 255366 297978
rect 255422 297922 255518 297978
rect 251178 292294 251274 292350
rect 251330 292294 251398 292350
rect 251454 292294 251522 292350
rect 251578 292294 251646 292350
rect 251702 292294 251798 292350
rect 251178 292226 251798 292294
rect 251178 292170 251274 292226
rect 251330 292170 251398 292226
rect 251454 292170 251522 292226
rect 251578 292170 251646 292226
rect 251702 292170 251798 292226
rect 251178 292102 251798 292170
rect 251178 292046 251274 292102
rect 251330 292046 251398 292102
rect 251454 292046 251522 292102
rect 251578 292046 251646 292102
rect 251702 292046 251798 292102
rect 251178 291978 251798 292046
rect 251178 291922 251274 291978
rect 251330 291922 251398 291978
rect 251454 291922 251522 291978
rect 251578 291922 251646 291978
rect 251702 291922 251798 291978
rect 224178 280294 224274 280350
rect 224330 280294 224398 280350
rect 224454 280294 224522 280350
rect 224578 280294 224646 280350
rect 224702 280294 224798 280350
rect 224178 280226 224798 280294
rect 224178 280170 224274 280226
rect 224330 280170 224398 280226
rect 224454 280170 224522 280226
rect 224578 280170 224646 280226
rect 224702 280170 224798 280226
rect 224178 280102 224798 280170
rect 224178 280046 224274 280102
rect 224330 280046 224398 280102
rect 224454 280046 224522 280102
rect 224578 280046 224646 280102
rect 224702 280046 224798 280102
rect 224178 279978 224798 280046
rect 224178 279922 224274 279978
rect 224330 279922 224398 279978
rect 224454 279922 224522 279978
rect 224578 279922 224646 279978
rect 224702 279922 224798 279978
rect 224178 262350 224798 279922
rect 225808 280350 226128 280384
rect 225808 280294 225878 280350
rect 225934 280294 226002 280350
rect 226058 280294 226128 280350
rect 225808 280226 226128 280294
rect 225808 280170 225878 280226
rect 225934 280170 226002 280226
rect 226058 280170 226128 280226
rect 225808 280102 226128 280170
rect 225808 280046 225878 280102
rect 225934 280046 226002 280102
rect 226058 280046 226128 280102
rect 225808 279978 226128 280046
rect 225808 279922 225878 279978
rect 225934 279922 226002 279978
rect 226058 279922 226128 279978
rect 225808 279888 226128 279922
rect 249452 275156 249508 275166
rect 241168 274350 241488 274384
rect 241168 274294 241238 274350
rect 241294 274294 241362 274350
rect 241418 274294 241488 274350
rect 241168 274226 241488 274294
rect 241168 274170 241238 274226
rect 241294 274170 241362 274226
rect 241418 274170 241488 274226
rect 241168 274102 241488 274170
rect 241168 274046 241238 274102
rect 241294 274046 241362 274102
rect 241418 274046 241488 274102
rect 241168 273978 241488 274046
rect 241168 273922 241238 273978
rect 241294 273922 241362 273978
rect 241418 273922 241488 273978
rect 241168 273888 241488 273922
rect 249452 268678 249508 275100
rect 249452 268612 249508 268622
rect 251178 274350 251798 291922
rect 251178 274294 251274 274350
rect 251330 274294 251398 274350
rect 251454 274294 251522 274350
rect 251578 274294 251646 274350
rect 251702 274294 251798 274350
rect 251178 274226 251798 274294
rect 251178 274170 251274 274226
rect 251330 274170 251398 274226
rect 251454 274170 251522 274226
rect 251578 274170 251646 274226
rect 251702 274170 251798 274226
rect 251178 274102 251798 274170
rect 251178 274046 251274 274102
rect 251330 274046 251398 274102
rect 251454 274046 251522 274102
rect 251578 274046 251646 274102
rect 251702 274046 251798 274102
rect 251178 273978 251798 274046
rect 251178 273922 251274 273978
rect 251330 273922 251398 273978
rect 251454 273922 251522 273978
rect 251578 273922 251646 273978
rect 251702 273922 251798 273978
rect 224178 262294 224274 262350
rect 224330 262294 224398 262350
rect 224454 262294 224522 262350
rect 224578 262294 224646 262350
rect 224702 262294 224798 262350
rect 224178 262226 224798 262294
rect 224178 262170 224274 262226
rect 224330 262170 224398 262226
rect 224454 262170 224522 262226
rect 224578 262170 224646 262226
rect 224702 262170 224798 262226
rect 224178 262102 224798 262170
rect 224178 262046 224274 262102
rect 224330 262046 224398 262102
rect 224454 262046 224522 262102
rect 224578 262046 224646 262102
rect 224702 262046 224798 262102
rect 224178 261978 224798 262046
rect 224178 261922 224274 261978
rect 224330 261922 224398 261978
rect 224454 261922 224522 261978
rect 224578 261922 224646 261978
rect 224702 261922 224798 261978
rect 224178 244350 224798 261922
rect 225808 262350 226128 262384
rect 225808 262294 225878 262350
rect 225934 262294 226002 262350
rect 226058 262294 226128 262350
rect 225808 262226 226128 262294
rect 225808 262170 225878 262226
rect 225934 262170 226002 262226
rect 226058 262170 226128 262226
rect 225808 262102 226128 262170
rect 225808 262046 225878 262102
rect 225934 262046 226002 262102
rect 226058 262046 226128 262102
rect 225808 261978 226128 262046
rect 225808 261922 225878 261978
rect 225934 261922 226002 261978
rect 226058 261922 226128 261978
rect 225808 261888 226128 261922
rect 241168 256350 241488 256384
rect 241168 256294 241238 256350
rect 241294 256294 241362 256350
rect 241418 256294 241488 256350
rect 241168 256226 241488 256294
rect 241168 256170 241238 256226
rect 241294 256170 241362 256226
rect 241418 256170 241488 256226
rect 241168 256102 241488 256170
rect 241168 256046 241238 256102
rect 241294 256046 241362 256102
rect 241418 256046 241488 256102
rect 241168 255978 241488 256046
rect 241168 255922 241238 255978
rect 241294 255922 241362 255978
rect 241418 255922 241488 255978
rect 241168 255888 241488 255922
rect 251178 256350 251798 273922
rect 252812 292516 252868 292526
rect 252812 258356 252868 292460
rect 252812 258290 252868 258300
rect 254898 280350 255518 297922
rect 264572 298676 264628 298686
rect 263788 290836 263844 290846
rect 263788 289828 263844 290780
rect 263788 289762 263844 289772
rect 263788 285796 263844 285806
rect 254898 280294 254994 280350
rect 255050 280294 255118 280350
rect 255174 280294 255242 280350
rect 255298 280294 255366 280350
rect 255422 280294 255518 280350
rect 254898 280226 255518 280294
rect 254898 280170 254994 280226
rect 255050 280170 255118 280226
rect 255174 280170 255242 280226
rect 255298 280170 255366 280226
rect 255422 280170 255518 280226
rect 254898 280102 255518 280170
rect 254898 280046 254994 280102
rect 255050 280046 255118 280102
rect 255174 280046 255242 280102
rect 255298 280046 255366 280102
rect 255422 280046 255518 280102
rect 254898 279978 255518 280046
rect 254898 279922 254994 279978
rect 255050 279922 255118 279978
rect 255174 279922 255242 279978
rect 255298 279922 255366 279978
rect 255422 279922 255518 279978
rect 254898 262350 255518 279922
rect 259532 285684 259588 285694
rect 259532 266420 259588 285628
rect 261212 284900 261268 284910
rect 261212 284452 261268 284844
rect 261212 284386 261268 284396
rect 263788 283220 263844 285740
rect 264572 285684 264628 298620
rect 287808 298350 288128 298384
rect 287808 298294 287878 298350
rect 287934 298294 288002 298350
rect 288058 298294 288128 298350
rect 287808 298226 288128 298294
rect 287808 298170 287878 298226
rect 287934 298170 288002 298226
rect 288058 298170 288128 298226
rect 287808 298102 288128 298170
rect 287808 298046 287878 298102
rect 287934 298046 288002 298102
rect 288058 298046 288128 298102
rect 287808 297978 288128 298046
rect 287808 297922 287878 297978
rect 287934 297922 288002 297978
rect 288058 297922 288128 297978
rect 287808 297888 288128 297922
rect 318528 298350 318848 298384
rect 318528 298294 318598 298350
rect 318654 298294 318722 298350
rect 318778 298294 318848 298350
rect 318528 298226 318848 298294
rect 318528 298170 318598 298226
rect 318654 298170 318722 298226
rect 318778 298170 318848 298226
rect 318528 298102 318848 298170
rect 318528 298046 318598 298102
rect 318654 298046 318722 298102
rect 318778 298046 318848 298102
rect 318528 297978 318848 298046
rect 318528 297922 318598 297978
rect 318654 297922 318722 297978
rect 318778 297922 318848 297978
rect 318528 297888 318848 297922
rect 272448 292350 272768 292384
rect 272448 292294 272518 292350
rect 272574 292294 272642 292350
rect 272698 292294 272768 292350
rect 272448 292226 272768 292294
rect 272448 292170 272518 292226
rect 272574 292170 272642 292226
rect 272698 292170 272768 292226
rect 272448 292102 272768 292170
rect 272448 292046 272518 292102
rect 272574 292046 272642 292102
rect 272698 292046 272768 292102
rect 272448 291978 272768 292046
rect 272448 291922 272518 291978
rect 272574 291922 272642 291978
rect 272698 291922 272768 291978
rect 272448 291888 272768 291922
rect 303168 292350 303488 292384
rect 303168 292294 303238 292350
rect 303294 292294 303362 292350
rect 303418 292294 303488 292350
rect 303168 292226 303488 292294
rect 303168 292170 303238 292226
rect 303294 292170 303362 292226
rect 303418 292170 303488 292226
rect 303168 292102 303488 292170
rect 303168 292046 303238 292102
rect 303294 292046 303362 292102
rect 303418 292046 303488 292102
rect 303168 291978 303488 292046
rect 303168 291922 303238 291978
rect 303294 291922 303362 291978
rect 303418 291922 303488 291978
rect 303168 291888 303488 291922
rect 264572 285618 264628 285628
rect 263788 283154 263844 283164
rect 287808 280350 288128 280384
rect 287808 280294 287878 280350
rect 287934 280294 288002 280350
rect 288058 280294 288128 280350
rect 287808 280226 288128 280294
rect 287808 280170 287878 280226
rect 287934 280170 288002 280226
rect 288058 280170 288128 280226
rect 287808 280102 288128 280170
rect 287808 280046 287878 280102
rect 287934 280046 288002 280102
rect 288058 280046 288128 280102
rect 287808 279978 288128 280046
rect 287808 279922 287878 279978
rect 287934 279922 288002 279978
rect 288058 279922 288128 279978
rect 287808 279888 288128 279922
rect 318528 280350 318848 280384
rect 318528 280294 318598 280350
rect 318654 280294 318722 280350
rect 318778 280294 318848 280350
rect 318528 280226 318848 280294
rect 318528 280170 318598 280226
rect 318654 280170 318722 280226
rect 318778 280170 318848 280226
rect 318528 280102 318848 280170
rect 318528 280046 318598 280102
rect 318654 280046 318722 280102
rect 318778 280046 318848 280102
rect 318528 279978 318848 280046
rect 318528 279922 318598 279978
rect 318654 279922 318722 279978
rect 318778 279922 318848 279978
rect 318528 279888 318848 279922
rect 263788 279636 263844 279646
rect 263340 279076 263396 279086
rect 263340 278038 263396 279020
rect 263788 278218 263844 279580
rect 263788 278152 263844 278162
rect 263340 277972 263396 277982
rect 262108 277396 262164 277406
rect 262108 276418 262164 277340
rect 262108 276352 262164 276362
rect 263788 276836 263844 276846
rect 262220 275716 262276 275726
rect 262220 272998 262276 275660
rect 263788 275698 263844 276780
rect 263788 275632 263844 275642
rect 272448 274350 272768 274384
rect 272448 274294 272518 274350
rect 272574 274294 272642 274350
rect 272698 274294 272768 274350
rect 272448 274226 272768 274294
rect 272448 274170 272518 274226
rect 272574 274170 272642 274226
rect 272698 274170 272768 274226
rect 272448 274102 272768 274170
rect 272448 274046 272518 274102
rect 272574 274046 272642 274102
rect 272698 274046 272768 274102
rect 272448 273978 272768 274046
rect 272448 273922 272518 273978
rect 272574 273922 272642 273978
rect 272698 273922 272768 273978
rect 272448 273888 272768 273922
rect 303168 274350 303488 274384
rect 303168 274294 303238 274350
rect 303294 274294 303362 274350
rect 303418 274294 303488 274350
rect 303168 274226 303488 274294
rect 303168 274170 303238 274226
rect 303294 274170 303362 274226
rect 303418 274170 303488 274226
rect 303168 274102 303488 274170
rect 303168 274046 303238 274102
rect 303294 274046 303362 274102
rect 303418 274046 303488 274102
rect 303168 273978 303488 274046
rect 303168 273922 303238 273978
rect 303294 273922 303362 273978
rect 303418 273922 303488 273978
rect 303168 273888 303488 273922
rect 262220 272932 262276 272942
rect 262108 272916 262164 272926
rect 262108 270298 262164 272860
rect 263788 272356 263844 272366
rect 263788 271558 263844 272300
rect 263788 271492 263844 271502
rect 263900 271796 263956 271806
rect 263900 270838 263956 271740
rect 263900 270772 263956 270782
rect 262108 270232 262164 270242
rect 263788 269556 263844 269566
rect 263788 268858 263844 269500
rect 263788 268792 263844 268802
rect 263788 268498 263844 268508
rect 263788 267876 263844 268442
rect 263788 267810 263844 267820
rect 259532 266354 259588 266364
rect 262444 267092 262500 267102
rect 262220 265748 262276 265758
rect 260316 265636 260372 265646
rect 254898 262294 254994 262350
rect 255050 262294 255118 262350
rect 255174 262294 255242 262350
rect 255298 262294 255366 262350
rect 255422 262294 255518 262350
rect 254898 262226 255518 262294
rect 254898 262170 254994 262226
rect 255050 262170 255118 262226
rect 255174 262170 255242 262226
rect 255298 262170 255366 262226
rect 255422 262170 255518 262226
rect 254898 262102 255518 262170
rect 254898 262046 254994 262102
rect 255050 262046 255118 262102
rect 255174 262046 255242 262102
rect 255298 262046 255366 262102
rect 255422 262046 255518 262102
rect 254898 261978 255518 262046
rect 254898 261922 254994 261978
rect 255050 261922 255118 261978
rect 255174 261922 255242 261978
rect 255298 261922 255366 261978
rect 255422 261922 255518 261978
rect 251178 256294 251274 256350
rect 251330 256294 251398 256350
rect 251454 256294 251522 256350
rect 251578 256294 251646 256350
rect 251702 256294 251798 256350
rect 251178 256226 251798 256294
rect 251178 256170 251274 256226
rect 251330 256170 251398 256226
rect 251454 256170 251522 256226
rect 251578 256170 251646 256226
rect 251702 256170 251798 256226
rect 251178 256102 251798 256170
rect 251178 256046 251274 256102
rect 251330 256046 251398 256102
rect 251454 256046 251522 256102
rect 251578 256046 251646 256102
rect 251702 256046 251798 256102
rect 251178 255978 251798 256046
rect 251178 255922 251274 255978
rect 251330 255922 251398 255978
rect 251454 255922 251522 255978
rect 251578 255922 251646 255978
rect 251702 255922 251798 255978
rect 224178 244294 224274 244350
rect 224330 244294 224398 244350
rect 224454 244294 224522 244350
rect 224578 244294 224646 244350
rect 224702 244294 224798 244350
rect 224178 244226 224798 244294
rect 224178 244170 224274 244226
rect 224330 244170 224398 244226
rect 224454 244170 224522 244226
rect 224578 244170 224646 244226
rect 224702 244170 224798 244226
rect 224178 244102 224798 244170
rect 224178 244046 224274 244102
rect 224330 244046 224398 244102
rect 224454 244046 224522 244102
rect 224578 244046 224646 244102
rect 224702 244046 224798 244102
rect 224178 243978 224798 244046
rect 224178 243922 224274 243978
rect 224330 243922 224398 243978
rect 224454 243922 224522 243978
rect 224578 243922 224646 243978
rect 224702 243922 224798 243978
rect 224178 226350 224798 243922
rect 248556 239876 248612 239886
rect 248556 234612 248612 239820
rect 248556 234546 248612 234556
rect 251178 238350 251798 255922
rect 251178 238294 251274 238350
rect 251330 238294 251398 238350
rect 251454 238294 251522 238350
rect 251578 238294 251646 238350
rect 251702 238294 251798 238350
rect 251178 238226 251798 238294
rect 251178 238170 251274 238226
rect 251330 238170 251398 238226
rect 251454 238170 251522 238226
rect 251578 238170 251646 238226
rect 251702 238170 251798 238226
rect 251178 238102 251798 238170
rect 251178 238046 251274 238102
rect 251330 238046 251398 238102
rect 251454 238046 251522 238102
rect 251578 238046 251646 238102
rect 251702 238046 251798 238102
rect 251178 237978 251798 238046
rect 251178 237922 251274 237978
rect 251330 237922 251398 237978
rect 251454 237922 251522 237978
rect 251578 237922 251646 237978
rect 251702 237922 251798 237978
rect 224178 226294 224274 226350
rect 224330 226294 224398 226350
rect 224454 226294 224522 226350
rect 224578 226294 224646 226350
rect 224702 226294 224798 226350
rect 224178 226226 224798 226294
rect 224178 226170 224274 226226
rect 224330 226170 224398 226226
rect 224454 226170 224522 226226
rect 224578 226170 224646 226226
rect 224702 226170 224798 226226
rect 224178 226102 224798 226170
rect 224178 226046 224274 226102
rect 224330 226046 224398 226102
rect 224454 226046 224522 226102
rect 224578 226046 224646 226102
rect 224702 226046 224798 226102
rect 224178 225978 224798 226046
rect 224178 225922 224274 225978
rect 224330 225922 224398 225978
rect 224454 225922 224522 225978
rect 224578 225922 224646 225978
rect 224702 225922 224798 225978
rect 224178 208350 224798 225922
rect 251178 220350 251798 237922
rect 251178 220294 251274 220350
rect 251330 220294 251398 220350
rect 251454 220294 251522 220350
rect 251578 220294 251646 220350
rect 251702 220294 251798 220350
rect 251178 220226 251798 220294
rect 251178 220170 251274 220226
rect 251330 220170 251398 220226
rect 251454 220170 251522 220226
rect 251578 220170 251646 220226
rect 251702 220170 251798 220226
rect 251178 220102 251798 220170
rect 251178 220046 251274 220102
rect 251330 220046 251398 220102
rect 251454 220046 251522 220102
rect 251578 220046 251646 220102
rect 251702 220046 251798 220102
rect 251178 219978 251798 220046
rect 251178 219922 251274 219978
rect 251330 219922 251398 219978
rect 251454 219922 251522 219978
rect 251578 219922 251646 219978
rect 251702 219922 251798 219978
rect 231532 212884 231588 212894
rect 231532 212436 231588 212828
rect 231532 212370 231588 212380
rect 231756 212772 231812 212782
rect 231756 212436 231812 212716
rect 231756 212370 231812 212380
rect 224178 208294 224274 208350
rect 224330 208294 224398 208350
rect 224454 208294 224522 208350
rect 224578 208294 224646 208350
rect 224702 208294 224798 208350
rect 224178 208226 224798 208294
rect 224178 208170 224274 208226
rect 224330 208170 224398 208226
rect 224454 208170 224522 208226
rect 224578 208170 224646 208226
rect 224702 208170 224798 208226
rect 224178 208102 224798 208170
rect 224178 208046 224274 208102
rect 224330 208046 224398 208102
rect 224454 208046 224522 208102
rect 224578 208046 224646 208102
rect 224702 208046 224798 208102
rect 224178 207978 224798 208046
rect 224178 207922 224274 207978
rect 224330 207922 224398 207978
rect 224454 207922 224522 207978
rect 224578 207922 224646 207978
rect 224702 207922 224798 207978
rect 224178 190350 224798 207922
rect 225808 208350 226128 208384
rect 225808 208294 225878 208350
rect 225934 208294 226002 208350
rect 226058 208294 226128 208350
rect 225808 208226 226128 208294
rect 225808 208170 225878 208226
rect 225934 208170 226002 208226
rect 226058 208170 226128 208226
rect 225808 208102 226128 208170
rect 225808 208046 225878 208102
rect 225934 208046 226002 208102
rect 226058 208046 226128 208102
rect 225808 207978 226128 208046
rect 225808 207922 225878 207978
rect 225934 207922 226002 207978
rect 226058 207922 226128 207978
rect 225808 207888 226128 207922
rect 241168 202350 241488 202384
rect 241168 202294 241238 202350
rect 241294 202294 241362 202350
rect 241418 202294 241488 202350
rect 241168 202226 241488 202294
rect 241168 202170 241238 202226
rect 241294 202170 241362 202226
rect 241418 202170 241488 202226
rect 241168 202102 241488 202170
rect 241168 202046 241238 202102
rect 241294 202046 241362 202102
rect 241418 202046 241488 202102
rect 241168 201978 241488 202046
rect 241168 201922 241238 201978
rect 241294 201922 241362 201978
rect 241418 201922 241488 201978
rect 241168 201888 241488 201922
rect 251178 202350 251798 219922
rect 254898 244350 255518 261922
rect 259980 264718 260036 264728
rect 259980 257236 260036 264662
rect 260316 261658 260372 265580
rect 260316 261592 260372 261602
rect 262108 262836 262164 262846
rect 262108 261044 262164 262780
rect 262220 261716 262276 265692
rect 262220 261650 262276 261660
rect 262332 263396 262388 263406
rect 262108 260978 262164 260988
rect 262332 259028 262388 263340
rect 262444 261156 262500 267036
rect 263788 267058 263844 267068
rect 263788 266756 263844 267002
rect 263788 266690 263844 266700
rect 263788 266518 263844 266528
rect 263788 266196 263844 266462
rect 263788 266130 263844 266140
rect 262444 261090 262500 261100
rect 262556 264898 262612 264908
rect 262332 258962 262388 258972
rect 259980 257170 260036 257180
rect 262556 256676 262612 264842
rect 264012 264516 264068 264526
rect 263788 260398 263844 260408
rect 263788 260036 263844 260342
rect 263788 259970 263844 259980
rect 263900 260218 263956 260228
rect 263900 259476 263956 260162
rect 263900 259410 263956 259420
rect 263788 258598 263844 258608
rect 263788 258356 263844 258542
rect 263788 258290 263844 258300
rect 263900 258418 263956 258428
rect 263900 257796 263956 258362
rect 263900 257730 263956 257740
rect 264012 257684 264068 264460
rect 287808 262350 288128 262384
rect 287808 262294 287878 262350
rect 287934 262294 288002 262350
rect 288058 262294 288128 262350
rect 287808 262226 288128 262294
rect 287808 262170 287878 262226
rect 287934 262170 288002 262226
rect 288058 262170 288128 262226
rect 287808 262102 288128 262170
rect 287808 262046 287878 262102
rect 287934 262046 288002 262102
rect 288058 262046 288128 262102
rect 287808 261978 288128 262046
rect 287808 261922 287878 261978
rect 287934 261922 288002 261978
rect 288058 261922 288128 261978
rect 287808 261888 288128 261922
rect 318528 262350 318848 262384
rect 318528 262294 318598 262350
rect 318654 262294 318722 262350
rect 318778 262294 318848 262350
rect 318528 262226 318848 262294
rect 318528 262170 318598 262226
rect 318654 262170 318722 262226
rect 318778 262170 318848 262226
rect 318528 262102 318848 262170
rect 318528 262046 318598 262102
rect 318654 262046 318722 262102
rect 318778 262046 318848 262102
rect 318528 261978 318848 262046
rect 318528 261922 318598 261978
rect 318654 261922 318722 261978
rect 318778 261922 318848 261978
rect 318528 261888 318848 261922
rect 264012 257618 264068 257628
rect 262556 256610 262612 256620
rect 272448 256350 272768 256384
rect 272448 256294 272518 256350
rect 272574 256294 272642 256350
rect 272698 256294 272768 256350
rect 272448 256226 272768 256294
rect 272448 256170 272518 256226
rect 272574 256170 272642 256226
rect 272698 256170 272768 256226
rect 272448 256102 272768 256170
rect 272448 256046 272518 256102
rect 272574 256046 272642 256102
rect 272698 256046 272768 256102
rect 272448 255978 272768 256046
rect 272448 255922 272518 255978
rect 272574 255922 272642 255978
rect 272698 255922 272768 255978
rect 272448 255888 272768 255922
rect 303168 256350 303488 256384
rect 303168 256294 303238 256350
rect 303294 256294 303362 256350
rect 303418 256294 303488 256350
rect 303168 256226 303488 256294
rect 303168 256170 303238 256226
rect 303294 256170 303362 256226
rect 303418 256170 303488 256226
rect 303168 256102 303488 256170
rect 303168 256046 303238 256102
rect 303294 256046 303362 256102
rect 303418 256046 303488 256102
rect 303168 255978 303488 256046
rect 303168 255922 303238 255978
rect 303294 255922 303362 255978
rect 303418 255922 303488 255978
rect 303168 255888 303488 255922
rect 263788 255358 263844 255368
rect 260316 254458 260372 254468
rect 260316 248836 260372 254402
rect 263788 253876 263844 255302
rect 263788 253810 263844 253820
rect 263788 253558 263844 253568
rect 263788 253316 263844 253502
rect 263788 253250 263844 253260
rect 263900 253378 263956 253388
rect 263900 252756 263956 253322
rect 263900 252690 263956 252700
rect 263788 251938 263844 251948
rect 263788 251076 263844 251882
rect 263788 251010 263844 251020
rect 263788 250516 263844 250526
rect 263788 250318 263844 250460
rect 263788 250252 263844 250262
rect 260316 248770 260372 248780
rect 254898 244294 254994 244350
rect 255050 244294 255118 244350
rect 255174 244294 255242 244350
rect 255298 244294 255366 244350
rect 255422 244294 255518 244350
rect 254898 244226 255518 244294
rect 254898 244170 254994 244226
rect 255050 244170 255118 244226
rect 255174 244170 255242 244226
rect 255298 244170 255366 244226
rect 255422 244170 255518 244226
rect 254898 244102 255518 244170
rect 254898 244046 254994 244102
rect 255050 244046 255118 244102
rect 255174 244046 255242 244102
rect 255298 244046 255366 244102
rect 255422 244046 255518 244102
rect 254898 243978 255518 244046
rect 254898 243922 254994 243978
rect 255050 243922 255118 243978
rect 255174 243922 255242 243978
rect 255298 243922 255366 243978
rect 255422 243922 255518 243978
rect 254898 226350 255518 243922
rect 287808 244350 288128 244384
rect 287808 244294 287878 244350
rect 287934 244294 288002 244350
rect 288058 244294 288128 244350
rect 287808 244226 288128 244294
rect 287808 244170 287878 244226
rect 287934 244170 288002 244226
rect 288058 244170 288128 244226
rect 287808 244102 288128 244170
rect 287808 244046 287878 244102
rect 287934 244046 288002 244102
rect 288058 244046 288128 244102
rect 287808 243978 288128 244046
rect 287808 243922 287878 243978
rect 287934 243922 288002 243978
rect 288058 243922 288128 243978
rect 287808 243888 288128 243922
rect 318528 244350 318848 244384
rect 318528 244294 318598 244350
rect 318654 244294 318722 244350
rect 318778 244294 318848 244350
rect 318528 244226 318848 244294
rect 318528 244170 318598 244226
rect 318654 244170 318722 244226
rect 318778 244170 318848 244226
rect 318528 244102 318848 244170
rect 318528 244046 318598 244102
rect 318654 244046 318722 244102
rect 318778 244046 318848 244102
rect 318528 243978 318848 244046
rect 318528 243922 318598 243978
rect 318654 243922 318722 243978
rect 318778 243922 318848 243978
rect 318528 243888 318848 243922
rect 263788 239316 263844 239326
rect 263788 236068 263844 239260
rect 263788 236002 263844 236012
rect 263900 238756 263956 238766
rect 257852 235396 257908 235406
rect 254898 226294 254994 226350
rect 255050 226294 255118 226350
rect 255174 226294 255242 226350
rect 255298 226294 255366 226350
rect 255422 226294 255518 226350
rect 254898 226226 255518 226294
rect 254898 226170 254994 226226
rect 255050 226170 255118 226226
rect 255174 226170 255242 226226
rect 255298 226170 255366 226226
rect 255422 226170 255518 226226
rect 254898 226102 255518 226170
rect 254898 226046 254994 226102
rect 255050 226046 255118 226102
rect 255174 226046 255242 226102
rect 255298 226046 255366 226102
rect 255422 226046 255518 226102
rect 254898 225978 255518 226046
rect 254898 225922 254994 225978
rect 255050 225922 255118 225978
rect 255174 225922 255242 225978
rect 255298 225922 255366 225978
rect 255422 225922 255518 225978
rect 252812 215908 252868 215918
rect 251178 202294 251274 202350
rect 251330 202294 251398 202350
rect 251454 202294 251522 202350
rect 251578 202294 251646 202350
rect 251702 202294 251798 202350
rect 251178 202226 251798 202294
rect 251178 202170 251274 202226
rect 251330 202170 251398 202226
rect 251454 202170 251522 202226
rect 251578 202170 251646 202226
rect 251702 202170 251798 202226
rect 251178 202102 251798 202170
rect 251178 202046 251274 202102
rect 251330 202046 251398 202102
rect 251454 202046 251522 202102
rect 251578 202046 251646 202102
rect 251702 202046 251798 202102
rect 251178 201978 251798 202046
rect 251178 201922 251274 201978
rect 251330 201922 251398 201978
rect 251454 201922 251522 201978
rect 251578 201922 251646 201978
rect 251702 201922 251798 201978
rect 248556 196756 248612 196766
rect 248556 196498 248612 196700
rect 248556 196432 248612 196442
rect 248556 194158 248612 194168
rect 224178 190294 224274 190350
rect 224330 190294 224398 190350
rect 224454 190294 224522 190350
rect 224578 190294 224646 190350
rect 224702 190294 224798 190350
rect 224178 190226 224798 190294
rect 224178 190170 224274 190226
rect 224330 190170 224398 190226
rect 224454 190170 224522 190226
rect 224578 190170 224646 190226
rect 224702 190170 224798 190226
rect 224178 190102 224798 190170
rect 224178 190046 224274 190102
rect 224330 190046 224398 190102
rect 224454 190046 224522 190102
rect 224578 190046 224646 190102
rect 224702 190046 224798 190102
rect 224178 189978 224798 190046
rect 224178 189922 224274 189978
rect 224330 189922 224398 189978
rect 224454 189922 224522 189978
rect 224578 189922 224646 189978
rect 224702 189922 224798 189978
rect 224178 172350 224798 189922
rect 225808 190350 226128 190384
rect 225808 190294 225878 190350
rect 225934 190294 226002 190350
rect 226058 190294 226128 190350
rect 225808 190226 226128 190294
rect 225808 190170 225878 190226
rect 225934 190170 226002 190226
rect 226058 190170 226128 190226
rect 225808 190102 226128 190170
rect 225808 190046 225878 190102
rect 225934 190046 226002 190102
rect 226058 190046 226128 190102
rect 225808 189978 226128 190046
rect 225808 189922 225878 189978
rect 225934 189922 226002 189978
rect 226058 189922 226128 189978
rect 225808 189888 226128 189922
rect 248556 184996 248612 194102
rect 248556 184930 248612 184940
rect 241168 184350 241488 184384
rect 241168 184294 241238 184350
rect 241294 184294 241362 184350
rect 241418 184294 241488 184350
rect 241168 184226 241488 184294
rect 241168 184170 241238 184226
rect 241294 184170 241362 184226
rect 241418 184170 241488 184226
rect 241168 184102 241488 184170
rect 241168 184046 241238 184102
rect 241294 184046 241362 184102
rect 241418 184046 241488 184102
rect 241168 183978 241488 184046
rect 241168 183922 241238 183978
rect 241294 183922 241362 183978
rect 241418 183922 241488 183978
rect 241168 183888 241488 183922
rect 251178 184350 251798 201922
rect 251916 209076 251972 209086
rect 251916 187124 251972 209020
rect 252812 190484 252868 215852
rect 252812 190418 252868 190428
rect 254898 208350 255518 225922
rect 254898 208294 254994 208350
rect 255050 208294 255118 208350
rect 255174 208294 255242 208350
rect 255298 208294 255366 208350
rect 255422 208294 255518 208350
rect 254898 208226 255518 208294
rect 254898 208170 254994 208226
rect 255050 208170 255118 208226
rect 255174 208170 255242 208226
rect 255298 208170 255366 208226
rect 255422 208170 255518 208226
rect 254898 208102 255518 208170
rect 254898 208046 254994 208102
rect 255050 208046 255118 208102
rect 255174 208046 255242 208102
rect 255298 208046 255366 208102
rect 255422 208046 255518 208102
rect 254898 207978 255518 208046
rect 254898 207922 254994 207978
rect 255050 207922 255118 207978
rect 255174 207922 255242 207978
rect 255298 207922 255366 207978
rect 255422 207922 255518 207978
rect 251916 187058 251972 187068
rect 254898 190350 255518 207922
rect 256172 234276 256228 234286
rect 256172 191828 256228 234220
rect 256172 191762 256228 191772
rect 254898 190294 254994 190350
rect 255050 190294 255118 190350
rect 255174 190294 255242 190350
rect 255298 190294 255366 190350
rect 255422 190294 255518 190350
rect 254898 190226 255518 190294
rect 254898 190170 254994 190226
rect 255050 190170 255118 190226
rect 255174 190170 255242 190226
rect 255298 190170 255366 190226
rect 255422 190170 255518 190226
rect 254898 190102 255518 190170
rect 254898 190046 254994 190102
rect 255050 190046 255118 190102
rect 255174 190046 255242 190102
rect 255298 190046 255366 190102
rect 255422 190046 255518 190102
rect 254898 189978 255518 190046
rect 254898 189922 254994 189978
rect 255050 189922 255118 189978
rect 255174 189922 255242 189978
rect 255298 189922 255366 189978
rect 255422 189922 255518 189978
rect 251178 184294 251274 184350
rect 251330 184294 251398 184350
rect 251454 184294 251522 184350
rect 251578 184294 251646 184350
rect 251702 184294 251798 184350
rect 251178 184226 251798 184294
rect 251178 184170 251274 184226
rect 251330 184170 251398 184226
rect 251454 184170 251522 184226
rect 251578 184170 251646 184226
rect 251702 184170 251798 184226
rect 251178 184102 251798 184170
rect 251178 184046 251274 184102
rect 251330 184046 251398 184102
rect 251454 184046 251522 184102
rect 251578 184046 251646 184102
rect 251702 184046 251798 184102
rect 251178 183978 251798 184046
rect 251178 183922 251274 183978
rect 251330 183922 251398 183978
rect 251454 183922 251522 183978
rect 251578 183922 251646 183978
rect 251702 183922 251798 183978
rect 224178 172294 224274 172350
rect 224330 172294 224398 172350
rect 224454 172294 224522 172350
rect 224578 172294 224646 172350
rect 224702 172294 224798 172350
rect 224178 172226 224798 172294
rect 224178 172170 224274 172226
rect 224330 172170 224398 172226
rect 224454 172170 224522 172226
rect 224578 172170 224646 172226
rect 224702 172170 224798 172226
rect 224178 172102 224798 172170
rect 224178 172046 224274 172102
rect 224330 172046 224398 172102
rect 224454 172046 224522 172102
rect 224578 172046 224646 172102
rect 224702 172046 224798 172102
rect 224178 171978 224798 172046
rect 224178 171922 224274 171978
rect 224330 171922 224398 171978
rect 224454 171922 224522 171978
rect 224578 171922 224646 171978
rect 224702 171922 224798 171978
rect 224178 154350 224798 171922
rect 224178 154294 224274 154350
rect 224330 154294 224398 154350
rect 224454 154294 224522 154350
rect 224578 154294 224646 154350
rect 224702 154294 224798 154350
rect 224178 154226 224798 154294
rect 224178 154170 224274 154226
rect 224330 154170 224398 154226
rect 224454 154170 224522 154226
rect 224578 154170 224646 154226
rect 224702 154170 224798 154226
rect 224178 154102 224798 154170
rect 224178 154046 224274 154102
rect 224330 154046 224398 154102
rect 224454 154046 224522 154102
rect 224578 154046 224646 154102
rect 224702 154046 224798 154102
rect 224178 153978 224798 154046
rect 224178 153922 224274 153978
rect 224330 153922 224398 153978
rect 224454 153922 224522 153978
rect 224578 153922 224646 153978
rect 224702 153922 224798 153978
rect 224178 136350 224798 153922
rect 251178 166350 251798 183922
rect 251178 166294 251274 166350
rect 251330 166294 251398 166350
rect 251454 166294 251522 166350
rect 251578 166294 251646 166350
rect 251702 166294 251798 166350
rect 251178 166226 251798 166294
rect 251178 166170 251274 166226
rect 251330 166170 251398 166226
rect 251454 166170 251522 166226
rect 251578 166170 251646 166226
rect 251702 166170 251798 166226
rect 251178 166102 251798 166170
rect 251178 166046 251274 166102
rect 251330 166046 251398 166102
rect 251454 166046 251522 166102
rect 251578 166046 251646 166102
rect 251702 166046 251798 166102
rect 251178 165978 251798 166046
rect 251178 165922 251274 165978
rect 251330 165922 251398 165978
rect 251454 165922 251522 165978
rect 251578 165922 251646 165978
rect 251702 165922 251798 165978
rect 251178 148350 251798 165922
rect 251178 148294 251274 148350
rect 251330 148294 251398 148350
rect 251454 148294 251522 148350
rect 251578 148294 251646 148350
rect 251702 148294 251798 148350
rect 251178 148226 251798 148294
rect 251178 148170 251274 148226
rect 251330 148170 251398 148226
rect 251454 148170 251522 148226
rect 251578 148170 251646 148226
rect 251702 148170 251798 148226
rect 251178 148102 251798 148170
rect 251178 148046 251274 148102
rect 251330 148046 251398 148102
rect 251454 148046 251522 148102
rect 251578 148046 251646 148102
rect 251702 148046 251798 148102
rect 251178 147978 251798 148046
rect 251178 147922 251274 147978
rect 251330 147922 251398 147978
rect 251454 147922 251522 147978
rect 251578 147922 251646 147978
rect 251702 147922 251798 147978
rect 250236 139524 250292 139534
rect 224178 136294 224274 136350
rect 224330 136294 224398 136350
rect 224454 136294 224522 136350
rect 224578 136294 224646 136350
rect 224702 136294 224798 136350
rect 224178 136226 224798 136294
rect 224178 136170 224274 136226
rect 224330 136170 224398 136226
rect 224454 136170 224522 136226
rect 224578 136170 224646 136226
rect 224702 136170 224798 136226
rect 224178 136102 224798 136170
rect 224178 136046 224274 136102
rect 224330 136046 224398 136102
rect 224454 136046 224522 136102
rect 224578 136046 224646 136102
rect 224702 136046 224798 136102
rect 224178 135978 224798 136046
rect 224178 135922 224274 135978
rect 224330 135922 224398 135978
rect 224454 135922 224522 135978
rect 224578 135922 224646 135978
rect 224702 135922 224798 135978
rect 224178 118350 224798 135922
rect 225808 136350 226128 136384
rect 225808 136294 225878 136350
rect 225934 136294 226002 136350
rect 226058 136294 226128 136350
rect 225808 136226 226128 136294
rect 225808 136170 225878 136226
rect 225934 136170 226002 136226
rect 226058 136170 226128 136226
rect 225808 136102 226128 136170
rect 225808 136046 225878 136102
rect 225934 136046 226002 136102
rect 226058 136046 226128 136102
rect 225808 135978 226128 136046
rect 225808 135922 225878 135978
rect 225934 135922 226002 135978
rect 226058 135922 226128 135978
rect 225808 135888 226128 135922
rect 250236 134596 250292 139468
rect 250236 134530 250292 134540
rect 241168 130350 241488 130384
rect 241168 130294 241238 130350
rect 241294 130294 241362 130350
rect 241418 130294 241488 130350
rect 241168 130226 241488 130294
rect 241168 130170 241238 130226
rect 241294 130170 241362 130226
rect 241418 130170 241488 130226
rect 241168 130102 241488 130170
rect 241168 130046 241238 130102
rect 241294 130046 241362 130102
rect 241418 130046 241488 130102
rect 241168 129978 241488 130046
rect 241168 129922 241238 129978
rect 241294 129922 241362 129978
rect 241418 129922 241488 129978
rect 241168 129888 241488 129922
rect 251178 130350 251798 147922
rect 251178 130294 251274 130350
rect 251330 130294 251398 130350
rect 251454 130294 251522 130350
rect 251578 130294 251646 130350
rect 251702 130294 251798 130350
rect 251178 130226 251798 130294
rect 251178 130170 251274 130226
rect 251330 130170 251398 130226
rect 251454 130170 251522 130226
rect 251578 130170 251646 130226
rect 251702 130170 251798 130226
rect 251178 130102 251798 130170
rect 251178 130046 251274 130102
rect 251330 130046 251398 130102
rect 251454 130046 251522 130102
rect 251578 130046 251646 130102
rect 251702 130046 251798 130102
rect 251178 129978 251798 130046
rect 251178 129922 251274 129978
rect 251330 129922 251398 129978
rect 251454 129922 251522 129978
rect 251578 129922 251646 129978
rect 251702 129922 251798 129978
rect 224178 118294 224274 118350
rect 224330 118294 224398 118350
rect 224454 118294 224522 118350
rect 224578 118294 224646 118350
rect 224702 118294 224798 118350
rect 224178 118226 224798 118294
rect 224178 118170 224274 118226
rect 224330 118170 224398 118226
rect 224454 118170 224522 118226
rect 224578 118170 224646 118226
rect 224702 118170 224798 118226
rect 224178 118102 224798 118170
rect 224178 118046 224274 118102
rect 224330 118046 224398 118102
rect 224454 118046 224522 118102
rect 224578 118046 224646 118102
rect 224702 118046 224798 118102
rect 224178 117978 224798 118046
rect 224178 117922 224274 117978
rect 224330 117922 224398 117978
rect 224454 117922 224522 117978
rect 224578 117922 224646 117978
rect 224702 117922 224798 117978
rect 224178 100350 224798 117922
rect 225808 118350 226128 118384
rect 225808 118294 225878 118350
rect 225934 118294 226002 118350
rect 226058 118294 226128 118350
rect 225808 118226 226128 118294
rect 225808 118170 225878 118226
rect 225934 118170 226002 118226
rect 226058 118170 226128 118226
rect 225808 118102 226128 118170
rect 225808 118046 225878 118102
rect 225934 118046 226002 118102
rect 226058 118046 226128 118102
rect 225808 117978 226128 118046
rect 225808 117922 225878 117978
rect 225934 117922 226002 117978
rect 226058 117922 226128 117978
rect 225808 117888 226128 117922
rect 241168 112350 241488 112384
rect 241168 112294 241238 112350
rect 241294 112294 241362 112350
rect 241418 112294 241488 112350
rect 241168 112226 241488 112294
rect 241168 112170 241238 112226
rect 241294 112170 241362 112226
rect 241418 112170 241488 112226
rect 241168 112102 241488 112170
rect 241168 112046 241238 112102
rect 241294 112046 241362 112102
rect 241418 112046 241488 112102
rect 241168 111978 241488 112046
rect 241168 111922 241238 111978
rect 241294 111922 241362 111978
rect 241418 111922 241488 111978
rect 241168 111888 241488 111922
rect 251178 112350 251798 129922
rect 252812 179956 252868 179966
rect 252812 125300 252868 179900
rect 254898 172350 255518 189922
rect 257852 189812 257908 235340
rect 263900 235396 263956 238700
rect 272448 238350 272768 238384
rect 272448 238294 272518 238350
rect 272574 238294 272642 238350
rect 272698 238294 272768 238350
rect 272448 238226 272768 238294
rect 272448 238170 272518 238226
rect 272574 238170 272642 238226
rect 272698 238170 272768 238226
rect 272448 238102 272768 238170
rect 272448 238046 272518 238102
rect 272574 238046 272642 238102
rect 272698 238046 272768 238102
rect 272448 237978 272768 238046
rect 272448 237922 272518 237978
rect 272574 237922 272642 237978
rect 272698 237922 272768 237978
rect 272448 237888 272768 237922
rect 303168 238350 303488 238384
rect 303168 238294 303238 238350
rect 303294 238294 303362 238350
rect 303418 238294 303488 238350
rect 303168 238226 303488 238294
rect 303168 238170 303238 238226
rect 303294 238170 303362 238226
rect 303418 238170 303488 238226
rect 303168 238102 303488 238170
rect 303168 238046 303238 238102
rect 303294 238046 303362 238102
rect 303418 238046 303488 238102
rect 303168 237978 303488 238046
rect 303168 237922 303238 237978
rect 303294 237922 303362 237978
rect 303418 237922 303488 237978
rect 303168 237888 303488 237922
rect 263900 235330 263956 235340
rect 264908 235956 264964 235966
rect 262892 235172 262948 235182
rect 261212 234836 261268 234846
rect 257964 233492 258020 233502
rect 257964 194516 258020 233436
rect 261100 213220 261156 213230
rect 261100 212212 261156 213164
rect 261100 212146 261156 212156
rect 257964 194450 258020 194460
rect 258076 206276 258132 206286
rect 257852 189746 257908 189756
rect 258076 189140 258132 206220
rect 261212 205940 261268 234780
rect 261212 205874 261268 205884
rect 262108 206836 262164 206846
rect 262108 205858 262164 206780
rect 262108 205792 262164 205802
rect 262892 195188 262948 235116
rect 263900 225876 263956 225886
rect 263788 225316 263844 225326
rect 263788 224308 263844 225260
rect 263788 224242 263844 224252
rect 263900 222628 263956 225820
rect 263900 222562 263956 222572
rect 263788 220276 263844 220286
rect 263788 219268 263844 220220
rect 263788 219202 263844 219212
rect 263788 218596 263844 218606
rect 263788 217588 263844 218540
rect 263788 217522 263844 217532
rect 263788 216356 263844 216366
rect 263788 214228 263844 216300
rect 264908 215908 264964 235900
rect 287808 226350 288128 226384
rect 287808 226294 287878 226350
rect 287934 226294 288002 226350
rect 288058 226294 288128 226350
rect 287808 226226 288128 226294
rect 287808 226170 287878 226226
rect 287934 226170 288002 226226
rect 288058 226170 288128 226226
rect 287808 226102 288128 226170
rect 287808 226046 287878 226102
rect 287934 226046 288002 226102
rect 288058 226046 288128 226102
rect 287808 225978 288128 226046
rect 287808 225922 287878 225978
rect 287934 225922 288002 225978
rect 288058 225922 288128 225978
rect 287808 225888 288128 225922
rect 318528 226350 318848 226384
rect 318528 226294 318598 226350
rect 318654 226294 318722 226350
rect 318778 226294 318848 226350
rect 318528 226226 318848 226294
rect 318528 226170 318598 226226
rect 318654 226170 318722 226226
rect 318778 226170 318848 226226
rect 318528 226102 318848 226170
rect 318528 226046 318598 226102
rect 318654 226046 318722 226102
rect 318778 226046 318848 226102
rect 318528 225978 318848 226046
rect 318528 225922 318598 225978
rect 318654 225922 318722 225978
rect 318778 225922 318848 225978
rect 318528 225888 318848 225922
rect 272448 220350 272768 220384
rect 272448 220294 272518 220350
rect 272574 220294 272642 220350
rect 272698 220294 272768 220350
rect 272448 220226 272768 220294
rect 272448 220170 272518 220226
rect 272574 220170 272642 220226
rect 272698 220170 272768 220226
rect 272448 220102 272768 220170
rect 272448 220046 272518 220102
rect 272574 220046 272642 220102
rect 272698 220046 272768 220102
rect 272448 219978 272768 220046
rect 272448 219922 272518 219978
rect 272574 219922 272642 219978
rect 272698 219922 272768 219978
rect 272448 219888 272768 219922
rect 303168 220350 303488 220384
rect 303168 220294 303238 220350
rect 303294 220294 303362 220350
rect 303418 220294 303488 220350
rect 303168 220226 303488 220294
rect 303168 220170 303238 220226
rect 303294 220170 303362 220226
rect 303418 220170 303488 220226
rect 303168 220102 303488 220170
rect 303168 220046 303238 220102
rect 303294 220046 303362 220102
rect 303418 220046 303488 220102
rect 303168 219978 303488 220046
rect 303168 219922 303238 219978
rect 303294 219922 303362 219978
rect 303418 219922 303488 219978
rect 303168 219888 303488 219922
rect 264908 215842 264964 215852
rect 263788 214162 263844 214172
rect 263900 215796 263956 215806
rect 263788 213556 263844 213566
rect 263788 212100 263844 213500
rect 263900 213332 263956 215740
rect 263900 213266 263956 213276
rect 263788 212034 263844 212044
rect 263788 210420 263844 210430
rect 263788 209636 263844 210364
rect 263788 209570 263844 209580
rect 287808 208350 288128 208384
rect 287808 208294 287878 208350
rect 287934 208294 288002 208350
rect 288058 208294 288128 208350
rect 287808 208226 288128 208294
rect 287808 208170 287878 208226
rect 287934 208170 288002 208226
rect 288058 208170 288128 208226
rect 287808 208102 288128 208170
rect 287808 208046 287878 208102
rect 287934 208046 288002 208102
rect 288058 208046 288128 208102
rect 287808 207978 288128 208046
rect 287808 207922 287878 207978
rect 287934 207922 288002 207978
rect 288058 207922 288128 207978
rect 287808 207888 288128 207922
rect 318528 208350 318848 208384
rect 318528 208294 318598 208350
rect 318654 208294 318722 208350
rect 318778 208294 318848 208350
rect 318528 208226 318848 208294
rect 318528 208170 318598 208226
rect 318654 208170 318722 208226
rect 318778 208170 318848 208226
rect 318528 208102 318848 208170
rect 318528 208046 318598 208102
rect 318654 208046 318722 208102
rect 318778 208046 318848 208102
rect 318528 207978 318848 208046
rect 318528 207922 318598 207978
rect 318654 207922 318722 207978
rect 318778 207922 318848 207978
rect 318528 207888 318848 207922
rect 264796 205716 264852 205726
rect 264572 205156 264628 205166
rect 263788 198996 263844 199006
rect 263788 198298 263844 198940
rect 263788 198232 263844 198242
rect 263900 197876 263956 197886
rect 263788 197316 263844 197326
rect 263788 196858 263844 197260
rect 263788 196792 263844 196802
rect 263900 196678 263956 197820
rect 263900 196612 263956 196622
rect 262892 195122 262948 195132
rect 263788 196196 263844 196206
rect 263788 195058 263844 196140
rect 263788 194992 263844 195002
rect 264012 193396 264068 193406
rect 262108 193258 262164 193268
rect 258076 189074 258132 189084
rect 258412 191156 258468 191166
rect 258412 186238 258468 191100
rect 262108 190036 262164 193202
rect 263788 192178 263844 192188
rect 263788 191716 263844 192122
rect 263788 191650 263844 191660
rect 262108 189970 262164 189980
rect 263788 189658 263844 189668
rect 263788 189476 263844 189602
rect 263788 189410 263844 189420
rect 263900 189478 263956 189488
rect 263900 188356 263956 189422
rect 263900 188290 263956 188300
rect 263900 187498 263956 187508
rect 258636 186676 258692 186686
rect 258636 186418 258692 186620
rect 258636 186352 258692 186362
rect 258412 186172 258468 186182
rect 263788 186058 263844 186068
rect 263788 185556 263844 186002
rect 263788 185490 263844 185500
rect 263900 183876 263956 187442
rect 264012 187318 264068 193340
rect 264572 191268 264628 205100
rect 264796 193844 264852 205660
rect 272448 202350 272768 202384
rect 272448 202294 272518 202350
rect 272574 202294 272642 202350
rect 272698 202294 272768 202350
rect 272448 202226 272768 202294
rect 272448 202170 272518 202226
rect 272574 202170 272642 202226
rect 272698 202170 272768 202226
rect 272448 202102 272768 202170
rect 272448 202046 272518 202102
rect 272574 202046 272642 202102
rect 272698 202046 272768 202102
rect 272448 201978 272768 202046
rect 272448 201922 272518 201978
rect 272574 201922 272642 201978
rect 272698 201922 272768 201978
rect 272448 201888 272768 201922
rect 303168 202350 303488 202384
rect 303168 202294 303238 202350
rect 303294 202294 303362 202350
rect 303418 202294 303488 202350
rect 303168 202226 303488 202294
rect 303168 202170 303238 202226
rect 303294 202170 303362 202226
rect 303418 202170 303488 202226
rect 303168 202102 303488 202170
rect 303168 202046 303238 202102
rect 303294 202046 303362 202102
rect 303418 202046 303488 202102
rect 303168 201978 303488 202046
rect 303168 201922 303238 201978
rect 303294 201922 303362 201978
rect 303418 201922 303488 201978
rect 303168 201888 303488 201922
rect 264796 193778 264852 193788
rect 264572 191202 264628 191212
rect 287808 190350 288128 190384
rect 287808 190294 287878 190350
rect 287934 190294 288002 190350
rect 288058 190294 288128 190350
rect 287808 190226 288128 190294
rect 287808 190170 287878 190226
rect 287934 190170 288002 190226
rect 288058 190170 288128 190226
rect 287808 190102 288128 190170
rect 287808 190046 287878 190102
rect 287934 190046 288002 190102
rect 288058 190046 288128 190102
rect 287808 189978 288128 190046
rect 287808 189922 287878 189978
rect 287934 189922 288002 189978
rect 288058 189922 288128 189978
rect 287808 189888 288128 189922
rect 318528 190350 318848 190384
rect 318528 190294 318598 190350
rect 318654 190294 318722 190350
rect 318778 190294 318848 190350
rect 318528 190226 318848 190294
rect 318528 190170 318598 190226
rect 318654 190170 318722 190226
rect 318778 190170 318848 190226
rect 318528 190102 318848 190170
rect 318528 190046 318598 190102
rect 318654 190046 318722 190102
rect 318778 190046 318848 190102
rect 318528 189978 318848 190046
rect 318528 189922 318598 189978
rect 318654 189922 318722 189978
rect 318778 189922 318848 189978
rect 318528 189888 318848 189922
rect 264012 187252 264068 187262
rect 272448 184350 272768 184384
rect 272448 184294 272518 184350
rect 272574 184294 272642 184350
rect 272698 184294 272768 184350
rect 272448 184226 272768 184294
rect 272448 184170 272518 184226
rect 272574 184170 272642 184226
rect 272698 184170 272768 184226
rect 272448 184102 272768 184170
rect 272448 184046 272518 184102
rect 272574 184046 272642 184102
rect 272698 184046 272768 184102
rect 272448 183978 272768 184046
rect 272448 183922 272518 183978
rect 272574 183922 272642 183978
rect 272698 183922 272768 183978
rect 272448 183888 272768 183922
rect 303168 184350 303488 184384
rect 303168 184294 303238 184350
rect 303294 184294 303362 184350
rect 303418 184294 303488 184350
rect 303168 184226 303488 184294
rect 303168 184170 303238 184226
rect 303294 184170 303362 184226
rect 303418 184170 303488 184226
rect 303168 184102 303488 184170
rect 303168 184046 303238 184102
rect 303294 184046 303362 184102
rect 303418 184046 303488 184102
rect 303168 183978 303488 184046
rect 303168 183922 303238 183978
rect 303294 183922 303362 183978
rect 303418 183922 303488 183978
rect 303168 183888 303488 183922
rect 263900 183810 263956 183820
rect 261436 182196 261492 182206
rect 257852 178836 257908 178846
rect 254898 172294 254994 172350
rect 255050 172294 255118 172350
rect 255174 172294 255242 172350
rect 255298 172294 255366 172350
rect 255422 172294 255518 172350
rect 254898 172226 255518 172294
rect 254898 172170 254994 172226
rect 255050 172170 255118 172226
rect 255174 172170 255242 172226
rect 255298 172170 255366 172226
rect 255422 172170 255518 172226
rect 254898 172102 255518 172170
rect 254898 172046 254994 172102
rect 255050 172046 255118 172102
rect 255174 172046 255242 172102
rect 255298 172046 255366 172102
rect 255422 172046 255518 172102
rect 254898 171978 255518 172046
rect 254898 171922 254994 171978
rect 255050 171922 255118 171978
rect 255174 171922 255242 171978
rect 255298 171922 255366 171978
rect 255422 171922 255518 171978
rect 254898 154350 255518 171922
rect 254898 154294 254994 154350
rect 255050 154294 255118 154350
rect 255174 154294 255242 154350
rect 255298 154294 255366 154350
rect 255422 154294 255518 154350
rect 254898 154226 255518 154294
rect 254898 154170 254994 154226
rect 255050 154170 255118 154226
rect 255174 154170 255242 154226
rect 255298 154170 255366 154226
rect 255422 154170 255518 154226
rect 254898 154102 255518 154170
rect 254898 154046 254994 154102
rect 255050 154046 255118 154102
rect 255174 154046 255242 154102
rect 255298 154046 255366 154102
rect 255422 154046 255518 154102
rect 254898 153978 255518 154046
rect 254898 153922 254994 153978
rect 255050 153922 255118 153978
rect 255174 153922 255242 153978
rect 255298 153922 255366 153978
rect 255422 153922 255518 153978
rect 254898 136350 255518 153922
rect 256396 178276 256452 178286
rect 256172 142100 256228 142110
rect 256172 141764 256228 142044
rect 256172 141698 256228 141708
rect 254898 136294 254994 136350
rect 255050 136294 255118 136350
rect 255174 136294 255242 136350
rect 255298 136294 255366 136350
rect 255422 136294 255518 136350
rect 254898 136226 255518 136294
rect 254898 136170 254994 136226
rect 255050 136170 255118 136226
rect 255174 136170 255242 136226
rect 255298 136170 255366 136226
rect 255422 136170 255518 136226
rect 254898 136102 255518 136170
rect 254898 136046 254994 136102
rect 255050 136046 255118 136102
rect 255174 136046 255242 136102
rect 255298 136046 255366 136102
rect 255422 136046 255518 136102
rect 254898 135978 255518 136046
rect 254898 135922 254994 135978
rect 255050 135922 255118 135978
rect 255174 135922 255242 135978
rect 255298 135922 255366 135978
rect 255422 135922 255518 135978
rect 252812 125234 252868 125244
rect 252924 128548 252980 128558
rect 251178 112294 251274 112350
rect 251330 112294 251398 112350
rect 251454 112294 251522 112350
rect 251578 112294 251646 112350
rect 251702 112294 251798 112350
rect 251178 112226 251798 112294
rect 251178 112170 251274 112226
rect 251330 112170 251398 112226
rect 251454 112170 251522 112226
rect 251578 112170 251646 112226
rect 251702 112170 251798 112226
rect 251178 112102 251798 112170
rect 251178 112046 251274 112102
rect 251330 112046 251398 112102
rect 251454 112046 251522 112102
rect 251578 112046 251646 112102
rect 251702 112046 251798 112102
rect 251178 111978 251798 112046
rect 251178 111922 251274 111978
rect 251330 111922 251398 111978
rect 251454 111922 251522 111978
rect 251578 111922 251646 111978
rect 251702 111922 251798 111978
rect 249452 109956 249508 109966
rect 230188 101780 230244 101790
rect 230188 100772 230244 101724
rect 230188 100706 230244 100716
rect 224178 100294 224274 100350
rect 224330 100294 224398 100350
rect 224454 100294 224522 100350
rect 224578 100294 224646 100350
rect 224702 100294 224798 100350
rect 224178 100226 224798 100294
rect 224178 100170 224274 100226
rect 224330 100170 224398 100226
rect 224454 100170 224522 100226
rect 224578 100170 224646 100226
rect 224702 100170 224798 100226
rect 224178 100102 224798 100170
rect 224178 100046 224274 100102
rect 224330 100046 224398 100102
rect 224454 100046 224522 100102
rect 224578 100046 224646 100102
rect 224702 100046 224798 100102
rect 224178 99978 224798 100046
rect 224178 99922 224274 99978
rect 224330 99922 224398 99978
rect 224454 99922 224522 99978
rect 224578 99922 224646 99978
rect 224702 99922 224798 99978
rect 224178 82350 224798 99922
rect 230188 92596 230244 92606
rect 230188 90244 230244 92540
rect 230188 90178 230244 90188
rect 224178 82294 224274 82350
rect 224330 82294 224398 82350
rect 224454 82294 224522 82350
rect 224578 82294 224646 82350
rect 224702 82294 224798 82350
rect 224178 82226 224798 82294
rect 224178 82170 224274 82226
rect 224330 82170 224398 82226
rect 224454 82170 224522 82226
rect 224578 82170 224646 82226
rect 224702 82170 224798 82226
rect 224178 82102 224798 82170
rect 224178 82046 224274 82102
rect 224330 82046 224398 82102
rect 224454 82046 224522 82102
rect 224578 82046 224646 82102
rect 224702 82046 224798 82102
rect 224178 81978 224798 82046
rect 224178 81922 224274 81978
rect 224330 81922 224398 81978
rect 224454 81922 224522 81978
rect 224578 81922 224646 81978
rect 224702 81922 224798 81978
rect 224178 64350 224798 81922
rect 249452 71540 249508 109900
rect 249452 71474 249508 71484
rect 251178 94350 251798 111922
rect 251178 94294 251274 94350
rect 251330 94294 251398 94350
rect 251454 94294 251522 94350
rect 251578 94294 251646 94350
rect 251702 94294 251798 94350
rect 251178 94226 251798 94294
rect 251178 94170 251274 94226
rect 251330 94170 251398 94226
rect 251454 94170 251522 94226
rect 251578 94170 251646 94226
rect 251702 94170 251798 94226
rect 251178 94102 251798 94170
rect 251178 94046 251274 94102
rect 251330 94046 251398 94102
rect 251454 94046 251522 94102
rect 251578 94046 251646 94102
rect 251702 94046 251798 94102
rect 251178 93978 251798 94046
rect 251178 93922 251274 93978
rect 251330 93922 251398 93978
rect 251454 93922 251522 93978
rect 251578 93922 251646 93978
rect 251702 93922 251798 93978
rect 251178 76350 251798 93922
rect 251178 76294 251274 76350
rect 251330 76294 251398 76350
rect 251454 76294 251522 76350
rect 251578 76294 251646 76350
rect 251702 76294 251798 76350
rect 251178 76226 251798 76294
rect 251178 76170 251274 76226
rect 251330 76170 251398 76226
rect 251454 76170 251522 76226
rect 251578 76170 251646 76226
rect 251702 76170 251798 76226
rect 251178 76102 251798 76170
rect 251178 76046 251274 76102
rect 251330 76046 251398 76102
rect 251454 76046 251522 76102
rect 251578 76046 251646 76102
rect 251702 76046 251798 76102
rect 251178 75978 251798 76046
rect 251178 75922 251274 75978
rect 251330 75922 251398 75978
rect 251454 75922 251522 75978
rect 251578 75922 251646 75978
rect 251702 75922 251798 75978
rect 224178 64294 224274 64350
rect 224330 64294 224398 64350
rect 224454 64294 224522 64350
rect 224578 64294 224646 64350
rect 224702 64294 224798 64350
rect 224178 64226 224798 64294
rect 224178 64170 224274 64226
rect 224330 64170 224398 64226
rect 224454 64170 224522 64226
rect 224578 64170 224646 64226
rect 224702 64170 224798 64226
rect 224178 64102 224798 64170
rect 224178 64046 224274 64102
rect 224330 64046 224398 64102
rect 224454 64046 224522 64102
rect 224578 64046 224646 64102
rect 224702 64046 224798 64102
rect 224178 63978 224798 64046
rect 224178 63922 224274 63978
rect 224330 63922 224398 63978
rect 224454 63922 224522 63978
rect 224578 63922 224646 63978
rect 224702 63922 224798 63978
rect 224178 46350 224798 63922
rect 225808 64350 226128 64384
rect 225808 64294 225878 64350
rect 225934 64294 226002 64350
rect 226058 64294 226128 64350
rect 225808 64226 226128 64294
rect 225808 64170 225878 64226
rect 225934 64170 226002 64226
rect 226058 64170 226128 64226
rect 225808 64102 226128 64170
rect 225808 64046 225878 64102
rect 225934 64046 226002 64102
rect 226058 64046 226128 64102
rect 225808 63978 226128 64046
rect 225808 63922 225878 63978
rect 225934 63922 226002 63978
rect 226058 63922 226128 63978
rect 225808 63888 226128 63922
rect 241168 58350 241488 58384
rect 241168 58294 241238 58350
rect 241294 58294 241362 58350
rect 241418 58294 241488 58350
rect 241168 58226 241488 58294
rect 241168 58170 241238 58226
rect 241294 58170 241362 58226
rect 241418 58170 241488 58226
rect 241168 58102 241488 58170
rect 241168 58046 241238 58102
rect 241294 58046 241362 58102
rect 241418 58046 241488 58102
rect 241168 57978 241488 58046
rect 241168 57922 241238 57978
rect 241294 57922 241362 57978
rect 241418 57922 241488 57978
rect 241168 57888 241488 57922
rect 251178 58350 251798 75922
rect 251178 58294 251274 58350
rect 251330 58294 251398 58350
rect 251454 58294 251522 58350
rect 251578 58294 251646 58350
rect 251702 58294 251798 58350
rect 251178 58226 251798 58294
rect 251178 58170 251274 58226
rect 251330 58170 251398 58226
rect 251454 58170 251522 58226
rect 251578 58170 251646 58226
rect 251702 58170 251798 58226
rect 251178 58102 251798 58170
rect 251178 58046 251274 58102
rect 251330 58046 251398 58102
rect 251454 58046 251522 58102
rect 251578 58046 251646 58102
rect 251702 58046 251798 58102
rect 251178 57978 251798 58046
rect 251178 57922 251274 57978
rect 251330 57922 251398 57978
rect 251454 57922 251522 57978
rect 251578 57922 251646 57978
rect 251702 57922 251798 57978
rect 224178 46294 224274 46350
rect 224330 46294 224398 46350
rect 224454 46294 224522 46350
rect 224578 46294 224646 46350
rect 224702 46294 224798 46350
rect 224178 46226 224798 46294
rect 224178 46170 224274 46226
rect 224330 46170 224398 46226
rect 224454 46170 224522 46226
rect 224578 46170 224646 46226
rect 224702 46170 224798 46226
rect 224178 46102 224798 46170
rect 224178 46046 224274 46102
rect 224330 46046 224398 46102
rect 224454 46046 224522 46102
rect 224578 46046 224646 46102
rect 224702 46046 224798 46102
rect 224178 45978 224798 46046
rect 224178 45922 224274 45978
rect 224330 45922 224398 45978
rect 224454 45922 224522 45978
rect 224578 45922 224646 45978
rect 224702 45922 224798 45978
rect 224178 28350 224798 45922
rect 225808 46350 226128 46384
rect 225808 46294 225878 46350
rect 225934 46294 226002 46350
rect 226058 46294 226128 46350
rect 225808 46226 226128 46294
rect 225808 46170 225878 46226
rect 225934 46170 226002 46226
rect 226058 46170 226128 46226
rect 225808 46102 226128 46170
rect 225808 46046 225878 46102
rect 225934 46046 226002 46102
rect 226058 46046 226128 46102
rect 225808 45978 226128 46046
rect 225808 45922 225878 45978
rect 225934 45922 226002 45978
rect 226058 45922 226128 45978
rect 225808 45888 226128 45922
rect 241168 40350 241488 40384
rect 241168 40294 241238 40350
rect 241294 40294 241362 40350
rect 241418 40294 241488 40350
rect 241168 40226 241488 40294
rect 241168 40170 241238 40226
rect 241294 40170 241362 40226
rect 241418 40170 241488 40226
rect 241168 40102 241488 40170
rect 241168 40046 241238 40102
rect 241294 40046 241362 40102
rect 241418 40046 241488 40102
rect 241168 39978 241488 40046
rect 241168 39922 241238 39978
rect 241294 39922 241362 39978
rect 241418 39922 241488 39978
rect 241168 39888 241488 39922
rect 251178 40350 251798 57922
rect 251916 122836 251972 122846
rect 251916 49476 251972 122780
rect 252812 120596 252868 120606
rect 252812 69972 252868 120540
rect 252924 117908 252980 128492
rect 252924 117842 252980 117852
rect 254492 120036 254548 120046
rect 254492 78372 254548 119980
rect 254492 78306 254548 78316
rect 254898 118350 255518 135922
rect 256396 121940 256452 178220
rect 257852 126644 257908 178780
rect 261324 150836 261380 150846
rect 259980 150276 260036 150286
rect 257852 126578 257908 126588
rect 259756 149716 259812 149726
rect 256396 121874 256452 121884
rect 259532 121716 259588 121726
rect 254898 118294 254994 118350
rect 255050 118294 255118 118350
rect 255174 118294 255242 118350
rect 255298 118294 255366 118350
rect 255422 118294 255518 118350
rect 254898 118226 255518 118294
rect 254898 118170 254994 118226
rect 255050 118170 255118 118226
rect 255174 118170 255242 118226
rect 255298 118170 255366 118226
rect 255422 118170 255518 118226
rect 254898 118102 255518 118170
rect 254898 118046 254994 118102
rect 255050 118046 255118 118102
rect 255174 118046 255242 118102
rect 255298 118046 255366 118102
rect 255422 118046 255518 118102
rect 254898 117978 255518 118046
rect 254898 117922 254994 117978
rect 255050 117922 255118 117978
rect 255174 117922 255242 117978
rect 255298 117922 255366 117978
rect 255422 117922 255518 117978
rect 254898 100350 255518 117922
rect 254898 100294 254994 100350
rect 255050 100294 255118 100350
rect 255174 100294 255242 100350
rect 255298 100294 255366 100350
rect 255422 100294 255518 100350
rect 254898 100226 255518 100294
rect 254898 100170 254994 100226
rect 255050 100170 255118 100226
rect 255174 100170 255242 100226
rect 255298 100170 255366 100226
rect 255422 100170 255518 100226
rect 254898 100102 255518 100170
rect 254898 100046 254994 100102
rect 255050 100046 255118 100102
rect 255174 100046 255242 100102
rect 255298 100046 255366 100102
rect 255422 100046 255518 100102
rect 254898 99978 255518 100046
rect 254898 99922 254994 99978
rect 255050 99922 255118 99978
rect 255174 99922 255242 99978
rect 255298 99922 255366 99978
rect 255422 99922 255518 99978
rect 254898 82350 255518 99922
rect 254898 82294 254994 82350
rect 255050 82294 255118 82350
rect 255174 82294 255242 82350
rect 255298 82294 255366 82350
rect 255422 82294 255518 82350
rect 254898 82226 255518 82294
rect 254898 82170 254994 82226
rect 255050 82170 255118 82226
rect 255174 82170 255242 82226
rect 255298 82170 255366 82226
rect 255422 82170 255518 82226
rect 254898 82102 255518 82170
rect 254898 82046 254994 82102
rect 255050 82046 255118 82102
rect 255174 82046 255242 82102
rect 255298 82046 255366 82102
rect 255422 82046 255518 82102
rect 254898 81978 255518 82046
rect 254898 81922 254994 81978
rect 255050 81922 255118 81978
rect 255174 81922 255242 81978
rect 255298 81922 255366 81978
rect 255422 81922 255518 81978
rect 252812 69906 252868 69916
rect 252924 74788 252980 74798
rect 252812 68068 252868 68078
rect 252812 67844 252868 68012
rect 252812 67778 252868 67788
rect 251916 49410 251972 49420
rect 252924 45444 252980 74732
rect 252924 45378 252980 45388
rect 254898 64350 255518 81922
rect 254898 64294 254994 64350
rect 255050 64294 255118 64350
rect 255174 64294 255242 64350
rect 255298 64294 255366 64350
rect 255422 64294 255518 64350
rect 254898 64226 255518 64294
rect 254898 64170 254994 64226
rect 255050 64170 255118 64226
rect 255174 64170 255242 64226
rect 255298 64170 255366 64226
rect 255422 64170 255518 64226
rect 254898 64102 255518 64170
rect 254898 64046 254994 64102
rect 255050 64046 255118 64102
rect 255174 64046 255242 64102
rect 255298 64046 255366 64102
rect 255422 64046 255518 64102
rect 254898 63978 255518 64046
rect 254898 63922 254994 63978
rect 255050 63922 255118 63978
rect 255174 63922 255242 63978
rect 255298 63922 255366 63978
rect 255422 63922 255518 63978
rect 254898 46350 255518 63922
rect 256172 121156 256228 121166
rect 256172 53508 256228 121100
rect 257852 118356 257908 118366
rect 257852 73332 257908 118300
rect 258076 113316 258132 113326
rect 257852 73266 257908 73276
rect 257964 85764 258020 85774
rect 256172 53442 256228 53452
rect 257964 50148 258020 85708
rect 258076 73220 258132 113260
rect 258076 73154 258132 73164
rect 258188 77364 258244 77374
rect 257964 50082 258020 50092
rect 258188 47460 258244 77308
rect 259532 52836 259588 121660
rect 259756 121268 259812 149660
rect 259980 122612 260036 150220
rect 259980 122546 260036 122556
rect 261212 146916 261268 146926
rect 259756 121202 259812 121212
rect 259980 120932 260036 120942
rect 259980 117478 260036 120876
rect 261212 119924 261268 146860
rect 261324 125972 261380 150780
rect 261324 125906 261380 125916
rect 261212 119858 261268 119868
rect 259980 117412 260036 117422
rect 261436 117348 261492 182140
rect 264572 181636 264628 181646
rect 261436 117282 261492 117292
rect 262892 179396 262948 179406
rect 259644 116116 259700 116126
rect 259644 71428 259700 116060
rect 262892 114548 262948 179340
rect 263788 176036 263844 176046
rect 263788 174020 263844 175980
rect 263788 173954 263844 173964
rect 263900 168756 263956 168766
rect 263788 168196 263844 168206
rect 263788 163828 263844 168140
rect 263788 163762 263844 163772
rect 263900 162148 263956 168700
rect 263900 162082 263956 162092
rect 263788 151396 263844 151406
rect 263788 150500 263844 151340
rect 263788 150434 263844 150444
rect 264012 139860 264068 139870
rect 263900 139748 263956 139758
rect 263788 137956 263844 137966
rect 263788 137818 263844 137900
rect 263788 137752 263844 137762
rect 263900 136836 263956 139692
rect 263900 136770 263956 136780
rect 264012 136276 264068 139804
rect 264012 136210 264068 136220
rect 263900 134036 263956 134046
rect 263788 133476 263844 133486
rect 263788 132958 263844 133420
rect 263788 132892 263844 132902
rect 263900 132778 263956 133980
rect 263900 132712 263956 132722
rect 263900 131338 263956 131348
rect 263788 130116 263844 130126
rect 263788 128638 263844 130060
rect 263900 129556 263956 131282
rect 263900 129490 263956 129500
rect 263788 128572 263844 128582
rect 263900 128996 263956 129006
rect 263788 128436 263844 128446
rect 263788 127198 263844 128380
rect 263900 127918 263956 128940
rect 264572 128548 264628 181580
rect 264684 177716 264740 177726
rect 264684 172228 264740 177660
rect 264684 172162 264740 172172
rect 287808 172350 288128 172384
rect 287808 172294 287878 172350
rect 287934 172294 288002 172350
rect 288058 172294 288128 172350
rect 287808 172226 288128 172294
rect 287808 172170 287878 172226
rect 287934 172170 288002 172226
rect 288058 172170 288128 172226
rect 287808 172102 288128 172170
rect 287808 172046 287878 172102
rect 287934 172046 288002 172102
rect 288058 172046 288128 172102
rect 287808 171978 288128 172046
rect 287808 171922 287878 171978
rect 287934 171922 288002 171978
rect 288058 171922 288128 171978
rect 287808 171888 288128 171922
rect 318528 172350 318848 172384
rect 318528 172294 318598 172350
rect 318654 172294 318722 172350
rect 318778 172294 318848 172350
rect 318528 172226 318848 172294
rect 318528 172170 318598 172226
rect 318654 172170 318722 172226
rect 318778 172170 318848 172226
rect 318528 172102 318848 172170
rect 318528 172046 318598 172102
rect 318654 172046 318722 172102
rect 318778 172046 318848 172102
rect 318528 171978 318848 172046
rect 318528 171922 318598 171978
rect 318654 171922 318722 171978
rect 318778 171922 318848 171978
rect 318528 171888 318848 171922
rect 272448 166350 272768 166384
rect 272448 166294 272518 166350
rect 272574 166294 272642 166350
rect 272698 166294 272768 166350
rect 272448 166226 272768 166294
rect 272448 166170 272518 166226
rect 272574 166170 272642 166226
rect 272698 166170 272768 166226
rect 272448 166102 272768 166170
rect 272448 166046 272518 166102
rect 272574 166046 272642 166102
rect 272698 166046 272768 166102
rect 272448 165978 272768 166046
rect 272448 165922 272518 165978
rect 272574 165922 272642 165978
rect 272698 165922 272768 165978
rect 272448 165888 272768 165922
rect 303168 166350 303488 166384
rect 303168 166294 303238 166350
rect 303294 166294 303362 166350
rect 303418 166294 303488 166350
rect 303168 166226 303488 166294
rect 303168 166170 303238 166226
rect 303294 166170 303362 166226
rect 303418 166170 303488 166226
rect 303168 166102 303488 166170
rect 303168 166046 303238 166102
rect 303294 166046 303362 166102
rect 303418 166046 303488 166102
rect 303168 165978 303488 166046
rect 303168 165922 303238 165978
rect 303294 165922 303362 165978
rect 303418 165922 303488 165978
rect 303168 165888 303488 165922
rect 287808 154350 288128 154384
rect 287808 154294 287878 154350
rect 287934 154294 288002 154350
rect 288058 154294 288128 154350
rect 287808 154226 288128 154294
rect 287808 154170 287878 154226
rect 287934 154170 288002 154226
rect 288058 154170 288128 154226
rect 287808 154102 288128 154170
rect 287808 154046 287878 154102
rect 287934 154046 288002 154102
rect 288058 154046 288128 154102
rect 287808 153978 288128 154046
rect 287808 153922 287878 153978
rect 287934 153922 288002 153978
rect 288058 153922 288128 153978
rect 287808 153888 288128 153922
rect 318528 154350 318848 154384
rect 318528 154294 318598 154350
rect 318654 154294 318722 154350
rect 318778 154294 318848 154350
rect 318528 154226 318848 154294
rect 318528 154170 318598 154226
rect 318654 154170 318722 154226
rect 318778 154170 318848 154226
rect 318528 154102 318848 154170
rect 318528 154046 318598 154102
rect 318654 154046 318722 154102
rect 318778 154046 318848 154102
rect 318528 153978 318848 154046
rect 318528 153922 318598 153978
rect 318654 153922 318722 153978
rect 318778 153922 318848 153978
rect 318528 153888 318848 153922
rect 264684 153076 264740 153086
rect 264684 147028 264740 153020
rect 272448 148350 272768 148384
rect 272448 148294 272518 148350
rect 272574 148294 272642 148350
rect 272698 148294 272768 148350
rect 272448 148226 272768 148294
rect 272448 148170 272518 148226
rect 272574 148170 272642 148226
rect 272698 148170 272768 148226
rect 272448 148102 272768 148170
rect 272448 148046 272518 148102
rect 272574 148046 272642 148102
rect 272698 148046 272768 148102
rect 272448 147978 272768 148046
rect 272448 147922 272518 147978
rect 272574 147922 272642 147978
rect 272698 147922 272768 147978
rect 272448 147888 272768 147922
rect 303168 148350 303488 148384
rect 303168 148294 303238 148350
rect 303294 148294 303362 148350
rect 303418 148294 303488 148350
rect 303168 148226 303488 148294
rect 303168 148170 303238 148226
rect 303294 148170 303362 148226
rect 303418 148170 303488 148226
rect 303168 148102 303488 148170
rect 303168 148046 303238 148102
rect 303294 148046 303362 148102
rect 303418 148046 303488 148102
rect 303168 147978 303488 148046
rect 303168 147922 303238 147978
rect 303294 147922 303362 147978
rect 303418 147922 303488 147978
rect 303168 147888 303488 147922
rect 264684 146962 264740 146972
rect 287808 136350 288128 136384
rect 287808 136294 287878 136350
rect 287934 136294 288002 136350
rect 288058 136294 288128 136350
rect 287808 136226 288128 136294
rect 287808 136170 287878 136226
rect 287934 136170 288002 136226
rect 288058 136170 288128 136226
rect 287808 136102 288128 136170
rect 287808 136046 287878 136102
rect 287934 136046 288002 136102
rect 288058 136046 288128 136102
rect 287808 135978 288128 136046
rect 287808 135922 287878 135978
rect 287934 135922 288002 135978
rect 288058 135922 288128 135978
rect 287808 135888 288128 135922
rect 318528 136350 318848 136384
rect 318528 136294 318598 136350
rect 318654 136294 318722 136350
rect 318778 136294 318848 136350
rect 318528 136226 318848 136294
rect 318528 136170 318598 136226
rect 318654 136170 318722 136226
rect 318778 136170 318848 136226
rect 318528 136102 318848 136170
rect 318528 136046 318598 136102
rect 318654 136046 318722 136102
rect 318778 136046 318848 136102
rect 318528 135978 318848 136046
rect 318528 135922 318598 135978
rect 318654 135922 318722 135978
rect 318778 135922 318848 135978
rect 318528 135888 318848 135922
rect 264796 131158 264852 131168
rect 264572 128482 264628 128492
rect 264684 130676 264740 130686
rect 263900 127852 263956 127862
rect 264012 127876 264068 127886
rect 263788 127142 263956 127198
rect 263788 126756 263844 126766
rect 263788 126118 263844 126700
rect 263788 126052 263844 126062
rect 263900 125218 263956 127142
rect 263900 125152 263956 125162
rect 264012 121798 264068 127820
rect 264012 121732 264068 121742
rect 264684 120932 264740 130620
rect 264796 124516 264852 131102
rect 272448 130350 272768 130384
rect 272448 130294 272518 130350
rect 272574 130294 272642 130350
rect 272698 130294 272768 130350
rect 272448 130226 272768 130294
rect 272448 130170 272518 130226
rect 272574 130170 272642 130226
rect 272698 130170 272768 130226
rect 272448 130102 272768 130170
rect 272448 130046 272518 130102
rect 272574 130046 272642 130102
rect 272698 130046 272768 130102
rect 272448 129978 272768 130046
rect 272448 129922 272518 129978
rect 272574 129922 272642 129978
rect 272698 129922 272768 129978
rect 272448 129888 272768 129922
rect 303168 130350 303488 130384
rect 303168 130294 303238 130350
rect 303294 130294 303362 130350
rect 303418 130294 303488 130350
rect 303168 130226 303488 130294
rect 303168 130170 303238 130226
rect 303294 130170 303362 130226
rect 303418 130170 303488 130226
rect 303168 130102 303488 130170
rect 303168 130046 303238 130102
rect 303294 130046 303362 130102
rect 303418 130046 303488 130102
rect 303168 129978 303488 130046
rect 303168 129922 303238 129978
rect 303294 129922 303362 129978
rect 303418 129922 303488 129978
rect 303168 129888 303488 129922
rect 264796 124450 264852 124460
rect 264684 120866 264740 120876
rect 287808 118350 288128 118384
rect 287808 118294 287878 118350
rect 287934 118294 288002 118350
rect 288058 118294 288128 118350
rect 287808 118226 288128 118294
rect 287808 118170 287878 118226
rect 287934 118170 288002 118226
rect 288058 118170 288128 118226
rect 287808 118102 288128 118170
rect 287808 118046 287878 118102
rect 287934 118046 288002 118102
rect 288058 118046 288128 118102
rect 287808 117978 288128 118046
rect 287808 117922 287878 117978
rect 287934 117922 288002 117978
rect 288058 117922 288128 117978
rect 287808 117888 288128 117922
rect 318528 118350 318848 118384
rect 318528 118294 318598 118350
rect 318654 118294 318722 118350
rect 318778 118294 318848 118350
rect 318528 118226 318848 118294
rect 318528 118170 318598 118226
rect 318654 118170 318722 118226
rect 318778 118170 318848 118226
rect 318528 118102 318848 118170
rect 318528 118046 318598 118102
rect 318654 118046 318722 118102
rect 318778 118046 318848 118102
rect 318528 117978 318848 118046
rect 318528 117922 318598 117978
rect 318654 117922 318722 117978
rect 318778 117922 318848 117978
rect 318528 117888 318848 117922
rect 262892 114482 262948 114492
rect 261436 114436 261492 114446
rect 259756 107156 259812 107166
rect 259756 84868 259812 107100
rect 261324 106036 261380 106046
rect 259756 84802 259812 84812
rect 261212 92036 261268 92046
rect 259644 71362 259700 71372
rect 259532 52770 259588 52780
rect 261212 52164 261268 91980
rect 261324 69748 261380 105980
rect 261436 91924 261492 114380
rect 261436 91858 261492 91868
rect 262892 113876 262948 113886
rect 262892 69860 262948 113820
rect 272448 112350 272768 112384
rect 272448 112294 272518 112350
rect 272574 112294 272642 112350
rect 272698 112294 272768 112350
rect 272448 112226 272768 112294
rect 272448 112170 272518 112226
rect 272574 112170 272642 112226
rect 272698 112170 272768 112226
rect 272448 112102 272768 112170
rect 272448 112046 272518 112102
rect 272574 112046 272642 112102
rect 272698 112046 272768 112102
rect 272448 111978 272768 112046
rect 272448 111922 272518 111978
rect 272574 111922 272642 111978
rect 272698 111922 272768 111978
rect 272448 111888 272768 111922
rect 303168 112350 303488 112384
rect 303168 112294 303238 112350
rect 303294 112294 303362 112350
rect 303418 112294 303488 112350
rect 303168 112226 303488 112294
rect 303168 112170 303238 112226
rect 303294 112170 303362 112226
rect 303418 112170 303488 112226
rect 303168 112102 303488 112170
rect 303168 112046 303238 112102
rect 303294 112046 303362 112102
rect 303418 112046 303488 112102
rect 303168 111978 303488 112046
rect 303168 111922 303238 111978
rect 303294 111922 303362 111978
rect 303418 111922 303488 111978
rect 303168 111888 303488 111922
rect 264684 111636 264740 111646
rect 264124 109396 264180 109406
rect 263788 104916 263844 104926
rect 263788 103348 263844 104860
rect 263788 103282 263844 103292
rect 263900 104356 263956 104366
rect 263900 101668 263956 104300
rect 263900 101602 263956 101612
rect 264012 103796 264068 103806
rect 264012 99988 264068 103740
rect 264124 103124 264180 109340
rect 264124 103058 264180 103068
rect 264572 103236 264628 103246
rect 264012 99922 264068 99932
rect 263788 98756 263844 98766
rect 263788 91700 263844 98700
rect 263788 91634 263844 91644
rect 263788 91476 263844 91486
rect 263788 85764 263844 91420
rect 264572 88340 264628 103180
rect 264684 96740 264740 111580
rect 265132 108836 265188 108846
rect 265020 99876 265076 99886
rect 264684 96674 264740 96684
rect 264796 99316 264852 99326
rect 264572 88274 264628 88284
rect 263788 85698 263844 85708
rect 264572 86996 264628 87006
rect 263788 80836 263844 80846
rect 263788 78260 263844 80780
rect 263788 78194 263844 78204
rect 263788 75796 263844 75806
rect 263788 73108 263844 75740
rect 264572 74788 264628 86940
rect 264796 86548 264852 99260
rect 265020 89908 265076 99820
rect 265132 98308 265188 108780
rect 287808 100350 288128 100384
rect 287808 100294 287878 100350
rect 287934 100294 288002 100350
rect 288058 100294 288128 100350
rect 287808 100226 288128 100294
rect 287808 100170 287878 100226
rect 287934 100170 288002 100226
rect 288058 100170 288128 100226
rect 287808 100102 288128 100170
rect 287808 100046 287878 100102
rect 287934 100046 288002 100102
rect 288058 100046 288128 100102
rect 287808 99978 288128 100046
rect 287808 99922 287878 99978
rect 287934 99922 288002 99978
rect 288058 99922 288128 99978
rect 287808 99888 288128 99922
rect 318528 100350 318848 100384
rect 318528 100294 318598 100350
rect 318654 100294 318722 100350
rect 318778 100294 318848 100350
rect 318528 100226 318848 100294
rect 318528 100170 318598 100226
rect 318654 100170 318722 100226
rect 318778 100170 318848 100226
rect 318528 100102 318848 100170
rect 318528 100046 318598 100102
rect 318654 100046 318722 100102
rect 318778 100046 318848 100102
rect 318528 99978 318848 100046
rect 318528 99922 318598 99978
rect 318654 99922 318722 99978
rect 318778 99922 318848 99978
rect 318528 99888 318848 99922
rect 265132 98242 265188 98252
rect 272448 94350 272768 94384
rect 272448 94294 272518 94350
rect 272574 94294 272642 94350
rect 272698 94294 272768 94350
rect 272448 94226 272768 94294
rect 272448 94170 272518 94226
rect 272574 94170 272642 94226
rect 272698 94170 272768 94226
rect 272448 94102 272768 94170
rect 272448 94046 272518 94102
rect 272574 94046 272642 94102
rect 272698 94046 272768 94102
rect 272448 93978 272768 94046
rect 272448 93922 272518 93978
rect 272574 93922 272642 93978
rect 272698 93922 272768 93978
rect 272448 93888 272768 93922
rect 303168 94350 303488 94384
rect 303168 94294 303238 94350
rect 303294 94294 303362 94350
rect 303418 94294 303488 94350
rect 303168 94226 303488 94294
rect 303168 94170 303238 94226
rect 303294 94170 303362 94226
rect 303418 94170 303488 94226
rect 303168 94102 303488 94170
rect 303168 94046 303238 94102
rect 303294 94046 303362 94102
rect 303418 94046 303488 94102
rect 303168 93978 303488 94046
rect 303168 93922 303238 93978
rect 303294 93922 303362 93978
rect 303418 93922 303488 93978
rect 303168 93888 303488 93922
rect 265020 89842 265076 89852
rect 264796 86482 264852 86492
rect 264908 87556 264964 87566
rect 264908 77364 264964 87500
rect 287808 82350 288128 82384
rect 287808 82294 287878 82350
rect 287934 82294 288002 82350
rect 288058 82294 288128 82350
rect 287808 82226 288128 82294
rect 287808 82170 287878 82226
rect 287934 82170 288002 82226
rect 288058 82170 288128 82226
rect 287808 82102 288128 82170
rect 287808 82046 287878 82102
rect 287934 82046 288002 82102
rect 288058 82046 288128 82102
rect 287808 81978 288128 82046
rect 287808 81922 287878 81978
rect 287934 81922 288002 81978
rect 288058 81922 288128 81978
rect 287808 81888 288128 81922
rect 318528 82350 318848 82384
rect 318528 82294 318598 82350
rect 318654 82294 318722 82350
rect 318778 82294 318848 82350
rect 318528 82226 318848 82294
rect 318528 82170 318598 82226
rect 318654 82170 318722 82226
rect 318778 82170 318848 82226
rect 318528 82102 318848 82170
rect 318528 82046 318598 82102
rect 318654 82046 318722 82102
rect 318778 82046 318848 82102
rect 318528 81978 318848 82046
rect 318528 81922 318598 81978
rect 318654 81922 318722 81978
rect 318778 81922 318848 81978
rect 318528 81888 318848 81922
rect 264908 77298 264964 77308
rect 272448 76350 272768 76384
rect 272448 76294 272518 76350
rect 272574 76294 272642 76350
rect 272698 76294 272768 76350
rect 272448 76226 272768 76294
rect 272448 76170 272518 76226
rect 272574 76170 272642 76226
rect 272698 76170 272768 76226
rect 272448 76102 272768 76170
rect 272448 76046 272518 76102
rect 272574 76046 272642 76102
rect 272698 76046 272768 76102
rect 272448 75978 272768 76046
rect 272448 75922 272518 75978
rect 272574 75922 272642 75978
rect 272698 75922 272768 75978
rect 272448 75888 272768 75922
rect 303168 76350 303488 76384
rect 303168 76294 303238 76350
rect 303294 76294 303362 76350
rect 303418 76294 303488 76350
rect 303168 76226 303488 76294
rect 303168 76170 303238 76226
rect 303294 76170 303362 76226
rect 303418 76170 303488 76226
rect 303168 76102 303488 76170
rect 303168 76046 303238 76102
rect 303294 76046 303362 76102
rect 303418 76046 303488 76102
rect 303168 75978 303488 76046
rect 303168 75922 303238 75978
rect 303294 75922 303362 75978
rect 303418 75922 303488 75978
rect 303168 75888 303488 75922
rect 264572 74722 264628 74732
rect 333452 73220 333508 569582
rect 343338 562350 343958 579922
rect 343338 562294 343434 562350
rect 343490 562294 343558 562350
rect 343614 562294 343682 562350
rect 343738 562294 343806 562350
rect 343862 562294 343958 562350
rect 343338 562226 343958 562294
rect 343338 562170 343434 562226
rect 343490 562170 343558 562226
rect 343614 562170 343682 562226
rect 343738 562170 343806 562226
rect 343862 562170 343958 562226
rect 343338 562102 343958 562170
rect 343338 562046 343434 562102
rect 343490 562046 343558 562102
rect 343614 562046 343682 562102
rect 343738 562046 343806 562102
rect 343862 562046 343958 562102
rect 343338 561978 343958 562046
rect 343338 561922 343434 561978
rect 343490 561922 343558 561978
rect 343614 561922 343682 561978
rect 343738 561922 343806 561978
rect 343862 561922 343958 561978
rect 340284 553252 340340 553262
rect 338492 549220 338548 549230
rect 336812 519988 336868 519998
rect 335244 516628 335300 516638
rect 334460 511924 334516 511934
rect 334348 510244 334404 510254
rect 334348 507556 334404 510188
rect 334460 509796 334516 511868
rect 334460 509730 334516 509740
rect 334348 507490 334404 507500
rect 335132 506660 335188 506670
rect 335132 476196 335188 506604
rect 335244 488516 335300 516572
rect 335468 510132 335524 510142
rect 335244 488450 335300 488460
rect 335356 504868 335412 504878
rect 335356 477316 335412 504812
rect 335468 483476 335524 510076
rect 335916 503524 335972 503534
rect 335916 501956 335972 503468
rect 335916 501890 335972 501900
rect 336812 492996 336868 519932
rect 337708 505428 337764 505438
rect 337708 501396 337764 505372
rect 338492 503636 338548 549164
rect 340172 543844 340228 543854
rect 338716 506548 338772 506558
rect 338492 503570 338548 503580
rect 338604 505092 338660 505102
rect 337708 501330 337764 501340
rect 336812 492930 336868 492940
rect 335468 483410 335524 483420
rect 335580 488068 335636 488078
rect 335356 477250 335412 477260
rect 335132 476130 335188 476140
rect 335356 475524 335412 475534
rect 334460 473698 334516 473708
rect 334460 473396 334516 473642
rect 334460 473330 334516 473340
rect 334348 471156 334404 471166
rect 334348 470458 334404 471100
rect 334460 470638 334516 470648
rect 334460 470530 334516 470540
rect 334460 470458 334516 470468
rect 334348 470402 334460 470458
rect 334460 470392 334516 470402
rect 334460 469558 334516 469568
rect 334460 468916 334516 469502
rect 334460 468850 334516 468860
rect 334460 466138 334516 466148
rect 334348 466082 334460 466138
rect 334348 460516 334404 466082
rect 334460 466072 334516 466082
rect 334460 465238 334516 465248
rect 334460 464436 334516 465182
rect 334460 464370 334516 464380
rect 334460 462898 334516 462908
rect 334460 461076 334516 462842
rect 334460 461010 334516 461020
rect 334348 460450 334404 460460
rect 335356 459956 335412 475468
rect 335580 474516 335636 488012
rect 335580 474450 335636 474460
rect 335804 483812 335860 483822
rect 335804 473956 335860 483756
rect 338604 481236 338660 505036
rect 338716 487396 338772 506492
rect 338716 487330 338772 487340
rect 340172 483812 340228 543788
rect 340284 504756 340340 553196
rect 341964 551684 342020 551694
rect 341852 545188 341908 545198
rect 340284 504690 340340 504700
rect 340396 511588 340452 511598
rect 340396 487956 340452 511532
rect 340396 487890 340452 487900
rect 340172 483746 340228 483756
rect 338604 481170 338660 481180
rect 339388 480538 339444 480548
rect 339388 475524 339444 480482
rect 341852 478436 341908 545132
rect 341964 508116 342020 551628
rect 343338 544350 343958 561922
rect 347058 598172 347678 598268
rect 347058 598116 347154 598172
rect 347210 598116 347278 598172
rect 347334 598116 347402 598172
rect 347458 598116 347526 598172
rect 347582 598116 347678 598172
rect 347058 598048 347678 598116
rect 347058 597992 347154 598048
rect 347210 597992 347278 598048
rect 347334 597992 347402 598048
rect 347458 597992 347526 598048
rect 347582 597992 347678 598048
rect 347058 597924 347678 597992
rect 347058 597868 347154 597924
rect 347210 597868 347278 597924
rect 347334 597868 347402 597924
rect 347458 597868 347526 597924
rect 347582 597868 347678 597924
rect 347058 597800 347678 597868
rect 347058 597744 347154 597800
rect 347210 597744 347278 597800
rect 347334 597744 347402 597800
rect 347458 597744 347526 597800
rect 347582 597744 347678 597800
rect 347058 586350 347678 597744
rect 347058 586294 347154 586350
rect 347210 586294 347278 586350
rect 347334 586294 347402 586350
rect 347458 586294 347526 586350
rect 347582 586294 347678 586350
rect 347058 586226 347678 586294
rect 347058 586170 347154 586226
rect 347210 586170 347278 586226
rect 347334 586170 347402 586226
rect 347458 586170 347526 586226
rect 347582 586170 347678 586226
rect 347058 586102 347678 586170
rect 347058 586046 347154 586102
rect 347210 586046 347278 586102
rect 347334 586046 347402 586102
rect 347458 586046 347526 586102
rect 347582 586046 347678 586102
rect 347058 585978 347678 586046
rect 347058 585922 347154 585978
rect 347210 585922 347278 585978
rect 347334 585922 347402 585978
rect 347458 585922 347526 585978
rect 347582 585922 347678 585978
rect 347058 568350 347678 585922
rect 347058 568294 347154 568350
rect 347210 568294 347278 568350
rect 347334 568294 347402 568350
rect 347458 568294 347526 568350
rect 347582 568294 347678 568350
rect 347058 568226 347678 568294
rect 347058 568170 347154 568226
rect 347210 568170 347278 568226
rect 347334 568170 347402 568226
rect 347458 568170 347526 568226
rect 347582 568170 347678 568226
rect 347058 568102 347678 568170
rect 347058 568046 347154 568102
rect 347210 568046 347278 568102
rect 347334 568046 347402 568102
rect 347458 568046 347526 568102
rect 347582 568046 347678 568102
rect 347058 567978 347678 568046
rect 347058 567922 347154 567978
rect 347210 567922 347278 567978
rect 347334 567922 347402 567978
rect 347458 567922 347526 567978
rect 347582 567922 347678 567978
rect 343338 544294 343434 544350
rect 343490 544294 343558 544350
rect 343614 544294 343682 544350
rect 343738 544294 343806 544350
rect 343862 544294 343958 544350
rect 343338 544226 343958 544294
rect 343338 544170 343434 544226
rect 343490 544170 343558 544226
rect 343614 544170 343682 544226
rect 343738 544170 343806 544226
rect 343862 544170 343958 544226
rect 343338 544102 343958 544170
rect 343338 544046 343434 544102
rect 343490 544046 343558 544102
rect 343614 544046 343682 544102
rect 343738 544046 343806 544102
rect 343862 544046 343958 544102
rect 343338 543978 343958 544046
rect 343338 543922 343434 543978
rect 343490 543922 343558 543978
rect 343614 543922 343682 543978
rect 343738 543922 343806 543978
rect 343862 543922 343958 543978
rect 343338 526350 343958 543922
rect 343338 526294 343434 526350
rect 343490 526294 343558 526350
rect 343614 526294 343682 526350
rect 343738 526294 343806 526350
rect 343862 526294 343958 526350
rect 343338 526226 343958 526294
rect 343338 526170 343434 526226
rect 343490 526170 343558 526226
rect 343614 526170 343682 526226
rect 343738 526170 343806 526226
rect 343862 526170 343958 526226
rect 343338 526102 343958 526170
rect 343338 526046 343434 526102
rect 343490 526046 343558 526102
rect 343614 526046 343682 526102
rect 343738 526046 343806 526102
rect 343862 526046 343958 526102
rect 343338 525978 343958 526046
rect 343338 525922 343434 525978
rect 343490 525922 343558 525978
rect 343614 525922 343682 525978
rect 343738 525922 343806 525978
rect 343862 525922 343958 525978
rect 341964 508050 342020 508060
rect 342076 513380 342132 513390
rect 342076 490196 342132 513324
rect 343338 508350 343958 525922
rect 342076 490130 342132 490140
rect 342188 508340 342244 508350
rect 342188 484036 342244 508284
rect 342188 483970 342244 483980
rect 343338 508294 343434 508350
rect 343490 508294 343558 508350
rect 343614 508294 343682 508350
rect 343738 508294 343806 508350
rect 343862 508294 343958 508350
rect 343338 508226 343958 508294
rect 343338 508170 343434 508226
rect 343490 508170 343558 508226
rect 343614 508170 343682 508226
rect 343738 508170 343806 508226
rect 343862 508170 343958 508226
rect 343338 508102 343958 508170
rect 343338 508046 343434 508102
rect 343490 508046 343558 508102
rect 343614 508046 343682 508102
rect 343738 508046 343806 508102
rect 343862 508046 343958 508102
rect 343338 507978 343958 508046
rect 343338 507922 343434 507978
rect 343490 507922 343558 507978
rect 343614 507922 343682 507978
rect 343738 507922 343806 507978
rect 343862 507922 343958 507978
rect 343338 490350 343958 507922
rect 345212 550564 345268 550574
rect 343338 490294 343434 490350
rect 343490 490294 343558 490350
rect 343614 490294 343682 490350
rect 343738 490294 343806 490350
rect 343862 490294 343958 490350
rect 343338 490226 343958 490294
rect 343338 490170 343434 490226
rect 343490 490170 343558 490226
rect 343614 490170 343682 490226
rect 343738 490170 343806 490226
rect 343862 490170 343958 490226
rect 343338 490102 343958 490170
rect 343338 490046 343434 490102
rect 343490 490046 343558 490102
rect 343614 490046 343682 490102
rect 343738 490046 343806 490102
rect 343862 490046 343958 490102
rect 343338 489978 343958 490046
rect 343338 489922 343434 489978
rect 343490 489922 343558 489978
rect 343614 489922 343682 489978
rect 343738 489922 343806 489978
rect 343862 489922 343958 489978
rect 341852 478370 341908 478380
rect 342076 478660 342132 478670
rect 339388 475458 339444 475468
rect 340172 476644 340228 476654
rect 335804 473890 335860 473900
rect 335356 459890 335412 459900
rect 336028 458052 336084 458062
rect 336028 452116 336084 457996
rect 336140 456372 336196 456382
rect 336140 452676 336196 456316
rect 337708 456148 337764 456158
rect 337708 453796 337764 456092
rect 337708 453730 337764 453740
rect 336140 452610 336196 452620
rect 336028 452050 336084 452060
rect 335132 451220 335188 451230
rect 334460 427588 334516 427598
rect 334460 423556 334516 427532
rect 334460 423490 334516 423500
rect 335132 420756 335188 451164
rect 336812 447860 336868 447870
rect 335804 446068 335860 446078
rect 335804 442596 335860 446012
rect 335916 444724 335972 444734
rect 335916 443156 335972 444668
rect 335916 443090 335972 443100
rect 335804 442530 335860 442540
rect 335132 420690 335188 420700
rect 335356 437668 335412 437678
rect 335356 419076 335412 437612
rect 335804 432628 335860 432638
rect 335804 426916 335860 432572
rect 335804 426850 335860 426860
rect 336812 424116 336868 447804
rect 338492 444612 338548 444622
rect 338492 429156 338548 444556
rect 338492 429090 338548 429100
rect 336812 424050 336868 424060
rect 340172 420196 340228 476588
rect 342076 444276 342132 478604
rect 343338 472350 343958 489922
rect 344092 501508 344148 501518
rect 344092 489636 344148 501452
rect 344092 489570 344148 489580
rect 345212 488068 345268 550508
rect 347058 550350 347678 567922
rect 374058 597212 374678 598268
rect 374058 597156 374154 597212
rect 374210 597156 374278 597212
rect 374334 597156 374402 597212
rect 374458 597156 374526 597212
rect 374582 597156 374678 597212
rect 374058 597088 374678 597156
rect 374058 597032 374154 597088
rect 374210 597032 374278 597088
rect 374334 597032 374402 597088
rect 374458 597032 374526 597088
rect 374582 597032 374678 597088
rect 374058 596964 374678 597032
rect 374058 596908 374154 596964
rect 374210 596908 374278 596964
rect 374334 596908 374402 596964
rect 374458 596908 374526 596964
rect 374582 596908 374678 596964
rect 374058 596840 374678 596908
rect 374058 596784 374154 596840
rect 374210 596784 374278 596840
rect 374334 596784 374402 596840
rect 374458 596784 374526 596840
rect 374582 596784 374678 596840
rect 374058 580350 374678 596784
rect 374058 580294 374154 580350
rect 374210 580294 374278 580350
rect 374334 580294 374402 580350
rect 374458 580294 374526 580350
rect 374582 580294 374678 580350
rect 374058 580226 374678 580294
rect 374058 580170 374154 580226
rect 374210 580170 374278 580226
rect 374334 580170 374402 580226
rect 374458 580170 374526 580226
rect 374582 580170 374678 580226
rect 374058 580102 374678 580170
rect 374058 580046 374154 580102
rect 374210 580046 374278 580102
rect 374334 580046 374402 580102
rect 374458 580046 374526 580102
rect 374582 580046 374678 580102
rect 374058 579978 374678 580046
rect 374058 579922 374154 579978
rect 374210 579922 374278 579978
rect 374334 579922 374402 579978
rect 374458 579922 374526 579978
rect 374582 579922 374678 579978
rect 356448 562350 356768 562384
rect 356448 562294 356518 562350
rect 356574 562294 356642 562350
rect 356698 562294 356768 562350
rect 356448 562226 356768 562294
rect 356448 562170 356518 562226
rect 356574 562170 356642 562226
rect 356698 562170 356768 562226
rect 356448 562102 356768 562170
rect 356448 562046 356518 562102
rect 356574 562046 356642 562102
rect 356698 562046 356768 562102
rect 356448 561978 356768 562046
rect 356448 561922 356518 561978
rect 356574 561922 356642 561978
rect 356698 561922 356768 561978
rect 356448 561888 356768 561922
rect 374058 562350 374678 579922
rect 374058 562294 374154 562350
rect 374210 562294 374278 562350
rect 374334 562294 374402 562350
rect 374458 562294 374526 562350
rect 374582 562294 374678 562350
rect 374058 562226 374678 562294
rect 374058 562170 374154 562226
rect 374210 562170 374278 562226
rect 374334 562170 374402 562226
rect 374458 562170 374526 562226
rect 374582 562170 374678 562226
rect 374058 562102 374678 562170
rect 374058 562046 374154 562102
rect 374210 562046 374278 562102
rect 374334 562046 374402 562102
rect 374458 562046 374526 562102
rect 374582 562046 374678 562102
rect 374058 561978 374678 562046
rect 374058 561922 374154 561978
rect 374210 561922 374278 561978
rect 374334 561922 374402 561978
rect 374458 561922 374526 561978
rect 374582 561922 374678 561978
rect 352716 555268 352772 555278
rect 352716 555172 352772 555182
rect 347788 553924 347844 553934
rect 347788 551684 347844 553868
rect 347788 551618 347844 551628
rect 347058 550294 347154 550350
rect 347210 550294 347278 550350
rect 347334 550294 347402 550350
rect 347458 550294 347526 550350
rect 347582 550294 347678 550350
rect 347058 550226 347678 550294
rect 347058 550170 347154 550226
rect 347210 550170 347278 550226
rect 347334 550170 347402 550226
rect 347458 550170 347526 550226
rect 347582 550170 347678 550226
rect 347058 550102 347678 550170
rect 347058 550046 347154 550102
rect 347210 550046 347278 550102
rect 347334 550046 347402 550102
rect 347458 550046 347526 550102
rect 347582 550046 347678 550102
rect 347058 549978 347678 550046
rect 347058 549922 347154 549978
rect 347210 549922 347278 549978
rect 347334 549922 347402 549978
rect 347458 549922 347526 549978
rect 347582 549922 347678 549978
rect 347058 532350 347678 549922
rect 347058 532294 347154 532350
rect 347210 532294 347278 532350
rect 347334 532294 347402 532350
rect 347458 532294 347526 532350
rect 347582 532294 347678 532350
rect 347058 532226 347678 532294
rect 347058 532170 347154 532226
rect 347210 532170 347278 532226
rect 347334 532170 347402 532226
rect 347458 532170 347526 532226
rect 347582 532170 347678 532226
rect 347058 532102 347678 532170
rect 347058 532046 347154 532102
rect 347210 532046 347278 532102
rect 347334 532046 347402 532102
rect 347458 532046 347526 532102
rect 347582 532046 347678 532102
rect 347058 531978 347678 532046
rect 347058 531922 347154 531978
rect 347210 531922 347278 531978
rect 347334 531922 347402 531978
rect 347458 531922 347526 531978
rect 347582 531922 347678 531978
rect 347058 514350 347678 531922
rect 347058 514294 347154 514350
rect 347210 514294 347278 514350
rect 347334 514294 347402 514350
rect 347458 514294 347526 514350
rect 347582 514294 347678 514350
rect 347058 514226 347678 514294
rect 347058 514170 347154 514226
rect 347210 514170 347278 514226
rect 347334 514170 347402 514226
rect 347458 514170 347526 514226
rect 347582 514170 347678 514226
rect 347058 514102 347678 514170
rect 347058 514046 347154 514102
rect 347210 514046 347278 514102
rect 347334 514046 347402 514102
rect 347458 514046 347526 514102
rect 347582 514046 347678 514102
rect 347058 513978 347678 514046
rect 347058 513922 347154 513978
rect 347210 513922 347278 513978
rect 347334 513922 347402 513978
rect 347458 513922 347526 513978
rect 347582 513922 347678 513978
rect 345548 513268 345604 513278
rect 345324 510020 345380 510030
rect 345324 491876 345380 509964
rect 345548 499156 345604 513212
rect 345548 499090 345604 499100
rect 345324 491810 345380 491820
rect 347058 496350 347678 513922
rect 347058 496294 347154 496350
rect 347210 496294 347278 496350
rect 347334 496294 347402 496350
rect 347458 496294 347526 496350
rect 347582 496294 347678 496350
rect 347058 496226 347678 496294
rect 347058 496170 347154 496226
rect 347210 496170 347278 496226
rect 347334 496170 347402 496226
rect 347458 496170 347526 496226
rect 347582 496170 347678 496226
rect 347058 496102 347678 496170
rect 347058 496046 347154 496102
rect 347210 496046 347278 496102
rect 347334 496046 347402 496102
rect 347458 496046 347526 496102
rect 347582 496046 347678 496102
rect 347058 495978 347678 496046
rect 347058 495922 347154 495978
rect 347210 495922 347278 495978
rect 347334 495922 347402 495978
rect 347458 495922 347526 495978
rect 347582 495922 347678 495978
rect 345212 488002 345268 488012
rect 347058 478350 347678 495922
rect 348572 551236 348628 551246
rect 348572 479556 348628 551180
rect 371808 550350 372128 550384
rect 371808 550294 371878 550350
rect 371934 550294 372002 550350
rect 372058 550294 372128 550350
rect 371808 550226 372128 550294
rect 371808 550170 371878 550226
rect 371934 550170 372002 550226
rect 372058 550170 372128 550226
rect 371808 550102 372128 550170
rect 371808 550046 371878 550102
rect 371934 550046 372002 550102
rect 372058 550046 372128 550102
rect 371808 549978 372128 550046
rect 371808 549922 371878 549978
rect 371934 549922 372002 549978
rect 372058 549922 372128 549978
rect 348684 549892 348740 549902
rect 371808 549888 372128 549922
rect 348684 503524 348740 549836
rect 356448 544350 356768 544384
rect 356448 544294 356518 544350
rect 356574 544294 356642 544350
rect 356698 544294 356768 544350
rect 356448 544226 356768 544294
rect 356448 544170 356518 544226
rect 356574 544170 356642 544226
rect 356698 544170 356768 544226
rect 356448 544102 356768 544170
rect 356448 544046 356518 544102
rect 356574 544046 356642 544102
rect 356698 544046 356768 544102
rect 356448 543978 356768 544046
rect 356448 543922 356518 543978
rect 356574 543922 356642 543978
rect 356698 543922 356768 543978
rect 356448 543888 356768 543922
rect 374058 544350 374678 561922
rect 374058 544294 374154 544350
rect 374210 544294 374278 544350
rect 374334 544294 374402 544350
rect 374458 544294 374526 544350
rect 374582 544294 374678 544350
rect 374058 544226 374678 544294
rect 374058 544170 374154 544226
rect 374210 544170 374278 544226
rect 374334 544170 374402 544226
rect 374458 544170 374526 544226
rect 374582 544170 374678 544226
rect 374058 544102 374678 544170
rect 374058 544046 374154 544102
rect 374210 544046 374278 544102
rect 374334 544046 374402 544102
rect 374458 544046 374526 544102
rect 374582 544046 374678 544102
rect 374058 543978 374678 544046
rect 374058 543922 374154 543978
rect 374210 543922 374278 543978
rect 374334 543922 374402 543978
rect 374458 543922 374526 543978
rect 374582 543922 374678 543978
rect 371808 532350 372128 532384
rect 371808 532294 371878 532350
rect 371934 532294 372002 532350
rect 372058 532294 372128 532350
rect 371808 532226 372128 532294
rect 371808 532170 371878 532226
rect 371934 532170 372002 532226
rect 372058 532170 372128 532226
rect 371808 532102 372128 532170
rect 371808 532046 371878 532102
rect 371934 532046 372002 532102
rect 372058 532046 372128 532102
rect 371808 531978 372128 532046
rect 371808 531922 371878 531978
rect 371934 531922 372002 531978
rect 372058 531922 372128 531978
rect 371808 531888 372128 531922
rect 354396 528052 354452 528062
rect 354396 526036 354452 527996
rect 354396 525970 354452 525980
rect 357756 527940 357812 527950
rect 348684 503458 348740 503468
rect 348796 523348 348852 523358
rect 348796 493556 348852 523292
rect 357756 522116 357812 527884
rect 357756 522050 357812 522060
rect 374058 526350 374678 543922
rect 374058 526294 374154 526350
rect 374210 526294 374278 526350
rect 374334 526294 374402 526350
rect 374458 526294 374526 526350
rect 374582 526294 374678 526350
rect 374058 526226 374678 526294
rect 374058 526170 374154 526226
rect 374210 526170 374278 526226
rect 374334 526170 374402 526226
rect 374458 526170 374526 526226
rect 374582 526170 374678 526226
rect 374058 526102 374678 526170
rect 374058 526046 374154 526102
rect 374210 526046 374278 526102
rect 374334 526046 374402 526102
rect 374458 526046 374526 526102
rect 374582 526046 374678 526102
rect 374058 525978 374678 526046
rect 374058 525922 374154 525978
rect 374210 525922 374278 525978
rect 374334 525922 374402 525978
rect 374458 525922 374526 525978
rect 374582 525922 374678 525978
rect 351932 522004 351988 522014
rect 350588 506884 350644 506894
rect 348796 493490 348852 493500
rect 348908 505204 348964 505214
rect 348908 485716 348964 505148
rect 348908 485650 348964 485660
rect 349020 503524 349076 503534
rect 349020 480116 349076 503468
rect 350588 484596 350644 506828
rect 350588 484530 350644 484540
rect 349020 480050 349076 480060
rect 348572 479490 348628 479500
rect 348796 480004 348852 480014
rect 347058 478294 347154 478350
rect 347210 478294 347278 478350
rect 347334 478294 347402 478350
rect 347458 478294 347526 478350
rect 347582 478294 347678 478350
rect 347058 478226 347678 478294
rect 347058 478170 347154 478226
rect 347210 478170 347278 478226
rect 347334 478170 347402 478226
rect 347458 478170 347526 478226
rect 347582 478170 347678 478226
rect 347058 478102 347678 478170
rect 347058 478046 347154 478102
rect 347210 478046 347278 478102
rect 347334 478046 347402 478102
rect 347458 478046 347526 478102
rect 347582 478046 347678 478102
rect 347058 477978 347678 478046
rect 347058 477922 347154 477978
rect 347210 477922 347278 477978
rect 347334 477922 347402 477978
rect 347458 477922 347526 477978
rect 347582 477922 347678 477978
rect 343338 472294 343434 472350
rect 343490 472294 343558 472350
rect 343614 472294 343682 472350
rect 343738 472294 343806 472350
rect 343862 472294 343958 472350
rect 343338 472226 343958 472294
rect 343338 472170 343434 472226
rect 343490 472170 343558 472226
rect 343614 472170 343682 472226
rect 343738 472170 343806 472226
rect 343862 472170 343958 472226
rect 343338 472102 343958 472170
rect 343338 472046 343434 472102
rect 343490 472046 343558 472102
rect 343614 472046 343682 472102
rect 343738 472046 343806 472102
rect 343862 472046 343958 472102
rect 343338 471978 343958 472046
rect 343338 471922 343434 471978
rect 343490 471922 343558 471978
rect 343614 471922 343682 471978
rect 343738 471922 343806 471978
rect 343862 471922 343958 471978
rect 343338 454350 343958 471922
rect 343338 454294 343434 454350
rect 343490 454294 343558 454350
rect 343614 454294 343682 454350
rect 343738 454294 343806 454350
rect 343862 454294 343958 454350
rect 343338 454226 343958 454294
rect 343338 454170 343434 454226
rect 343490 454170 343558 454226
rect 343614 454170 343682 454226
rect 343738 454170 343806 454226
rect 343862 454170 343958 454226
rect 343338 454102 343958 454170
rect 343338 454046 343434 454102
rect 343490 454046 343558 454102
rect 343614 454046 343682 454102
rect 343738 454046 343806 454102
rect 343862 454046 343958 454102
rect 343338 453978 343958 454046
rect 343338 453922 343434 453978
rect 343490 453922 343558 453978
rect 343614 453922 343682 453978
rect 343738 453922 343806 453978
rect 343862 453922 343958 453978
rect 342076 444210 342132 444220
rect 342188 449652 342244 449662
rect 340172 420130 340228 420140
rect 342188 419636 342244 449596
rect 342300 446292 342356 446302
rect 342300 425236 342356 446236
rect 342300 425170 342356 425180
rect 343338 436350 343958 453922
rect 345212 473844 345268 473854
rect 345212 449876 345268 473788
rect 345212 449810 345268 449820
rect 347058 460350 347678 477922
rect 348684 479332 348740 479342
rect 347058 460294 347154 460350
rect 347210 460294 347278 460350
rect 347334 460294 347402 460350
rect 347458 460294 347526 460350
rect 347582 460294 347678 460350
rect 347058 460226 347678 460294
rect 347058 460170 347154 460226
rect 347210 460170 347278 460226
rect 347334 460170 347402 460226
rect 347458 460170 347526 460226
rect 347582 460170 347678 460226
rect 347058 460102 347678 460170
rect 347058 460046 347154 460102
rect 347210 460046 347278 460102
rect 347334 460046 347402 460102
rect 347458 460046 347526 460102
rect 347582 460046 347678 460102
rect 347058 459978 347678 460046
rect 347058 459922 347154 459978
rect 347210 459922 347278 459978
rect 347334 459922 347402 459978
rect 347458 459922 347526 459978
rect 347582 459922 347678 459978
rect 344428 446628 344484 446638
rect 344428 444836 344484 446572
rect 344428 444770 344484 444780
rect 343338 436294 343434 436350
rect 343490 436294 343558 436350
rect 343614 436294 343682 436350
rect 343738 436294 343806 436350
rect 343862 436294 343958 436350
rect 343338 436226 343958 436294
rect 343338 436170 343434 436226
rect 343490 436170 343558 436226
rect 343614 436170 343682 436226
rect 343738 436170 343806 436226
rect 343862 436170 343958 436226
rect 343338 436102 343958 436170
rect 343338 436046 343434 436102
rect 343490 436046 343558 436102
rect 343614 436046 343682 436102
rect 343738 436046 343806 436102
rect 343862 436046 343958 436102
rect 343338 435978 343958 436046
rect 343338 435922 343434 435978
rect 343490 435922 343558 435978
rect 343614 435922 343682 435978
rect 343738 435922 343806 435978
rect 343862 435922 343958 435978
rect 342188 419570 342244 419580
rect 335356 419010 335412 419020
rect 343338 418350 343958 435922
rect 343338 418294 343434 418350
rect 343490 418294 343558 418350
rect 343614 418294 343682 418350
rect 343738 418294 343806 418350
rect 343862 418294 343958 418350
rect 343338 418226 343958 418294
rect 343338 418170 343434 418226
rect 343490 418170 343558 418226
rect 343614 418170 343682 418226
rect 343738 418170 343806 418226
rect 343862 418170 343958 418226
rect 343338 418102 343958 418170
rect 343338 418046 343434 418102
rect 343490 418046 343558 418102
rect 343614 418046 343682 418102
rect 343738 418046 343806 418102
rect 343862 418046 343958 418102
rect 343338 417978 343958 418046
rect 343338 417922 343434 417978
rect 343490 417922 343558 417978
rect 343614 417922 343682 417978
rect 343738 417922 343806 417978
rect 343862 417922 343958 417978
rect 334460 415156 334516 415166
rect 334460 415018 334516 415100
rect 334460 414952 334516 414962
rect 334460 414596 334516 414606
rect 334460 413758 334516 414540
rect 334460 413692 334516 413702
rect 334460 413578 334516 413588
rect 334460 413476 334516 413522
rect 334460 413410 334516 413420
rect 334348 412356 334404 412366
rect 334348 411778 334404 412300
rect 334460 411958 334516 411968
rect 334460 411796 334516 411902
rect 334460 411730 334516 411740
rect 334348 411712 334404 411722
rect 334460 411236 334516 411246
rect 334460 410698 334516 411180
rect 334460 410632 334516 410642
rect 334348 410116 334404 410126
rect 334348 409108 334404 410060
rect 338604 410116 338660 410126
rect 334460 409618 334516 409628
rect 334460 409556 334516 409562
rect 334460 409490 334516 409500
rect 334348 409042 334404 409052
rect 334460 408178 334516 408188
rect 334460 407876 334516 408122
rect 334460 407810 334516 407820
rect 338492 408100 338548 408110
rect 334460 407458 334516 407468
rect 334348 407402 334460 407458
rect 334348 401156 334404 407402
rect 334460 407392 334516 407402
rect 336252 406738 336308 406748
rect 336028 405636 336084 405646
rect 336028 404758 336084 405580
rect 336028 404692 336084 404702
rect 334460 403956 334516 403966
rect 334460 403318 334516 403900
rect 334460 403252 334516 403262
rect 334460 403138 334516 403148
rect 334460 402836 334516 403082
rect 334460 402770 334516 402780
rect 334348 401090 334404 401100
rect 334460 399718 334516 399728
rect 334460 398916 334516 399662
rect 336252 399476 336308 406682
rect 336252 399410 336308 399420
rect 334460 398850 334516 398860
rect 336812 399028 336868 399038
rect 334460 398098 334516 398108
rect 334348 398042 334460 398098
rect 334348 396676 334404 398042
rect 334460 398032 334516 398042
rect 334460 397918 334516 397928
rect 334460 397236 334516 397862
rect 334460 397170 334516 397180
rect 334348 396610 334404 396620
rect 334460 396478 334516 396488
rect 334348 396298 334404 396308
rect 334348 395556 334404 396242
rect 334460 396116 334516 396422
rect 334460 396050 334516 396060
rect 334348 395490 334404 395500
rect 334460 394678 334516 394688
rect 334348 394622 334460 394678
rect 334348 393876 334404 394622
rect 334460 394612 334516 394622
rect 334460 394498 334516 394508
rect 334460 394436 334516 394442
rect 334460 394370 334516 394380
rect 334348 393810 334404 393820
rect 334460 393058 334516 393068
rect 334348 392756 334404 392766
rect 334348 391618 334404 392700
rect 334460 392196 334516 393002
rect 334460 392130 334516 392140
rect 334460 391618 334516 391628
rect 334348 391562 334460 391618
rect 334460 391552 334516 391562
rect 336812 386596 336868 398972
rect 336812 386530 336868 386540
rect 335244 380548 335300 380558
rect 335132 378868 335188 378878
rect 334572 368788 334628 368798
rect 334348 367108 334404 367118
rect 334348 364756 334404 367052
rect 334348 364690 334404 364700
rect 334460 365540 334516 365550
rect 334460 363076 334516 365484
rect 334460 363010 334516 363020
rect 334572 362516 334628 368732
rect 335132 363636 335188 378812
rect 335244 369796 335300 380492
rect 336140 375508 336196 375518
rect 336140 370356 336196 375452
rect 336140 370290 336196 370300
rect 335244 369730 335300 369740
rect 335132 363570 335188 363580
rect 334572 362450 334628 362460
rect 335916 362068 335972 362078
rect 335916 357476 335972 362012
rect 338492 358036 338548 408044
rect 338604 387716 338660 410060
rect 341852 406084 341908 406094
rect 340508 403284 340564 403294
rect 340508 388276 340564 403228
rect 340508 388210 340564 388220
rect 338604 387650 338660 387660
rect 341852 360276 341908 406028
rect 341852 360210 341908 360220
rect 343338 400350 343958 417922
rect 347058 442350 347678 459922
rect 347058 442294 347154 442350
rect 347210 442294 347278 442350
rect 347334 442294 347402 442350
rect 347458 442294 347526 442350
rect 347582 442294 347678 442350
rect 347058 442226 347678 442294
rect 347058 442170 347154 442226
rect 347210 442170 347278 442226
rect 347334 442170 347402 442226
rect 347458 442170 347526 442226
rect 347582 442170 347678 442226
rect 347058 442102 347678 442170
rect 347058 442046 347154 442102
rect 347210 442046 347278 442102
rect 347334 442046 347402 442102
rect 347458 442046 347526 442102
rect 347582 442046 347678 442102
rect 347058 441978 347678 442046
rect 347058 441922 347154 441978
rect 347210 441922 347278 441978
rect 347334 441922 347402 441978
rect 347458 441922 347526 441978
rect 347582 441922 347678 441978
rect 347058 424350 347678 441922
rect 347058 424294 347154 424350
rect 347210 424294 347278 424350
rect 347334 424294 347402 424350
rect 347458 424294 347526 424350
rect 347582 424294 347678 424350
rect 347058 424226 347678 424294
rect 347058 424170 347154 424226
rect 347210 424170 347278 424226
rect 347334 424170 347402 424226
rect 347458 424170 347526 424226
rect 347582 424170 347678 424226
rect 347058 424102 347678 424170
rect 347058 424046 347154 424102
rect 347210 424046 347278 424102
rect 347334 424046 347402 424102
rect 347458 424046 347526 424102
rect 347582 424046 347678 424102
rect 347058 423978 347678 424046
rect 347058 423922 347154 423978
rect 347210 423922 347278 423978
rect 347334 423922 347402 423978
rect 347458 423922 347526 423978
rect 347582 423922 347678 423978
rect 347058 406350 347678 423922
rect 348572 473956 348628 473966
rect 348572 421316 348628 473900
rect 348684 473844 348740 479276
rect 348684 473778 348740 473788
rect 348796 446068 348852 479948
rect 351932 475076 351988 521948
rect 355292 520212 355348 520222
rect 353612 518308 353668 518318
rect 352156 506772 352212 506782
rect 352156 481796 352212 506716
rect 352268 504980 352324 504990
rect 352268 491316 352324 504924
rect 353612 495012 353668 518252
rect 353724 516740 353780 516750
rect 353724 497476 353780 516684
rect 355292 512036 355348 520156
rect 355292 511970 355348 511980
rect 354396 511700 354452 511710
rect 354396 510356 354452 511644
rect 354396 510290 354452 510300
rect 353836 509908 353892 509918
rect 353836 499716 353892 509852
rect 353836 499650 353892 499660
rect 374058 508350 374678 525922
rect 374058 508294 374154 508350
rect 374210 508294 374278 508350
rect 374334 508294 374402 508350
rect 374458 508294 374526 508350
rect 374582 508294 374678 508350
rect 374058 508226 374678 508294
rect 374058 508170 374154 508226
rect 374210 508170 374278 508226
rect 374334 508170 374402 508226
rect 374458 508170 374526 508226
rect 374582 508170 374678 508226
rect 374058 508102 374678 508170
rect 374058 508046 374154 508102
rect 374210 508046 374278 508102
rect 374334 508046 374402 508102
rect 374458 508046 374526 508102
rect 374582 508046 374678 508102
rect 374058 507978 374678 508046
rect 374058 507922 374154 507978
rect 374210 507922 374278 507978
rect 374334 507922 374402 507978
rect 374458 507922 374526 507978
rect 374582 507922 374678 507978
rect 353724 497410 353780 497420
rect 353612 494946 353668 494956
rect 352268 491250 352324 491260
rect 356448 490350 356768 490384
rect 356448 490294 356518 490350
rect 356574 490294 356642 490350
rect 356698 490294 356768 490350
rect 356448 490226 356768 490294
rect 356448 490170 356518 490226
rect 356574 490170 356642 490226
rect 356698 490170 356768 490226
rect 356448 490102 356768 490170
rect 356448 490046 356518 490102
rect 356574 490046 356642 490102
rect 356698 490046 356768 490102
rect 356448 489978 356768 490046
rect 356448 489922 356518 489978
rect 356574 489922 356642 489978
rect 356698 489922 356768 489978
rect 356448 489888 356768 489922
rect 374058 490350 374678 507922
rect 374058 490294 374154 490350
rect 374210 490294 374278 490350
rect 374334 490294 374402 490350
rect 374458 490294 374526 490350
rect 374582 490294 374678 490350
rect 374058 490226 374678 490294
rect 374058 490170 374154 490226
rect 374210 490170 374278 490226
rect 374334 490170 374402 490226
rect 374458 490170 374526 490226
rect 374582 490170 374678 490226
rect 374058 490102 374678 490170
rect 374058 490046 374154 490102
rect 374210 490046 374278 490102
rect 374334 490046 374402 490102
rect 374458 490046 374526 490102
rect 374582 490046 374678 490102
rect 374058 489978 374678 490046
rect 374058 489922 374154 489978
rect 374210 489922 374278 489978
rect 374334 489922 374402 489978
rect 374458 489922 374526 489978
rect 374582 489922 374678 489978
rect 352716 483364 352772 483374
rect 352716 483058 352772 483308
rect 352716 482992 352772 483002
rect 352156 481730 352212 481740
rect 371808 478350 372128 478384
rect 371808 478294 371878 478350
rect 371934 478294 372002 478350
rect 372058 478294 372128 478350
rect 371808 478226 372128 478294
rect 371808 478170 371878 478226
rect 371934 478170 372002 478226
rect 372058 478170 372128 478226
rect 371808 478102 372128 478170
rect 371808 478046 371878 478102
rect 371934 478046 372002 478102
rect 372058 478046 372128 478102
rect 371808 477978 372128 478046
rect 371808 477922 371878 477978
rect 371934 477922 372002 477978
rect 372058 477922 372128 477978
rect 371808 477888 372128 477922
rect 351932 475010 351988 475020
rect 356448 472350 356768 472384
rect 356448 472294 356518 472350
rect 356574 472294 356642 472350
rect 356698 472294 356768 472350
rect 356448 472226 356768 472294
rect 356448 472170 356518 472226
rect 356574 472170 356642 472226
rect 356698 472170 356768 472226
rect 356448 472102 356768 472170
rect 356448 472046 356518 472102
rect 356574 472046 356642 472102
rect 356698 472046 356768 472102
rect 356448 471978 356768 472046
rect 356448 471922 356518 471978
rect 356574 471922 356642 471978
rect 356698 471922 356768 471978
rect 356448 471888 356768 471922
rect 374058 472350 374678 489922
rect 374058 472294 374154 472350
rect 374210 472294 374278 472350
rect 374334 472294 374402 472350
rect 374458 472294 374526 472350
rect 374582 472294 374678 472350
rect 374058 472226 374678 472294
rect 374058 472170 374154 472226
rect 374210 472170 374278 472226
rect 374334 472170 374402 472226
rect 374458 472170 374526 472226
rect 374582 472170 374678 472226
rect 374058 472102 374678 472170
rect 374058 472046 374154 472102
rect 374210 472046 374278 472102
rect 374334 472046 374402 472102
rect 374458 472046 374526 472102
rect 374582 472046 374678 472102
rect 374058 471978 374678 472046
rect 374058 471922 374154 471978
rect 374210 471922 374278 471978
rect 374334 471922 374402 471978
rect 374458 471922 374526 471978
rect 374582 471922 374678 471978
rect 351036 471716 351092 471726
rect 351036 468658 351092 471660
rect 351036 468592 351092 468602
rect 371808 460350 372128 460384
rect 371808 460294 371878 460350
rect 371934 460294 372002 460350
rect 372058 460294 372128 460350
rect 371808 460226 372128 460294
rect 371808 460170 371878 460226
rect 371934 460170 372002 460226
rect 372058 460170 372128 460226
rect 371808 460102 372128 460170
rect 371808 460046 371878 460102
rect 371934 460046 372002 460102
rect 372058 460046 372128 460102
rect 371808 459978 372128 460046
rect 371808 459922 371878 459978
rect 371934 459922 372002 459978
rect 372058 459922 372128 459978
rect 371808 459888 372128 459922
rect 354396 458164 354452 458174
rect 354396 456708 354452 458108
rect 354396 456642 354452 456652
rect 354396 456260 354452 456270
rect 354396 450436 354452 456204
rect 354396 450370 354452 450380
rect 374058 454350 374678 471922
rect 374058 454294 374154 454350
rect 374210 454294 374278 454350
rect 374334 454294 374402 454350
rect 374458 454294 374526 454350
rect 374582 454294 374678 454350
rect 374058 454226 374678 454294
rect 374058 454170 374154 454226
rect 374210 454170 374278 454226
rect 374334 454170 374402 454226
rect 374458 454170 374526 454226
rect 374582 454170 374678 454226
rect 374058 454102 374678 454170
rect 374058 454046 374154 454102
rect 374210 454046 374278 454102
rect 374334 454046 374402 454102
rect 374458 454046 374526 454102
rect 374582 454046 374678 454102
rect 374058 453978 374678 454046
rect 374058 453922 374154 453978
rect 374210 453922 374278 453978
rect 374334 453922 374402 453978
rect 374458 453922 374526 453978
rect 374582 453922 374678 453978
rect 348796 446002 348852 446012
rect 351932 449764 351988 449774
rect 348572 421250 348628 421260
rect 348796 421540 348852 421550
rect 347058 406294 347154 406350
rect 347210 406294 347278 406350
rect 347334 406294 347402 406350
rect 347458 406294 347526 406350
rect 347582 406294 347678 406350
rect 347058 406226 347678 406294
rect 347058 406170 347154 406226
rect 347210 406170 347278 406226
rect 347334 406170 347402 406226
rect 347458 406170 347526 406226
rect 347582 406170 347678 406226
rect 347058 406102 347678 406170
rect 347058 406046 347154 406102
rect 347210 406046 347278 406102
rect 347334 406046 347402 406102
rect 347458 406046 347526 406102
rect 347582 406046 347678 406102
rect 347058 405978 347678 406046
rect 347058 405922 347154 405978
rect 347210 405922 347278 405978
rect 347334 405922 347402 405978
rect 347458 405922 347526 405978
rect 347582 405922 347678 405978
rect 343338 400294 343434 400350
rect 343490 400294 343558 400350
rect 343614 400294 343682 400350
rect 343738 400294 343806 400350
rect 343862 400294 343958 400350
rect 343338 400226 343958 400294
rect 343338 400170 343434 400226
rect 343490 400170 343558 400226
rect 343614 400170 343682 400226
rect 343738 400170 343806 400226
rect 343862 400170 343958 400226
rect 343338 400102 343958 400170
rect 343338 400046 343434 400102
rect 343490 400046 343558 400102
rect 343614 400046 343682 400102
rect 343738 400046 343806 400102
rect 343862 400046 343958 400102
rect 343338 399978 343958 400046
rect 343338 399922 343434 399978
rect 343490 399922 343558 399978
rect 343614 399922 343682 399978
rect 343738 399922 343806 399978
rect 343862 399922 343958 399978
rect 343338 382350 343958 399922
rect 343338 382294 343434 382350
rect 343490 382294 343558 382350
rect 343614 382294 343682 382350
rect 343738 382294 343806 382350
rect 343862 382294 343958 382350
rect 343338 382226 343958 382294
rect 343338 382170 343434 382226
rect 343490 382170 343558 382226
rect 343614 382170 343682 382226
rect 343738 382170 343806 382226
rect 343862 382170 343958 382226
rect 343338 382102 343958 382170
rect 343338 382046 343434 382102
rect 343490 382046 343558 382102
rect 343614 382046 343682 382102
rect 343738 382046 343806 382102
rect 343862 382046 343958 382102
rect 343338 381978 343958 382046
rect 343338 381922 343434 381978
rect 343490 381922 343558 381978
rect 343614 381922 343682 381978
rect 343738 381922 343806 381978
rect 343862 381922 343958 381978
rect 343338 364350 343958 381922
rect 343338 364294 343434 364350
rect 343490 364294 343558 364350
rect 343614 364294 343682 364350
rect 343738 364294 343806 364350
rect 343862 364294 343958 364350
rect 343338 364226 343958 364294
rect 343338 364170 343434 364226
rect 343490 364170 343558 364226
rect 343614 364170 343682 364226
rect 343738 364170 343806 364226
rect 343862 364170 343958 364226
rect 343338 364102 343958 364170
rect 343338 364046 343434 364102
rect 343490 364046 343558 364102
rect 343614 364046 343682 364102
rect 343738 364046 343806 364102
rect 343862 364046 343958 364102
rect 343338 363978 343958 364046
rect 343338 363922 343434 363978
rect 343490 363922 343558 363978
rect 343614 363922 343682 363978
rect 343738 363922 343806 363978
rect 343862 363922 343958 363978
rect 338492 357970 338548 357980
rect 335916 357410 335972 357420
rect 334460 350756 334516 350766
rect 334460 349498 334516 350700
rect 334460 349432 334516 349442
rect 343338 346350 343958 363922
rect 345212 402724 345268 402734
rect 345212 360836 345268 402668
rect 345212 360770 345268 360780
rect 347058 388350 347678 405922
rect 347788 409444 347844 409454
rect 347788 403284 347844 409388
rect 347788 403218 347844 403228
rect 348796 399028 348852 421484
rect 350252 420058 350308 420068
rect 350252 401716 350308 420002
rect 351932 416276 351988 449708
rect 352156 449428 352212 449438
rect 352156 430612 352212 449372
rect 355292 447748 355348 447758
rect 352156 430546 352212 430556
rect 353612 446404 353668 446414
rect 353612 425796 353668 446348
rect 355292 435876 355348 447692
rect 355292 435810 355348 435820
rect 370412 446180 370468 446190
rect 370412 429716 370468 446124
rect 370412 429650 370468 429660
rect 374058 436350 374678 453922
rect 374058 436294 374154 436350
rect 374210 436294 374278 436350
rect 374334 436294 374402 436350
rect 374458 436294 374526 436350
rect 374582 436294 374678 436350
rect 374058 436226 374678 436294
rect 374058 436170 374154 436226
rect 374210 436170 374278 436226
rect 374334 436170 374402 436226
rect 374458 436170 374526 436226
rect 374582 436170 374678 436226
rect 374058 436102 374678 436170
rect 374058 436046 374154 436102
rect 374210 436046 374278 436102
rect 374334 436046 374402 436102
rect 374458 436046 374526 436102
rect 374582 436046 374678 436102
rect 374058 435978 374678 436046
rect 374058 435922 374154 435978
rect 374210 435922 374278 435978
rect 374334 435922 374402 435978
rect 374458 435922 374526 435978
rect 374582 435922 374678 435978
rect 353612 425730 353668 425740
rect 356448 418350 356768 418384
rect 356448 418294 356518 418350
rect 356574 418294 356642 418350
rect 356698 418294 356768 418350
rect 356448 418226 356768 418294
rect 356448 418170 356518 418226
rect 356574 418170 356642 418226
rect 356698 418170 356768 418226
rect 356448 418102 356768 418170
rect 356448 418046 356518 418102
rect 356574 418046 356642 418102
rect 356698 418046 356768 418102
rect 356448 417978 356768 418046
rect 356448 417922 356518 417978
rect 356574 417922 356642 417978
rect 356698 417922 356768 417978
rect 356448 417888 356768 417922
rect 374058 418350 374678 435922
rect 374058 418294 374154 418350
rect 374210 418294 374278 418350
rect 374334 418294 374402 418350
rect 374458 418294 374526 418350
rect 374582 418294 374678 418350
rect 374058 418226 374678 418294
rect 374058 418170 374154 418226
rect 374210 418170 374278 418226
rect 374334 418170 374402 418226
rect 374458 418170 374526 418226
rect 374582 418170 374678 418226
rect 374058 418102 374678 418170
rect 374058 418046 374154 418102
rect 374210 418046 374278 418102
rect 374334 418046 374402 418102
rect 374458 418046 374526 418102
rect 374582 418046 374678 418102
rect 374058 417978 374678 418046
rect 374058 417922 374154 417978
rect 374210 417922 374278 417978
rect 374334 417922 374402 417978
rect 374458 417922 374526 417978
rect 374582 417922 374678 417978
rect 351932 416210 351988 416220
rect 351036 412916 351092 412926
rect 351036 409798 351092 412860
rect 352716 411598 352772 411608
rect 352716 411460 352772 411542
rect 352716 411394 352772 411404
rect 351036 409732 351092 409742
rect 350252 401650 350308 401660
rect 350364 409108 350420 409118
rect 348796 398962 348852 398972
rect 350364 391438 350420 409052
rect 371808 406350 372128 406384
rect 371808 406294 371878 406350
rect 371934 406294 372002 406350
rect 372058 406294 372128 406350
rect 371808 406226 372128 406294
rect 371808 406170 371878 406226
rect 371934 406170 372002 406226
rect 372058 406170 372128 406226
rect 371808 406102 372128 406170
rect 371808 406046 371878 406102
rect 371934 406046 372002 406102
rect 372058 406046 372128 406102
rect 371808 405978 372128 406046
rect 371808 405922 371878 405978
rect 371934 405922 372002 405978
rect 372058 405922 372128 405978
rect 371808 405888 372128 405922
rect 374058 404318 374678 417922
rect 377778 598172 378398 598268
rect 377778 598116 377874 598172
rect 377930 598116 377998 598172
rect 378054 598116 378122 598172
rect 378178 598116 378246 598172
rect 378302 598116 378398 598172
rect 377778 598048 378398 598116
rect 377778 597992 377874 598048
rect 377930 597992 377998 598048
rect 378054 597992 378122 598048
rect 378178 597992 378246 598048
rect 378302 597992 378398 598048
rect 377778 597924 378398 597992
rect 377778 597868 377874 597924
rect 377930 597868 377998 597924
rect 378054 597868 378122 597924
rect 378178 597868 378246 597924
rect 378302 597868 378398 597924
rect 377778 597800 378398 597868
rect 377778 597744 377874 597800
rect 377930 597744 377998 597800
rect 378054 597744 378122 597800
rect 378178 597744 378246 597800
rect 378302 597744 378398 597800
rect 377778 586350 378398 597744
rect 377778 586294 377874 586350
rect 377930 586294 377998 586350
rect 378054 586294 378122 586350
rect 378178 586294 378246 586350
rect 378302 586294 378398 586350
rect 377778 586226 378398 586294
rect 377778 586170 377874 586226
rect 377930 586170 377998 586226
rect 378054 586170 378122 586226
rect 378178 586170 378246 586226
rect 378302 586170 378398 586226
rect 377778 586102 378398 586170
rect 377778 586046 377874 586102
rect 377930 586046 377998 586102
rect 378054 586046 378122 586102
rect 378178 586046 378246 586102
rect 378302 586046 378398 586102
rect 377778 585978 378398 586046
rect 377778 585922 377874 585978
rect 377930 585922 377998 585978
rect 378054 585922 378122 585978
rect 378178 585922 378246 585978
rect 378302 585922 378398 585978
rect 377778 568350 378398 585922
rect 377778 568294 377874 568350
rect 377930 568294 377998 568350
rect 378054 568294 378122 568350
rect 378178 568294 378246 568350
rect 378302 568294 378398 568350
rect 377778 568226 378398 568294
rect 377778 568170 377874 568226
rect 377930 568170 377998 568226
rect 378054 568170 378122 568226
rect 378178 568170 378246 568226
rect 378302 568170 378398 568226
rect 377778 568102 378398 568170
rect 377778 568046 377874 568102
rect 377930 568046 377998 568102
rect 378054 568046 378122 568102
rect 378178 568046 378246 568102
rect 378302 568046 378398 568102
rect 377778 567978 378398 568046
rect 377778 567922 377874 567978
rect 377930 567922 377998 567978
rect 378054 567922 378122 567978
rect 378178 567922 378246 567978
rect 378302 567922 378398 567978
rect 377778 550350 378398 567922
rect 404778 597212 405398 598268
rect 404778 597156 404874 597212
rect 404930 597156 404998 597212
rect 405054 597156 405122 597212
rect 405178 597156 405246 597212
rect 405302 597156 405398 597212
rect 404778 597088 405398 597156
rect 404778 597032 404874 597088
rect 404930 597032 404998 597088
rect 405054 597032 405122 597088
rect 405178 597032 405246 597088
rect 405302 597032 405398 597088
rect 404778 596964 405398 597032
rect 404778 596908 404874 596964
rect 404930 596908 404998 596964
rect 405054 596908 405122 596964
rect 405178 596908 405246 596964
rect 405302 596908 405398 596964
rect 404778 596840 405398 596908
rect 404778 596784 404874 596840
rect 404930 596784 404998 596840
rect 405054 596784 405122 596840
rect 405178 596784 405246 596840
rect 405302 596784 405398 596840
rect 404778 580350 405398 596784
rect 404778 580294 404874 580350
rect 404930 580294 404998 580350
rect 405054 580294 405122 580350
rect 405178 580294 405246 580350
rect 405302 580294 405398 580350
rect 404778 580226 405398 580294
rect 404778 580170 404874 580226
rect 404930 580170 404998 580226
rect 405054 580170 405122 580226
rect 405178 580170 405246 580226
rect 405302 580170 405398 580226
rect 404778 580102 405398 580170
rect 404778 580046 404874 580102
rect 404930 580046 404998 580102
rect 405054 580046 405122 580102
rect 405178 580046 405246 580102
rect 405302 580046 405398 580102
rect 404778 579978 405398 580046
rect 404778 579922 404874 579978
rect 404930 579922 404998 579978
rect 405054 579922 405122 579978
rect 405178 579922 405246 579978
rect 405302 579922 405398 579978
rect 387168 562350 387488 562384
rect 387168 562294 387238 562350
rect 387294 562294 387362 562350
rect 387418 562294 387488 562350
rect 387168 562226 387488 562294
rect 387168 562170 387238 562226
rect 387294 562170 387362 562226
rect 387418 562170 387488 562226
rect 387168 562102 387488 562170
rect 387168 562046 387238 562102
rect 387294 562046 387362 562102
rect 387418 562046 387488 562102
rect 387168 561978 387488 562046
rect 387168 561922 387238 561978
rect 387294 561922 387362 561978
rect 387418 561922 387488 561978
rect 387168 561888 387488 561922
rect 404778 562350 405398 579922
rect 404778 562294 404874 562350
rect 404930 562294 404998 562350
rect 405054 562294 405122 562350
rect 405178 562294 405246 562350
rect 405302 562294 405398 562350
rect 404778 562226 405398 562294
rect 404778 562170 404874 562226
rect 404930 562170 404998 562226
rect 405054 562170 405122 562226
rect 405178 562170 405246 562226
rect 405302 562170 405398 562226
rect 404778 562102 405398 562170
rect 404778 562046 404874 562102
rect 404930 562046 404998 562102
rect 405054 562046 405122 562102
rect 405178 562046 405246 562102
rect 405302 562046 405398 562102
rect 404778 561978 405398 562046
rect 404778 561922 404874 561978
rect 404930 561922 404998 561978
rect 405054 561922 405122 561978
rect 405178 561922 405246 561978
rect 405302 561922 405398 561978
rect 396844 551908 396900 551918
rect 377778 550294 377874 550350
rect 377930 550294 377998 550350
rect 378054 550294 378122 550350
rect 378178 550294 378246 550350
rect 378302 550294 378398 550350
rect 377778 550226 378398 550294
rect 377778 550170 377874 550226
rect 377930 550170 377998 550226
rect 378054 550170 378122 550226
rect 378178 550170 378246 550226
rect 378302 550170 378398 550226
rect 377778 550102 378398 550170
rect 377778 550046 377874 550102
rect 377930 550046 377998 550102
rect 378054 550046 378122 550102
rect 378178 550046 378246 550102
rect 378302 550046 378398 550102
rect 377778 549978 378398 550046
rect 377778 549922 377874 549978
rect 377930 549922 377998 549978
rect 378054 549922 378122 549978
rect 378178 549922 378246 549978
rect 378302 549922 378398 549978
rect 377778 532350 378398 549922
rect 394828 551236 394884 551246
rect 393372 547204 393428 547214
rect 387168 544350 387488 544384
rect 387168 544294 387238 544350
rect 387294 544294 387362 544350
rect 387418 544294 387488 544350
rect 387168 544226 387488 544294
rect 387168 544170 387238 544226
rect 387294 544170 387362 544226
rect 387418 544170 387488 544226
rect 387168 544102 387488 544170
rect 387168 544046 387238 544102
rect 387294 544046 387362 544102
rect 387418 544046 387488 544102
rect 387168 543978 387488 544046
rect 387168 543922 387238 543978
rect 387294 543922 387362 543978
rect 387418 543922 387488 543978
rect 387168 543888 387488 543922
rect 377778 532294 377874 532350
rect 377930 532294 377998 532350
rect 378054 532294 378122 532350
rect 378178 532294 378246 532350
rect 378302 532294 378398 532350
rect 377778 532226 378398 532294
rect 377778 532170 377874 532226
rect 377930 532170 377998 532226
rect 378054 532170 378122 532226
rect 378178 532170 378246 532226
rect 378302 532170 378398 532226
rect 377778 532102 378398 532170
rect 377778 532046 377874 532102
rect 377930 532046 377998 532102
rect 378054 532046 378122 532102
rect 378178 532046 378246 532102
rect 378302 532046 378398 532102
rect 377778 531978 378398 532046
rect 377778 531922 377874 531978
rect 377930 531922 377998 531978
rect 378054 531922 378122 531978
rect 378178 531922 378246 531978
rect 378302 531922 378398 531978
rect 377778 514350 378398 531922
rect 377778 514294 377874 514350
rect 377930 514294 377998 514350
rect 378054 514294 378122 514350
rect 378178 514294 378246 514350
rect 378302 514294 378398 514350
rect 377778 514226 378398 514294
rect 377778 514170 377874 514226
rect 377930 514170 377998 514226
rect 378054 514170 378122 514226
rect 378178 514170 378246 514226
rect 378302 514170 378398 514226
rect 377778 514102 378398 514170
rect 377778 514046 377874 514102
rect 377930 514046 377998 514102
rect 378054 514046 378122 514102
rect 378178 514046 378246 514102
rect 378302 514046 378398 514102
rect 377778 513978 378398 514046
rect 377778 513922 377874 513978
rect 377930 513922 377998 513978
rect 378054 513922 378122 513978
rect 378178 513922 378246 513978
rect 378302 513922 378398 513978
rect 377778 496350 378398 513922
rect 380492 520100 380548 520110
rect 380492 513716 380548 520044
rect 380492 513650 380548 513660
rect 393372 506660 393428 547148
rect 394828 510244 394884 551180
rect 394828 510178 394884 510188
rect 394940 544516 394996 544526
rect 393372 506594 393428 506604
rect 394940 504868 394996 544460
rect 394940 504802 394996 504812
rect 395612 543284 395668 543294
rect 377778 496294 377874 496350
rect 377930 496294 377998 496350
rect 378054 496294 378122 496350
rect 378178 496294 378246 496350
rect 378302 496294 378398 496350
rect 377778 496226 378398 496294
rect 377778 496170 377874 496226
rect 377930 496170 377998 496226
rect 378054 496170 378122 496226
rect 378178 496170 378246 496226
rect 378302 496170 378398 496226
rect 377778 496102 378398 496170
rect 377778 496046 377874 496102
rect 377930 496046 377998 496102
rect 378054 496046 378122 496102
rect 378178 496046 378246 496102
rect 378302 496046 378398 496102
rect 377778 495978 378398 496046
rect 377778 495922 377874 495978
rect 377930 495922 377998 495978
rect 378054 495922 378122 495978
rect 378178 495922 378246 495978
rect 378302 495922 378398 495978
rect 377778 478350 378398 495922
rect 393932 503188 393988 503198
rect 393932 495796 393988 503132
rect 395612 503076 395668 543228
rect 396732 542724 396788 542734
rect 396620 542500 396676 542510
rect 396620 505428 396676 542444
rect 396732 522004 396788 542668
rect 396732 521938 396788 521948
rect 396620 505362 396676 505372
rect 396844 503524 396900 551852
rect 402332 548548 402388 548558
rect 398972 543844 399028 543854
rect 398972 515956 399028 543788
rect 398972 515890 399028 515900
rect 402332 511924 402388 548492
rect 402332 511858 402388 511868
rect 404778 544350 405398 561922
rect 404778 544294 404874 544350
rect 404930 544294 404998 544350
rect 405054 544294 405122 544350
rect 405178 544294 405246 544350
rect 405302 544294 405398 544350
rect 404778 544226 405398 544294
rect 404778 544170 404874 544226
rect 404930 544170 404998 544226
rect 405054 544170 405122 544226
rect 405178 544170 405246 544226
rect 405302 544170 405398 544226
rect 404778 544102 405398 544170
rect 404778 544046 404874 544102
rect 404930 544046 404998 544102
rect 405054 544046 405122 544102
rect 405178 544046 405246 544102
rect 405302 544046 405398 544102
rect 404778 543978 405398 544046
rect 404778 543922 404874 543978
rect 404930 543922 404998 543978
rect 405054 543922 405122 543978
rect 405178 543922 405246 543978
rect 405302 543922 405398 543978
rect 404778 526350 405398 543922
rect 404778 526294 404874 526350
rect 404930 526294 404998 526350
rect 405054 526294 405122 526350
rect 405178 526294 405246 526350
rect 405302 526294 405398 526350
rect 404778 526226 405398 526294
rect 404778 526170 404874 526226
rect 404930 526170 404998 526226
rect 405054 526170 405122 526226
rect 405178 526170 405246 526226
rect 405302 526170 405398 526226
rect 404778 526102 405398 526170
rect 404778 526046 404874 526102
rect 404930 526046 404998 526102
rect 405054 526046 405122 526102
rect 405178 526046 405246 526102
rect 405302 526046 405398 526102
rect 404778 525978 405398 526046
rect 404778 525922 404874 525978
rect 404930 525922 404998 525978
rect 405054 525922 405122 525978
rect 405178 525922 405246 525978
rect 405302 525922 405398 525978
rect 404778 508350 405398 525922
rect 404778 508294 404874 508350
rect 404930 508294 404998 508350
rect 405054 508294 405122 508350
rect 405178 508294 405246 508350
rect 405302 508294 405398 508350
rect 404778 508226 405398 508294
rect 404778 508170 404874 508226
rect 404930 508170 404998 508226
rect 405054 508170 405122 508226
rect 405178 508170 405246 508226
rect 405302 508170 405398 508226
rect 404778 508102 405398 508170
rect 404778 508046 404874 508102
rect 404930 508046 404998 508102
rect 405054 508046 405122 508102
rect 405178 508046 405246 508102
rect 405302 508046 405398 508102
rect 404778 507978 405398 508046
rect 404778 507922 404874 507978
rect 404930 507922 404998 507978
rect 405054 507922 405122 507978
rect 405178 507922 405246 507978
rect 405302 507922 405398 507978
rect 396844 503458 396900 503468
rect 402332 506660 402388 506670
rect 395612 503010 395668 503020
rect 402332 496916 402388 506604
rect 402332 496850 402388 496860
rect 393932 495730 393988 495740
rect 387168 490350 387488 490384
rect 387168 490294 387238 490350
rect 387294 490294 387362 490350
rect 387418 490294 387488 490350
rect 387168 490226 387488 490294
rect 387168 490170 387238 490226
rect 387294 490170 387362 490226
rect 387418 490170 387488 490226
rect 387168 490102 387488 490170
rect 387168 490046 387238 490102
rect 387294 490046 387362 490102
rect 387418 490046 387488 490102
rect 387168 489978 387488 490046
rect 387168 489922 387238 489978
rect 387294 489922 387362 489978
rect 387418 489922 387488 489978
rect 387168 489888 387488 489922
rect 404778 490350 405398 507922
rect 404778 490294 404874 490350
rect 404930 490294 404998 490350
rect 405054 490294 405122 490350
rect 405178 490294 405246 490350
rect 405302 490294 405398 490350
rect 404778 490226 405398 490294
rect 404778 490170 404874 490226
rect 404930 490170 404998 490226
rect 405054 490170 405122 490226
rect 405178 490170 405246 490226
rect 405302 490170 405398 490226
rect 404778 490102 405398 490170
rect 404778 490046 404874 490102
rect 404930 490046 404998 490102
rect 405054 490046 405122 490102
rect 405178 490046 405246 490102
rect 405302 490046 405398 490102
rect 404778 489978 405398 490046
rect 404778 489922 404874 489978
rect 404930 489922 404998 489978
rect 405054 489922 405122 489978
rect 405178 489922 405246 489978
rect 405302 489922 405398 489978
rect 396844 483364 396900 483374
rect 396732 482692 396788 482702
rect 377778 478294 377874 478350
rect 377930 478294 377998 478350
rect 378054 478294 378122 478350
rect 378178 478294 378246 478350
rect 378302 478294 378398 478350
rect 377778 478226 378398 478294
rect 377778 478170 377874 478226
rect 377930 478170 377998 478226
rect 378054 478170 378122 478226
rect 378178 478170 378246 478226
rect 378302 478170 378398 478226
rect 377778 478102 378398 478170
rect 377778 478046 377874 478102
rect 377930 478046 377998 478102
rect 378054 478046 378122 478102
rect 378178 478046 378246 478102
rect 378302 478046 378398 478102
rect 377778 477978 378398 478046
rect 377778 477922 377874 477978
rect 377930 477922 377998 477978
rect 378054 477922 378122 477978
rect 378178 477922 378246 477978
rect 378302 477922 378398 477978
rect 377778 460350 378398 477922
rect 394828 480004 394884 480014
rect 393372 475972 393428 475982
rect 387168 472350 387488 472384
rect 387168 472294 387238 472350
rect 387294 472294 387362 472350
rect 387418 472294 387488 472350
rect 387168 472226 387488 472294
rect 387168 472170 387238 472226
rect 387294 472170 387362 472226
rect 387418 472170 387488 472226
rect 387168 472102 387488 472170
rect 387168 472046 387238 472102
rect 387294 472046 387362 472102
rect 387418 472046 387488 472102
rect 387168 471978 387488 472046
rect 387168 471922 387238 471978
rect 387294 471922 387362 471978
rect 387418 471922 387488 471978
rect 387168 471888 387488 471922
rect 377778 460294 377874 460350
rect 377930 460294 377998 460350
rect 378054 460294 378122 460350
rect 378178 460294 378246 460350
rect 378302 460294 378398 460350
rect 377778 460226 378398 460294
rect 377778 460170 377874 460226
rect 377930 460170 377998 460226
rect 378054 460170 378122 460226
rect 378178 460170 378246 460226
rect 378302 460170 378398 460226
rect 377778 460102 378398 460170
rect 377778 460046 377874 460102
rect 377930 460046 377998 460102
rect 378054 460046 378122 460102
rect 378178 460046 378246 460102
rect 378302 460046 378398 460102
rect 377778 459978 378398 460046
rect 377778 459922 377874 459978
rect 377930 459922 377998 459978
rect 378054 459922 378122 459978
rect 378178 459922 378246 459978
rect 378302 459922 378398 459978
rect 377778 442350 378398 459922
rect 392476 457156 392532 457166
rect 392364 449540 392420 449550
rect 377778 442294 377874 442350
rect 377930 442294 377998 442350
rect 378054 442294 378122 442350
rect 378178 442294 378246 442350
rect 378302 442294 378398 442350
rect 377778 442226 378398 442294
rect 377778 442170 377874 442226
rect 377930 442170 377998 442226
rect 378054 442170 378122 442226
rect 378178 442170 378246 442226
rect 378302 442170 378398 442226
rect 377778 442102 378398 442170
rect 377778 442046 377874 442102
rect 377930 442046 377998 442102
rect 378054 442046 378122 442102
rect 378178 442046 378246 442102
rect 378302 442046 378398 442102
rect 377778 441978 378398 442046
rect 377778 441922 377874 441978
rect 377930 441922 377998 441978
rect 378054 441922 378122 441978
rect 378178 441922 378246 441978
rect 378302 441922 378398 441978
rect 377778 424350 378398 441922
rect 391356 446068 391412 446078
rect 391356 440356 391412 446012
rect 391356 440290 391412 440300
rect 392364 439796 392420 449484
rect 392476 447636 392532 457100
rect 393372 451220 393428 475916
rect 393372 451154 393428 451164
rect 392476 447570 392532 447580
rect 392364 439730 392420 439740
rect 394828 437668 394884 479948
rect 394940 479332 394996 479342
rect 394940 444724 394996 479276
rect 396508 478660 396564 478670
rect 395612 475412 395668 475422
rect 395052 471940 395108 471950
rect 395052 449316 395108 471884
rect 395052 449250 395108 449260
rect 395612 447076 395668 475356
rect 395612 447010 395668 447020
rect 396508 446628 396564 478604
rect 396620 476644 396676 476654
rect 396620 449764 396676 476588
rect 396732 457156 396788 482636
rect 396844 475412 396900 483308
rect 404012 477988 404068 477998
rect 396844 475346 396900 475356
rect 400652 475972 400708 475982
rect 396732 457090 396788 457100
rect 396844 473284 396900 473294
rect 396620 449698 396676 449708
rect 396844 449652 396900 473228
rect 398972 462868 399028 462878
rect 398972 450996 399028 462812
rect 398972 450930 399028 450940
rect 396844 449586 396900 449596
rect 396508 446562 396564 446572
rect 394940 444658 394996 444668
rect 394828 437602 394884 437612
rect 400652 426692 400708 475916
rect 402332 473956 402388 473966
rect 402332 428036 402388 473900
rect 404012 428596 404068 477932
rect 404012 428530 404068 428540
rect 404778 472350 405398 489922
rect 404778 472294 404874 472350
rect 404930 472294 404998 472350
rect 405054 472294 405122 472350
rect 405178 472294 405246 472350
rect 405302 472294 405398 472350
rect 404778 472226 405398 472294
rect 404778 472170 404874 472226
rect 404930 472170 404998 472226
rect 405054 472170 405122 472226
rect 405178 472170 405246 472226
rect 405302 472170 405398 472226
rect 404778 472102 405398 472170
rect 404778 472046 404874 472102
rect 404930 472046 404998 472102
rect 405054 472046 405122 472102
rect 405178 472046 405246 472102
rect 405302 472046 405398 472102
rect 404778 471978 405398 472046
rect 404778 471922 404874 471978
rect 404930 471922 404998 471978
rect 405054 471922 405122 471978
rect 405178 471922 405246 471978
rect 405302 471922 405398 471978
rect 404778 454350 405398 471922
rect 404778 454294 404874 454350
rect 404930 454294 404998 454350
rect 405054 454294 405122 454350
rect 405178 454294 405246 454350
rect 405302 454294 405398 454350
rect 404778 454226 405398 454294
rect 404778 454170 404874 454226
rect 404930 454170 404998 454226
rect 405054 454170 405122 454226
rect 405178 454170 405246 454226
rect 405302 454170 405398 454226
rect 404778 454102 405398 454170
rect 404778 454046 404874 454102
rect 404930 454046 404998 454102
rect 405054 454046 405122 454102
rect 405178 454046 405246 454102
rect 405302 454046 405398 454102
rect 404778 453978 405398 454046
rect 404778 453922 404874 453978
rect 404930 453922 404998 453978
rect 405054 453922 405122 453978
rect 405178 453922 405246 453978
rect 405302 453922 405398 453978
rect 404778 436350 405398 453922
rect 404778 436294 404874 436350
rect 404930 436294 404998 436350
rect 405054 436294 405122 436350
rect 405178 436294 405246 436350
rect 405302 436294 405398 436350
rect 404778 436226 405398 436294
rect 404778 436170 404874 436226
rect 404930 436170 404998 436226
rect 405054 436170 405122 436226
rect 405178 436170 405246 436226
rect 405302 436170 405398 436226
rect 404778 436102 405398 436170
rect 404778 436046 404874 436102
rect 404930 436046 404998 436102
rect 405054 436046 405122 436102
rect 405178 436046 405246 436102
rect 405302 436046 405398 436102
rect 404778 435978 405398 436046
rect 404778 435922 404874 435978
rect 404930 435922 404998 435978
rect 405054 435922 405122 435978
rect 405178 435922 405246 435978
rect 405302 435922 405398 435978
rect 402332 427970 402388 427980
rect 400652 426626 400708 426636
rect 377778 424294 377874 424350
rect 377930 424294 377998 424350
rect 378054 424294 378122 424350
rect 378178 424294 378246 424350
rect 378302 424294 378398 424350
rect 377778 424226 378398 424294
rect 377778 424170 377874 424226
rect 377930 424170 377998 424226
rect 378054 424170 378122 424226
rect 378178 424170 378246 424226
rect 378302 424170 378398 424226
rect 377778 424102 378398 424170
rect 377778 424046 377874 424102
rect 377930 424046 377998 424102
rect 378054 424046 378122 424102
rect 378178 424046 378246 424102
rect 378302 424046 378398 424102
rect 377778 423978 378398 424046
rect 377778 423922 377874 423978
rect 377930 423922 377998 423978
rect 378054 423922 378122 423978
rect 378178 423922 378246 423978
rect 378302 423922 378398 423978
rect 377778 406350 378398 423922
rect 396620 421540 396676 421550
rect 395612 419972 395668 419982
rect 387168 418350 387488 418384
rect 387168 418294 387238 418350
rect 387294 418294 387362 418350
rect 387418 418294 387488 418350
rect 387168 418226 387488 418294
rect 387168 418170 387238 418226
rect 387294 418170 387362 418226
rect 387418 418170 387488 418226
rect 387168 418102 387488 418170
rect 387168 418046 387238 418102
rect 387294 418046 387362 418102
rect 387418 418046 387488 418102
rect 387168 417978 387488 418046
rect 387168 417922 387238 417978
rect 387294 417922 387362 417978
rect 387418 417922 387488 417978
rect 387168 417888 387488 417922
rect 377778 406294 377874 406350
rect 377930 406294 377998 406350
rect 378054 406294 378122 406350
rect 378178 406294 378246 406350
rect 378302 406294 378398 406350
rect 377778 406226 378398 406294
rect 377778 406170 377874 406226
rect 377930 406170 377998 406226
rect 378054 406170 378122 406226
rect 378178 406170 378246 406226
rect 378302 406170 378398 406226
rect 377778 406102 378398 406170
rect 377778 406046 377874 406102
rect 377930 406046 377998 406102
rect 378054 406046 378122 406102
rect 378178 406046 378246 406102
rect 378302 406046 378398 406102
rect 377778 405978 378398 406046
rect 377778 405922 377874 405978
rect 377930 405922 377998 405978
rect 378054 405922 378122 405978
rect 378178 405922 378246 405978
rect 378302 405922 378398 405978
rect 351036 402418 351092 402428
rect 351036 398356 351092 402362
rect 356448 400350 356768 400384
rect 356448 400294 356518 400350
rect 356574 400294 356642 400350
rect 356698 400294 356768 400350
rect 356448 400226 356768 400294
rect 356448 400170 356518 400226
rect 356574 400170 356642 400226
rect 356698 400170 356768 400226
rect 356448 400102 356768 400170
rect 356448 400046 356518 400102
rect 356574 400046 356642 400102
rect 356698 400046 356768 400102
rect 356448 399978 356768 400046
rect 356448 399922 356518 399978
rect 356574 399922 356642 399978
rect 356698 399922 356768 399978
rect 356448 399888 356768 399922
rect 351036 398290 351092 398300
rect 350364 391372 350420 391382
rect 347058 388294 347154 388350
rect 347210 388294 347278 388350
rect 347334 388294 347402 388350
rect 347458 388294 347526 388350
rect 347582 388294 347678 388350
rect 347058 388226 347678 388294
rect 371808 388389 372128 388446
rect 371808 388333 371836 388389
rect 371892 388333 371940 388389
rect 371996 388333 372044 388389
rect 372100 388333 372128 388389
rect 371808 388276 372128 388333
rect 347058 388170 347154 388226
rect 347210 388170 347278 388226
rect 347334 388170 347402 388226
rect 347458 388170 347526 388226
rect 347582 388170 347678 388226
rect 347058 388102 347678 388170
rect 347058 388046 347154 388102
rect 347210 388046 347278 388102
rect 347334 388046 347402 388102
rect 347458 388046 347526 388102
rect 347582 388046 347678 388102
rect 347058 387978 347678 388046
rect 347058 387922 347154 387978
rect 347210 387922 347278 387978
rect 347334 387922 347402 387978
rect 347458 387922 347526 387978
rect 347582 387922 347678 387978
rect 347058 370350 347678 387922
rect 349468 387716 349524 387726
rect 347788 387268 347844 387278
rect 347788 383236 347844 387212
rect 349468 384580 349524 387660
rect 371308 385700 371364 385710
rect 367052 385364 367108 385374
rect 367052 385028 367108 385308
rect 367052 384962 367108 384972
rect 349468 384514 349524 384524
rect 347788 383170 347844 383180
rect 371308 381556 371364 385644
rect 371308 381490 371364 381500
rect 374058 382350 374678 399570
rect 374058 382294 374154 382350
rect 374210 382294 374278 382350
rect 374334 382294 374402 382350
rect 374458 382294 374526 382350
rect 374582 382294 374678 382350
rect 374058 382226 374678 382294
rect 374058 382170 374154 382226
rect 374210 382170 374278 382226
rect 374334 382170 374402 382226
rect 374458 382170 374526 382226
rect 374582 382170 374678 382226
rect 374058 382102 374678 382170
rect 374058 382046 374154 382102
rect 374210 382046 374278 382102
rect 374334 382046 374402 382102
rect 374458 382046 374526 382102
rect 374582 382046 374678 382102
rect 374058 381978 374678 382046
rect 374058 381922 374154 381978
rect 374210 381922 374278 381978
rect 374334 381922 374402 381978
rect 374458 381922 374526 381978
rect 374582 381922 374678 381978
rect 347058 370294 347154 370350
rect 347210 370294 347278 370350
rect 347334 370294 347402 370350
rect 347458 370294 347526 370350
rect 347582 370294 347678 370350
rect 347058 370226 347678 370294
rect 347058 370170 347154 370226
rect 347210 370170 347278 370226
rect 347334 370170 347402 370226
rect 347458 370170 347526 370226
rect 347582 370170 347678 370226
rect 347058 370102 347678 370170
rect 347058 370046 347154 370102
rect 347210 370046 347278 370102
rect 347334 370046 347402 370102
rect 347458 370046 347526 370102
rect 347582 370046 347678 370102
rect 347058 369978 347678 370046
rect 347058 369922 347154 369978
rect 347210 369922 347278 369978
rect 347334 369922 347402 369978
rect 347458 369922 347526 369978
rect 347582 369922 347678 369978
rect 343338 346294 343434 346350
rect 343490 346294 343558 346350
rect 343614 346294 343682 346350
rect 343738 346294 343806 346350
rect 343862 346294 343958 346350
rect 343338 346226 343958 346294
rect 343338 346170 343434 346226
rect 343490 346170 343558 346226
rect 343614 346170 343682 346226
rect 343738 346170 343806 346226
rect 343862 346170 343958 346226
rect 343338 346102 343958 346170
rect 343338 346046 343434 346102
rect 343490 346046 343558 346102
rect 343614 346046 343682 346102
rect 343738 346046 343806 346102
rect 343862 346046 343958 346102
rect 343338 345978 343958 346046
rect 343338 345922 343434 345978
rect 343490 345922 343558 345978
rect 343614 345922 343682 345978
rect 343738 345922 343806 345978
rect 343862 345922 343958 345978
rect 334460 345716 334516 345726
rect 334348 345156 334404 345166
rect 334348 343558 334404 345100
rect 334460 344458 334516 345660
rect 334460 344392 334516 344402
rect 334348 343492 334404 343502
rect 334460 344278 334516 344288
rect 334460 343476 334516 344222
rect 334460 343410 334516 343420
rect 334348 342356 334404 342366
rect 334348 341398 334404 342300
rect 334348 341332 334404 341342
rect 334460 341578 334516 341588
rect 334460 341236 334516 341522
rect 334460 341170 334516 341180
rect 334348 340676 334404 340686
rect 334348 339418 334404 340620
rect 334460 340116 334516 340126
rect 334460 339778 334516 340060
rect 334460 339712 334516 339722
rect 334460 339418 334516 339428
rect 334348 339362 334460 339418
rect 334460 339352 334516 339362
rect 334348 338996 334404 339006
rect 334348 337978 334404 338940
rect 341852 338996 341908 339006
rect 338604 338698 338660 338708
rect 334348 337912 334404 337922
rect 337708 338436 337764 338446
rect 334460 337876 334516 337886
rect 334460 337798 334516 337820
rect 334460 337732 334516 337742
rect 334460 337618 334516 337628
rect 334348 337316 334404 337326
rect 334348 336178 334404 337260
rect 334460 336756 334516 337562
rect 334460 336690 334516 336700
rect 334460 336358 334516 336368
rect 334460 336196 334516 336302
rect 334460 336130 334516 336140
rect 334348 336112 334404 336122
rect 334460 335998 334516 336008
rect 334460 335076 334516 335942
rect 334460 335010 334516 335020
rect 334460 334738 334516 334748
rect 334460 334516 334516 334682
rect 334460 334450 334516 334460
rect 334460 333658 334516 333668
rect 334460 333396 334516 333602
rect 334460 333330 334516 333340
rect 334460 332578 334516 332588
rect 334460 331716 334516 332522
rect 334460 331650 334516 331660
rect 337708 330958 337764 338380
rect 337708 330892 337764 330902
rect 334460 330778 334516 330788
rect 334460 330036 334516 330722
rect 334460 329970 334516 329980
rect 338492 330260 338548 330270
rect 334460 329338 334516 329348
rect 334460 327796 334516 329282
rect 334460 327730 334516 327740
rect 334460 327538 334516 327548
rect 334348 327482 334460 327538
rect 334348 326116 334404 327482
rect 334460 327472 334516 327482
rect 334460 327358 334516 327368
rect 334460 327236 334516 327302
rect 334460 327170 334516 327180
rect 334348 326050 334404 326060
rect 334460 325918 334516 325928
rect 334460 324436 334516 325862
rect 334460 324370 334516 324380
rect 334460 324118 334516 324128
rect 334348 323938 334404 323948
rect 334348 322756 334404 323882
rect 334460 323876 334516 324062
rect 334460 323810 334516 323820
rect 334348 322690 334404 322700
rect 334460 322498 334516 322508
rect 334460 321636 334516 322442
rect 334460 321570 334516 321580
rect 334460 320878 334516 320888
rect 334460 319956 334516 320822
rect 334460 319890 334516 319900
rect 334460 319078 334516 319088
rect 334460 318836 334516 319022
rect 334460 318770 334516 318780
rect 338492 299796 338548 330204
rect 338604 328916 338660 338642
rect 338604 328850 338660 328860
rect 341852 300916 341908 338940
rect 341852 300850 341908 300860
rect 343338 328350 343958 345922
rect 347058 352350 347678 369922
rect 374058 364350 374678 381922
rect 374058 364294 374154 364350
rect 374210 364294 374278 364350
rect 374334 364294 374402 364350
rect 374458 364294 374526 364350
rect 374582 364294 374678 364350
rect 374058 364226 374678 364294
rect 374058 364170 374154 364226
rect 374210 364170 374278 364226
rect 374334 364170 374402 364226
rect 374458 364170 374526 364226
rect 374582 364170 374678 364226
rect 374058 364102 374678 364170
rect 374058 364046 374154 364102
rect 374210 364046 374278 364102
rect 374334 364046 374402 364102
rect 374458 364046 374526 364102
rect 374582 364046 374678 364102
rect 374058 363978 374678 364046
rect 374058 363922 374154 363978
rect 374210 363922 374278 363978
rect 374334 363922 374402 363978
rect 374458 363922 374526 363978
rect 374582 363922 374678 363978
rect 351036 353108 351092 353118
rect 351036 352436 351092 353052
rect 351036 352370 351092 352380
rect 352604 352884 352660 352894
rect 347058 352294 347154 352350
rect 347210 352294 347278 352350
rect 347334 352294 347402 352350
rect 347458 352294 347526 352350
rect 347582 352294 347678 352350
rect 347058 352226 347678 352294
rect 347058 352170 347154 352226
rect 347210 352170 347278 352226
rect 347334 352170 347402 352226
rect 347458 352170 347526 352226
rect 347582 352170 347678 352226
rect 347058 352102 347678 352170
rect 347058 352046 347154 352102
rect 347210 352046 347278 352102
rect 347334 352046 347402 352102
rect 347458 352046 347526 352102
rect 347582 352046 347678 352102
rect 347058 351978 347678 352046
rect 347058 351922 347154 351978
rect 347210 351922 347278 351978
rect 347334 351922 347402 351978
rect 347458 351922 347526 351978
rect 347582 351922 347678 351978
rect 345212 339668 345268 339678
rect 344428 332038 344484 332048
rect 344428 329476 344484 331982
rect 344428 329410 344484 329420
rect 343338 328294 343434 328350
rect 343490 328294 343558 328350
rect 343614 328294 343682 328350
rect 343738 328294 343806 328350
rect 343862 328294 343958 328350
rect 343338 328226 343958 328294
rect 343338 328170 343434 328226
rect 343490 328170 343558 328226
rect 343614 328170 343682 328226
rect 343738 328170 343806 328226
rect 343862 328170 343958 328226
rect 343338 328102 343958 328170
rect 343338 328046 343434 328102
rect 343490 328046 343558 328102
rect 343614 328046 343682 328102
rect 343738 328046 343806 328102
rect 343862 328046 343958 328102
rect 343338 327978 343958 328046
rect 343338 327922 343434 327978
rect 343490 327922 343558 327978
rect 343614 327922 343682 327978
rect 343738 327922 343806 327978
rect 343862 327922 343958 327978
rect 343338 310350 343958 327922
rect 343338 310294 343434 310350
rect 343490 310294 343558 310350
rect 343614 310294 343682 310350
rect 343738 310294 343806 310350
rect 343862 310294 343958 310350
rect 343338 310226 343958 310294
rect 343338 310170 343434 310226
rect 343490 310170 343558 310226
rect 343614 310170 343682 310226
rect 343738 310170 343806 310226
rect 343862 310170 343958 310226
rect 343338 310102 343958 310170
rect 343338 310046 343434 310102
rect 343490 310046 343558 310102
rect 343614 310046 343682 310102
rect 343738 310046 343806 310102
rect 343862 310046 343958 310102
rect 343338 309978 343958 310046
rect 343338 309922 343434 309978
rect 343490 309922 343558 309978
rect 343614 309922 343682 309978
rect 343738 309922 343806 309978
rect 343862 309922 343958 309978
rect 338492 299730 338548 299740
rect 343338 292350 343958 309922
rect 345212 305396 345268 339612
rect 345212 305330 345268 305340
rect 347058 334350 347678 351922
rect 352604 351316 352660 352828
rect 371808 352350 372128 352384
rect 371808 352294 371878 352350
rect 371934 352294 372002 352350
rect 372058 352294 372128 352350
rect 371808 352226 372128 352294
rect 371808 352170 371878 352226
rect 371934 352170 372002 352226
rect 372058 352170 372128 352226
rect 371808 352102 372128 352170
rect 371808 352046 371878 352102
rect 371934 352046 372002 352102
rect 372058 352046 372128 352102
rect 371808 351978 372128 352046
rect 371808 351922 371878 351978
rect 371934 351922 372002 351978
rect 372058 351922 372128 351978
rect 371808 351888 372128 351922
rect 352604 351250 352660 351260
rect 347058 334294 347154 334350
rect 347210 334294 347278 334350
rect 347334 334294 347402 334350
rect 347458 334294 347526 334350
rect 347582 334294 347678 334350
rect 347058 334226 347678 334294
rect 347058 334170 347154 334226
rect 347210 334170 347278 334226
rect 347334 334170 347402 334226
rect 347458 334170 347526 334226
rect 347582 334170 347678 334226
rect 347058 334102 347678 334170
rect 347058 334046 347154 334102
rect 347210 334046 347278 334102
rect 347334 334046 347402 334102
rect 347458 334046 347526 334102
rect 347582 334046 347678 334102
rect 347058 333978 347678 334046
rect 347058 333922 347154 333978
rect 347210 333922 347278 333978
rect 347334 333922 347402 333978
rect 347458 333922 347526 333978
rect 347582 333922 347678 333978
rect 347058 316350 347678 333922
rect 350252 348778 350308 348788
rect 350252 326676 350308 348722
rect 356448 346350 356768 346384
rect 356448 346294 356518 346350
rect 356574 346294 356642 346350
rect 356698 346294 356768 346350
rect 356448 346226 356768 346294
rect 356448 346170 356518 346226
rect 356574 346170 356642 346226
rect 356698 346170 356768 346226
rect 356448 346102 356768 346170
rect 356448 346046 356518 346102
rect 356574 346046 356642 346102
rect 356698 346046 356768 346102
rect 356448 345978 356768 346046
rect 356448 345922 356518 345978
rect 356574 345922 356642 345978
rect 356698 345922 356768 345978
rect 356448 345888 356768 345922
rect 374058 346350 374678 363922
rect 374058 346294 374154 346350
rect 374210 346294 374278 346350
rect 374334 346294 374402 346350
rect 374458 346294 374526 346350
rect 374582 346294 374678 346350
rect 374058 346226 374678 346294
rect 374058 346170 374154 346226
rect 374210 346170 374278 346226
rect 374334 346170 374402 346226
rect 374458 346170 374526 346226
rect 374582 346170 374678 346226
rect 374058 346102 374678 346170
rect 374058 346046 374154 346102
rect 374210 346046 374278 346102
rect 374334 346046 374402 346102
rect 374458 346046 374526 346102
rect 374582 346046 374678 346102
rect 374058 345978 374678 346046
rect 374058 345922 374154 345978
rect 374210 345922 374278 345978
rect 374334 345922 374402 345978
rect 374458 345922 374526 345978
rect 374582 345922 374678 345978
rect 352604 341236 352660 341246
rect 352716 341218 352772 341228
rect 352660 341180 352716 341218
rect 352604 341162 352716 341180
rect 352716 341152 352772 341162
rect 351148 339598 351204 339608
rect 351148 335636 351204 339542
rect 351148 335570 351204 335580
rect 371808 334350 372128 334384
rect 371808 334294 371878 334350
rect 371934 334294 372002 334350
rect 372058 334294 372128 334350
rect 371808 334226 372128 334294
rect 371808 334170 371878 334226
rect 371934 334170 372002 334226
rect 372058 334170 372128 334226
rect 371808 334102 372128 334170
rect 371808 334046 371878 334102
rect 371934 334046 372002 334102
rect 372058 334046 372128 334102
rect 371808 333978 372128 334046
rect 371808 333922 371878 333978
rect 371934 333922 372002 333978
rect 372058 333922 372128 333978
rect 371808 333888 372128 333922
rect 356448 328350 356768 328384
rect 356448 328294 356518 328350
rect 356574 328294 356642 328350
rect 356698 328294 356768 328350
rect 356448 328226 356768 328294
rect 356448 328170 356518 328226
rect 356574 328170 356642 328226
rect 356698 328170 356768 328226
rect 356448 328102 356768 328170
rect 356448 328046 356518 328102
rect 356574 328046 356642 328102
rect 356698 328046 356768 328102
rect 356448 327978 356768 328046
rect 356448 327922 356518 327978
rect 356574 327922 356642 327978
rect 356698 327922 356768 327978
rect 356448 327888 356768 327922
rect 374058 328350 374678 345922
rect 374058 328294 374154 328350
rect 374210 328294 374278 328350
rect 374334 328294 374402 328350
rect 374458 328294 374526 328350
rect 374582 328294 374678 328350
rect 374058 328226 374678 328294
rect 374058 328170 374154 328226
rect 374210 328170 374278 328226
rect 374334 328170 374402 328226
rect 374458 328170 374526 328226
rect 374582 328170 374678 328226
rect 374058 328102 374678 328170
rect 374058 328046 374154 328102
rect 374210 328046 374278 328102
rect 374334 328046 374402 328102
rect 374458 328046 374526 328102
rect 374582 328046 374678 328102
rect 374058 327978 374678 328046
rect 374058 327922 374154 327978
rect 374210 327922 374278 327978
rect 374334 327922 374402 327978
rect 374458 327922 374526 327978
rect 374582 327922 374678 327978
rect 350252 326610 350308 326620
rect 347058 316294 347154 316350
rect 347210 316294 347278 316350
rect 347334 316294 347402 316350
rect 347458 316294 347526 316350
rect 347582 316294 347678 316350
rect 347058 316226 347678 316294
rect 347058 316170 347154 316226
rect 347210 316170 347278 316226
rect 347334 316170 347402 316226
rect 347458 316170 347526 316226
rect 347582 316170 347678 316226
rect 347058 316102 347678 316170
rect 347058 316046 347154 316102
rect 347210 316046 347278 316102
rect 347334 316046 347402 316102
rect 347458 316046 347526 316102
rect 347582 316046 347678 316102
rect 347058 315978 347678 316046
rect 347058 315922 347154 315978
rect 347210 315922 347278 315978
rect 347334 315922 347402 315978
rect 347458 315922 347526 315978
rect 347582 315922 347678 315978
rect 343338 292294 343434 292350
rect 343490 292294 343558 292350
rect 343614 292294 343682 292350
rect 343738 292294 343806 292350
rect 343862 292294 343958 292350
rect 343338 292226 343958 292294
rect 343338 292170 343434 292226
rect 343490 292170 343558 292226
rect 343614 292170 343682 292226
rect 343738 292170 343806 292226
rect 343862 292170 343958 292226
rect 343338 292102 343958 292170
rect 343338 292046 343434 292102
rect 343490 292046 343558 292102
rect 343614 292046 343682 292102
rect 343738 292046 343806 292102
rect 343862 292046 343958 292102
rect 343338 291978 343958 292046
rect 343338 291922 343434 291978
rect 343490 291922 343558 291978
rect 343614 291922 343682 291978
rect 343738 291922 343806 291978
rect 343862 291922 343958 291978
rect 335916 290836 335972 290846
rect 335916 289828 335972 290780
rect 335916 289762 335972 289772
rect 334460 288148 334516 288158
rect 334460 287924 334516 288092
rect 334460 287858 334516 287868
rect 342636 284116 342692 284126
rect 342636 283220 342692 284060
rect 342636 283154 342692 283164
rect 334460 281652 334516 281662
rect 334460 279636 334516 281596
rect 334460 279570 334516 279580
rect 334460 278516 334516 278526
rect 334348 278038 334404 278048
rect 334348 275716 334404 277982
rect 334460 277318 334516 278460
rect 334460 277252 334516 277262
rect 334348 275650 334404 275660
rect 334460 276836 334516 276846
rect 334460 275698 334516 276780
rect 334460 275632 334516 275642
rect 336924 275156 336980 275166
rect 334572 274596 334628 274606
rect 334460 274036 334516 274046
rect 334348 273476 334404 273486
rect 334348 272278 334404 273420
rect 334460 272998 334516 273980
rect 334460 272932 334516 272942
rect 334348 272212 334404 272222
rect 334460 272356 334516 272366
rect 334460 271558 334516 272300
rect 334460 271492 334516 271502
rect 334460 270116 334516 270126
rect 334460 268858 334516 270060
rect 334572 269758 334628 274540
rect 334572 269692 334628 269702
rect 334460 268792 334516 268802
rect 335692 268996 335748 269006
rect 334348 268436 334404 268446
rect 334348 267418 334404 268380
rect 334348 267352 334404 267362
rect 334460 267958 334516 267968
rect 334460 267316 334516 267902
rect 334460 267250 334516 267260
rect 334460 266518 334516 266528
rect 334460 266196 334516 266462
rect 334460 266130 334516 266140
rect 334572 266338 334628 266348
rect 334460 265438 334516 265448
rect 334460 264516 334516 265382
rect 334460 264450 334516 264460
rect 334460 263956 334516 263966
rect 334460 263818 334516 263900
rect 334460 263752 334516 263762
rect 334460 263638 334516 263648
rect 334460 262836 334516 263582
rect 334460 262770 334516 262780
rect 334460 261716 334516 261726
rect 334460 260758 334516 261660
rect 334460 260692 334516 260702
rect 334460 260596 334516 260616
rect 334460 260512 334516 260522
rect 334460 260398 334516 260408
rect 334460 260036 334516 260342
rect 334460 259970 334516 259980
rect 334460 258958 334516 258968
rect 334460 258850 334516 258860
rect 334460 258598 334516 258608
rect 334348 258542 334460 258598
rect 334348 257796 334404 258542
rect 334460 258532 334516 258542
rect 334460 258356 334516 258366
rect 334460 258238 334516 258300
rect 334460 258172 334516 258182
rect 334348 257730 334404 257740
rect 334572 255556 334628 266282
rect 335692 266308 335748 268940
rect 336924 267058 336980 275100
rect 343338 274350 343958 291922
rect 343338 274294 343434 274350
rect 343490 274294 343558 274350
rect 343614 274294 343682 274350
rect 343738 274294 343806 274350
rect 343862 274294 343958 274350
rect 343338 274226 343958 274294
rect 343338 274170 343434 274226
rect 343490 274170 343558 274226
rect 343614 274170 343682 274226
rect 343738 274170 343806 274226
rect 343862 274170 343958 274226
rect 343338 274102 343958 274170
rect 343338 274046 343434 274102
rect 343490 274046 343558 274102
rect 343614 274046 343682 274102
rect 343738 274046 343806 274102
rect 343862 274046 343958 274102
rect 343338 273978 343958 274046
rect 343338 273922 343434 273978
rect 343490 273922 343558 273978
rect 343614 273922 343682 273978
rect 343738 273922 343806 273978
rect 343862 273922 343958 273978
rect 336924 266992 336980 267002
rect 338492 267764 338548 267774
rect 335692 266242 335748 266252
rect 334572 255490 334628 255500
rect 336812 265748 336868 265758
rect 334684 255358 334740 255368
rect 334460 255178 334516 255188
rect 334348 254998 334404 255008
rect 334348 253876 334404 254942
rect 334460 254996 334516 255122
rect 334460 254930 334516 254940
rect 334684 254436 334740 255302
rect 334684 254370 334740 254380
rect 334348 253810 334404 253820
rect 334460 253558 334516 253568
rect 334460 252756 334516 253502
rect 334460 252690 334516 252700
rect 334460 251938 334516 251948
rect 334348 251758 334404 251768
rect 334348 250516 334404 251702
rect 334460 251636 334516 251882
rect 334460 251570 334516 251580
rect 334348 250450 334404 250460
rect 334460 250138 334516 250148
rect 334460 248836 334516 250082
rect 334460 248770 334516 248780
rect 334460 248518 334516 248528
rect 334460 248276 334516 248462
rect 334460 248210 334516 248220
rect 336028 246260 336084 246270
rect 336028 243796 336084 246204
rect 336812 244356 336868 265692
rect 338492 247156 338548 267708
rect 338492 247090 338548 247100
rect 343338 256350 343958 273922
rect 347058 298350 347678 315922
rect 351932 320516 351988 320526
rect 351932 314038 351988 320460
rect 351932 313972 351988 313982
rect 347058 298294 347154 298350
rect 347210 298294 347278 298350
rect 347334 298294 347402 298350
rect 347458 298294 347526 298350
rect 347582 298294 347678 298350
rect 347058 298226 347678 298294
rect 347058 298170 347154 298226
rect 347210 298170 347278 298226
rect 347334 298170 347402 298226
rect 347458 298170 347526 298226
rect 347582 298170 347678 298226
rect 347058 298102 347678 298170
rect 347058 298046 347154 298102
rect 347210 298046 347278 298102
rect 347334 298046 347402 298102
rect 347458 298046 347526 298102
rect 347582 298046 347678 298102
rect 347058 297978 347678 298046
rect 347058 297922 347154 297978
rect 347210 297922 347278 297978
rect 347334 297922 347402 297978
rect 347458 297922 347526 297978
rect 347582 297922 347678 297978
rect 347058 280350 347678 297922
rect 374058 310350 374678 327922
rect 374058 310294 374154 310350
rect 374210 310294 374278 310350
rect 374334 310294 374402 310350
rect 374458 310294 374526 310350
rect 374582 310294 374678 310350
rect 374058 310226 374678 310294
rect 374058 310170 374154 310226
rect 374210 310170 374278 310226
rect 374334 310170 374402 310226
rect 374458 310170 374526 310226
rect 374582 310170 374678 310226
rect 374058 310102 374678 310170
rect 374058 310046 374154 310102
rect 374210 310046 374278 310102
rect 374334 310046 374402 310102
rect 374458 310046 374526 310102
rect 374582 310046 374678 310102
rect 374058 309978 374678 310046
rect 374058 309922 374154 309978
rect 374210 309922 374278 309978
rect 374334 309922 374402 309978
rect 374458 309922 374526 309978
rect 374582 309922 374678 309978
rect 374058 292350 374678 309922
rect 374058 292294 374154 292350
rect 374210 292294 374278 292350
rect 374334 292294 374402 292350
rect 374458 292294 374526 292350
rect 374582 292294 374678 292350
rect 374058 292226 374678 292294
rect 374058 292170 374154 292226
rect 374210 292170 374278 292226
rect 374334 292170 374402 292226
rect 374458 292170 374526 292226
rect 374582 292170 374678 292226
rect 374058 292102 374678 292170
rect 374058 292046 374154 292102
rect 374210 292046 374278 292102
rect 374334 292046 374402 292102
rect 374458 292046 374526 292102
rect 374582 292046 374678 292102
rect 374058 291978 374678 292046
rect 374058 291922 374154 291978
rect 374210 291922 374278 291978
rect 374334 291922 374402 291978
rect 374458 291922 374526 291978
rect 374582 291922 374678 291978
rect 352716 286916 352772 286926
rect 352716 283108 352772 286860
rect 352716 283042 352772 283052
rect 347058 280294 347154 280350
rect 347210 280294 347278 280350
rect 347334 280294 347402 280350
rect 347458 280294 347526 280350
rect 347582 280294 347678 280350
rect 347058 280226 347678 280294
rect 347058 280170 347154 280226
rect 347210 280170 347278 280226
rect 347334 280170 347402 280226
rect 347458 280170 347526 280226
rect 347582 280170 347678 280226
rect 347058 280102 347678 280170
rect 347058 280046 347154 280102
rect 347210 280046 347278 280102
rect 347334 280046 347402 280102
rect 347458 280046 347526 280102
rect 347582 280046 347678 280102
rect 347058 279978 347678 280046
rect 347058 279922 347154 279978
rect 347210 279922 347278 279978
rect 347334 279922 347402 279978
rect 347458 279922 347526 279978
rect 347582 279922 347678 279978
rect 343338 256294 343434 256350
rect 343490 256294 343558 256350
rect 343614 256294 343682 256350
rect 343738 256294 343806 256350
rect 343862 256294 343958 256350
rect 343338 256226 343958 256294
rect 343338 256170 343434 256226
rect 343490 256170 343558 256226
rect 343614 256170 343682 256226
rect 343738 256170 343806 256226
rect 343862 256170 343958 256226
rect 343338 256102 343958 256170
rect 343338 256046 343434 256102
rect 343490 256046 343558 256102
rect 343614 256046 343682 256102
rect 343738 256046 343806 256102
rect 343862 256046 343958 256102
rect 343338 255978 343958 256046
rect 343338 255922 343434 255978
rect 343490 255922 343558 255978
rect 343614 255922 343682 255978
rect 343738 255922 343806 255978
rect 343862 255922 343958 255978
rect 336812 244290 336868 244300
rect 336028 243730 336084 243740
rect 335916 239876 335972 239886
rect 335692 238756 335748 238766
rect 335132 237076 335188 237086
rect 335132 224308 335188 237020
rect 335132 224242 335188 224252
rect 335692 219268 335748 238700
rect 335916 231028 335972 239820
rect 335916 230962 335972 230972
rect 343338 238350 343958 255922
rect 345212 267092 345268 267102
rect 345212 244916 345268 267036
rect 347058 262350 347678 279922
rect 371808 280350 372128 280384
rect 371808 280294 371878 280350
rect 371934 280294 372002 280350
rect 372058 280294 372128 280350
rect 371808 280226 372128 280294
rect 371808 280170 371878 280226
rect 371934 280170 372002 280226
rect 372058 280170 372128 280226
rect 371808 280102 372128 280170
rect 371808 280046 371878 280102
rect 371934 280046 372002 280102
rect 372058 280046 372128 280102
rect 371808 279978 372128 280046
rect 371808 279922 371878 279978
rect 371934 279922 372002 279978
rect 372058 279922 372128 279978
rect 371808 279888 372128 279922
rect 356448 274350 356768 274384
rect 356448 274294 356518 274350
rect 356574 274294 356642 274350
rect 356698 274294 356768 274350
rect 356448 274226 356768 274294
rect 356448 274170 356518 274226
rect 356574 274170 356642 274226
rect 356698 274170 356768 274226
rect 356448 274102 356768 274170
rect 356448 274046 356518 274102
rect 356574 274046 356642 274102
rect 356698 274046 356768 274102
rect 356448 273978 356768 274046
rect 356448 273922 356518 273978
rect 356574 273922 356642 273978
rect 356698 273922 356768 273978
rect 356448 273888 356768 273922
rect 374058 274350 374678 291922
rect 374058 274294 374154 274350
rect 374210 274294 374278 274350
rect 374334 274294 374402 274350
rect 374458 274294 374526 274350
rect 374582 274294 374678 274350
rect 374058 274226 374678 274294
rect 374058 274170 374154 274226
rect 374210 274170 374278 274226
rect 374334 274170 374402 274226
rect 374458 274170 374526 274226
rect 374582 274170 374678 274226
rect 374058 274102 374678 274170
rect 374058 274046 374154 274102
rect 374210 274046 374278 274102
rect 374334 274046 374402 274102
rect 374458 274046 374526 274102
rect 374582 274046 374678 274102
rect 374058 273978 374678 274046
rect 374058 273922 374154 273978
rect 374210 273922 374278 273978
rect 374334 273922 374402 273978
rect 374458 273922 374526 273978
rect 374582 273922 374678 273978
rect 351036 272916 351092 272926
rect 351036 271738 351092 272860
rect 351036 271672 351092 271682
rect 352716 269578 352772 269588
rect 352716 268436 352772 269522
rect 352716 268370 352772 268380
rect 351932 267238 351988 267248
rect 347788 266308 347844 266318
rect 347788 265258 347844 266252
rect 347788 265192 347844 265202
rect 347058 262294 347154 262350
rect 347210 262294 347278 262350
rect 347334 262294 347402 262350
rect 347458 262294 347526 262350
rect 347582 262294 347678 262350
rect 347058 262226 347678 262294
rect 347058 262170 347154 262226
rect 347210 262170 347278 262226
rect 347334 262170 347402 262226
rect 347458 262170 347526 262226
rect 347582 262170 347678 262226
rect 347058 262102 347678 262170
rect 347058 262046 347154 262102
rect 347210 262046 347278 262102
rect 347334 262046 347402 262102
rect 347458 262046 347526 262102
rect 347582 262046 347678 262102
rect 347058 261978 347678 262046
rect 347058 261922 347154 261978
rect 347210 261922 347278 261978
rect 347334 261922 347402 261978
rect 347458 261922 347526 261978
rect 347582 261922 347678 261978
rect 346892 259700 346948 259710
rect 346892 246596 346948 259644
rect 346892 246530 346948 246540
rect 345212 244850 345268 244860
rect 345996 244468 346052 244478
rect 345996 240996 346052 244412
rect 345996 240930 346052 240940
rect 347058 244350 347678 261922
rect 348572 264404 348628 264414
rect 348572 246260 348628 264348
rect 348572 246194 348628 246204
rect 348796 261044 348852 261054
rect 348796 246036 348852 260988
rect 351036 258778 351092 258788
rect 351036 256116 351092 258722
rect 351932 256676 351988 267182
rect 371808 262350 372128 262384
rect 371808 262294 371878 262350
rect 371934 262294 372002 262350
rect 372058 262294 372128 262350
rect 371808 262226 372128 262294
rect 371808 262170 371878 262226
rect 371934 262170 372002 262226
rect 372058 262170 372128 262226
rect 371808 262102 372128 262170
rect 371808 262046 371878 262102
rect 371934 262046 372002 262102
rect 372058 262046 372128 262102
rect 371808 261978 372128 262046
rect 371808 261922 371878 261978
rect 371934 261922 372002 261978
rect 372058 261922 372128 261978
rect 371808 261888 372128 261922
rect 351932 256610 351988 256620
rect 351036 256050 351092 256060
rect 356448 256350 356768 256384
rect 356448 256294 356518 256350
rect 356574 256294 356642 256350
rect 356698 256294 356768 256350
rect 356448 256226 356768 256294
rect 356448 256170 356518 256226
rect 356574 256170 356642 256226
rect 356698 256170 356768 256226
rect 356448 256102 356768 256170
rect 356448 256046 356518 256102
rect 356574 256046 356642 256102
rect 356698 256046 356768 256102
rect 356448 255978 356768 256046
rect 356448 255922 356518 255978
rect 356574 255922 356642 255978
rect 356698 255922 356768 255978
rect 356448 255888 356768 255922
rect 374058 256350 374678 273922
rect 374058 256294 374154 256350
rect 374210 256294 374278 256350
rect 374334 256294 374402 256350
rect 374458 256294 374526 256350
rect 374582 256294 374678 256350
rect 374058 256226 374678 256294
rect 374058 256170 374154 256226
rect 374210 256170 374278 256226
rect 374334 256170 374402 256226
rect 374458 256170 374526 256226
rect 374582 256170 374678 256226
rect 374058 256102 374678 256170
rect 374058 256046 374154 256102
rect 374210 256046 374278 256102
rect 374334 256046 374402 256102
rect 374458 256046 374526 256102
rect 374582 256046 374678 256102
rect 374058 255978 374678 256046
rect 374058 255922 374154 255978
rect 374210 255922 374278 255978
rect 374334 255922 374402 255978
rect 374458 255922 374526 255978
rect 374582 255922 374678 255978
rect 351036 251076 351092 251086
rect 351036 250318 351092 251020
rect 351036 250252 351092 250262
rect 348796 245970 348852 245980
rect 351036 247716 351092 247726
rect 351036 245812 351092 247660
rect 351036 245746 351092 245756
rect 347058 244294 347154 244350
rect 347210 244294 347278 244350
rect 347334 244294 347402 244350
rect 347458 244294 347526 244350
rect 347582 244294 347678 244350
rect 347058 244226 347678 244294
rect 347058 244170 347154 244226
rect 347210 244170 347278 244226
rect 347334 244170 347402 244226
rect 347458 244170 347526 244226
rect 347582 244170 347678 244226
rect 347058 244102 347678 244170
rect 347058 244046 347154 244102
rect 347210 244046 347278 244102
rect 347334 244046 347402 244102
rect 347458 244046 347526 244102
rect 347582 244046 347678 244102
rect 347058 243978 347678 244046
rect 347058 243922 347154 243978
rect 347210 243922 347278 243978
rect 347334 243922 347402 243978
rect 347458 243922 347526 243978
rect 347582 243922 347678 243978
rect 343338 238294 343434 238350
rect 343490 238294 343558 238350
rect 343614 238294 343682 238350
rect 343738 238294 343806 238350
rect 343862 238294 343958 238350
rect 343338 238226 343958 238294
rect 343338 238170 343434 238226
rect 343490 238170 343558 238226
rect 343614 238170 343682 238226
rect 343738 238170 343806 238226
rect 343862 238170 343958 238226
rect 343338 238102 343958 238170
rect 343338 238046 343434 238102
rect 343490 238046 343558 238102
rect 343614 238046 343682 238102
rect 343738 238046 343806 238102
rect 343862 238046 343958 238102
rect 343338 237978 343958 238046
rect 343338 237922 343434 237978
rect 343490 237922 343558 237978
rect 343614 237922 343682 237978
rect 343738 237922 343806 237978
rect 343862 237922 343958 237978
rect 338492 225316 338548 225326
rect 335692 219202 335748 219212
rect 335916 220836 335972 220846
rect 335916 217588 335972 220780
rect 335916 217522 335972 217532
rect 336028 216356 336084 216366
rect 336028 214340 336084 216300
rect 336028 214274 336084 214284
rect 337036 215236 337092 215246
rect 334460 212884 334516 212894
rect 334460 212660 334516 212828
rect 334460 212594 334516 212604
rect 334460 206276 334516 206286
rect 334460 205138 334516 206220
rect 334460 205072 334516 205082
rect 334460 204596 334516 204606
rect 334460 203338 334516 204540
rect 334460 203272 334516 203282
rect 334460 202356 334516 202366
rect 334460 200818 334516 202300
rect 334460 200752 334516 200762
rect 334460 200676 334516 200686
rect 334460 200098 334516 200620
rect 334460 200032 334516 200042
rect 334460 198996 334516 199006
rect 334460 198298 334516 198940
rect 334460 198232 334516 198242
rect 334348 197876 334404 197886
rect 334348 196678 334404 197820
rect 334460 197316 334516 197326
rect 334460 196858 334516 197260
rect 334460 196792 334516 196802
rect 334460 196678 334516 196688
rect 334348 196622 334460 196678
rect 334460 196612 334516 196622
rect 337036 196532 337092 215180
rect 338492 214228 338548 225260
rect 343338 220350 343958 237922
rect 343338 220294 343434 220350
rect 343490 220294 343558 220350
rect 343614 220294 343682 220350
rect 343738 220294 343806 220350
rect 343862 220294 343958 220350
rect 343338 220226 343958 220294
rect 343338 220170 343434 220226
rect 343490 220170 343558 220226
rect 343614 220170 343682 220226
rect 343738 220170 343806 220226
rect 343862 220170 343958 220226
rect 343338 220102 343958 220170
rect 343338 220046 343434 220102
rect 343490 220046 343558 220102
rect 343614 220046 343682 220102
rect 343738 220046 343806 220102
rect 343862 220046 343958 220102
rect 343338 219978 343958 220046
rect 343338 219922 343434 219978
rect 343490 219922 343558 219978
rect 343614 219922 343682 219978
rect 343738 219922 343806 219978
rect 343862 219922 343958 219978
rect 338492 214162 338548 214172
rect 339276 219156 339332 219166
rect 339276 213220 339332 219100
rect 340396 214676 340452 214686
rect 339276 213154 339332 213164
rect 340172 213556 340228 213566
rect 337036 196466 337092 196476
rect 338492 211876 338548 211886
rect 334460 196196 334516 196206
rect 334460 195058 334516 196140
rect 334460 194992 334516 195002
rect 334460 194878 334516 194888
rect 334348 194822 334460 194878
rect 334348 193956 334404 194822
rect 334460 194812 334516 194822
rect 334460 194516 334516 194526
rect 334460 193978 334516 194460
rect 334460 193912 334516 193922
rect 334348 193890 334404 193900
rect 334460 193396 334516 193406
rect 334460 193258 334516 193340
rect 334460 193192 334516 193202
rect 334348 192724 334404 192734
rect 334348 190596 334404 192668
rect 334460 192358 334516 192368
rect 334460 192276 334516 192302
rect 334460 192210 334516 192220
rect 338492 191156 338548 211820
rect 340172 194516 340228 213500
rect 340172 194450 340228 194460
rect 340284 210196 340340 210206
rect 340284 192500 340340 210140
rect 340396 195188 340452 214620
rect 340620 214116 340676 214126
rect 340620 195860 340676 214060
rect 343338 202350 343958 219922
rect 347058 226350 347678 243922
rect 347058 226294 347154 226350
rect 347210 226294 347278 226350
rect 347334 226294 347402 226350
rect 347458 226294 347526 226350
rect 347582 226294 347678 226350
rect 347058 226226 347678 226294
rect 347058 226170 347154 226226
rect 347210 226170 347278 226226
rect 347334 226170 347402 226226
rect 347458 226170 347526 226226
rect 347582 226170 347678 226226
rect 347058 226102 347678 226170
rect 347058 226046 347154 226102
rect 347210 226046 347278 226102
rect 347334 226046 347402 226102
rect 347458 226046 347526 226102
rect 347582 226046 347678 226102
rect 347058 225978 347678 226046
rect 347058 225922 347154 225978
rect 347210 225922 347278 225978
rect 347334 225922 347402 225978
rect 347458 225922 347526 225978
rect 347582 225922 347678 225978
rect 345996 210532 346052 210542
rect 345996 203476 346052 210476
rect 345996 203410 346052 203420
rect 347058 208350 347678 225922
rect 374058 238350 374678 255922
rect 374058 238294 374154 238350
rect 374210 238294 374278 238350
rect 374334 238294 374402 238350
rect 374458 238294 374526 238350
rect 374582 238294 374678 238350
rect 374058 238226 374678 238294
rect 374058 238170 374154 238226
rect 374210 238170 374278 238226
rect 374334 238170 374402 238226
rect 374458 238170 374526 238226
rect 374582 238170 374678 238226
rect 374058 238102 374678 238170
rect 374058 238046 374154 238102
rect 374210 238046 374278 238102
rect 374334 238046 374402 238102
rect 374458 238046 374526 238102
rect 374582 238046 374678 238102
rect 374058 237978 374678 238046
rect 374058 237922 374154 237978
rect 374210 237922 374278 237978
rect 374334 237922 374402 237978
rect 374458 237922 374526 237978
rect 374582 237922 374678 237978
rect 351932 221396 351988 221406
rect 351932 211204 351988 221340
rect 374058 220350 374678 237922
rect 374058 220294 374154 220350
rect 374210 220294 374278 220350
rect 374334 220294 374402 220350
rect 374458 220294 374526 220350
rect 374582 220294 374678 220350
rect 374058 220226 374678 220294
rect 374058 220170 374154 220226
rect 374210 220170 374278 220226
rect 374334 220170 374402 220226
rect 374458 220170 374526 220226
rect 374582 220170 374678 220226
rect 374058 220102 374678 220170
rect 374058 220046 374154 220102
rect 374210 220046 374278 220102
rect 374334 220046 374402 220102
rect 374458 220046 374526 220102
rect 374582 220046 374678 220102
rect 374058 219978 374678 220046
rect 374058 219922 374154 219978
rect 374210 219922 374278 219978
rect 374334 219922 374402 219978
rect 374458 219922 374526 219978
rect 374582 219922 374678 219978
rect 356188 218036 356244 218046
rect 356188 214452 356244 217980
rect 356188 214386 356244 214396
rect 370860 212884 370916 212894
rect 370860 212436 370916 212828
rect 370860 212370 370916 212380
rect 351932 211138 351988 211148
rect 351148 210644 351204 210654
rect 351036 210420 351092 210430
rect 351036 209076 351092 210364
rect 351036 209010 351092 209020
rect 347058 208294 347154 208350
rect 347210 208294 347278 208350
rect 347334 208294 347402 208350
rect 347458 208294 347526 208350
rect 347582 208294 347678 208350
rect 347058 208226 347678 208294
rect 347058 208170 347154 208226
rect 347210 208170 347278 208226
rect 347334 208170 347402 208226
rect 347458 208170 347526 208226
rect 347582 208170 347678 208226
rect 347058 208102 347678 208170
rect 347058 208046 347154 208102
rect 347210 208046 347278 208102
rect 347334 208046 347402 208102
rect 347458 208046 347526 208102
rect 347582 208046 347678 208102
rect 347058 207978 347678 208046
rect 347058 207922 347154 207978
rect 347210 207922 347278 207978
rect 347334 207922 347402 207978
rect 347458 207922 347526 207978
rect 347582 207922 347678 207978
rect 343338 202294 343434 202350
rect 343490 202294 343558 202350
rect 343614 202294 343682 202350
rect 343738 202294 343806 202350
rect 343862 202294 343958 202350
rect 343338 202226 343958 202294
rect 343338 202170 343434 202226
rect 343490 202170 343558 202226
rect 343614 202170 343682 202226
rect 343738 202170 343806 202226
rect 343862 202170 343958 202226
rect 343338 202102 343958 202170
rect 343338 202046 343434 202102
rect 343490 202046 343558 202102
rect 343614 202046 343682 202102
rect 343738 202046 343806 202102
rect 343862 202046 343958 202102
rect 343338 201978 343958 202046
rect 343338 201922 343434 201978
rect 343490 201922 343558 201978
rect 343614 201922 343682 201978
rect 343738 201922 343806 201978
rect 343862 201922 343958 201978
rect 340620 195794 340676 195804
rect 341852 201796 341908 201806
rect 340396 195122 340452 195132
rect 340284 192434 340340 192444
rect 338492 191090 338548 191100
rect 334348 190530 334404 190540
rect 336028 190036 336084 190046
rect 335132 188938 335188 188948
rect 335132 183316 335188 188882
rect 336028 186418 336084 189980
rect 341852 188038 341908 201740
rect 341852 187972 341908 187982
rect 336028 186352 336084 186362
rect 336140 187318 336196 187328
rect 336140 184436 336196 187262
rect 342636 186676 342692 186686
rect 342636 186238 342692 186620
rect 342636 186172 342692 186182
rect 336140 184370 336196 184380
rect 335132 183250 335188 183260
rect 343338 184350 343958 201922
rect 347058 190350 347678 207922
rect 351148 207956 351204 210588
rect 351148 207890 351204 207900
rect 371808 208350 372128 208384
rect 371808 208294 371878 208350
rect 371934 208294 372002 208350
rect 372058 208294 372128 208350
rect 371808 208226 372128 208294
rect 371808 208170 371878 208226
rect 371934 208170 372002 208226
rect 372058 208170 372128 208226
rect 371808 208102 372128 208170
rect 371808 208046 371878 208102
rect 371934 208046 372002 208102
rect 372058 208046 372128 208102
rect 371808 207978 372128 208046
rect 371808 207922 371878 207978
rect 371934 207922 372002 207978
rect 372058 207922 372128 207978
rect 371808 207888 372128 207922
rect 356448 202350 356768 202384
rect 356448 202294 356518 202350
rect 356574 202294 356642 202350
rect 356698 202294 356768 202350
rect 356448 202226 356768 202294
rect 356448 202170 356518 202226
rect 356574 202170 356642 202226
rect 356698 202170 356768 202226
rect 356448 202102 356768 202170
rect 356448 202046 356518 202102
rect 356574 202046 356642 202102
rect 356698 202046 356768 202102
rect 356448 201978 356768 202046
rect 356448 201922 356518 201978
rect 356574 201922 356642 201978
rect 356698 201922 356768 201978
rect 356448 201888 356768 201922
rect 374058 202350 374678 219922
rect 377778 388350 378398 405922
rect 394828 410116 394884 410126
rect 387168 400350 387488 400384
rect 387168 400294 387238 400350
rect 387294 400294 387362 400350
rect 387418 400294 387488 400350
rect 387168 400226 387488 400294
rect 387168 400170 387238 400226
rect 387294 400170 387362 400226
rect 387418 400170 387488 400226
rect 387168 400102 387488 400170
rect 387168 400046 387238 400102
rect 387294 400046 387362 400102
rect 387418 400046 387488 400102
rect 387168 399978 387488 400046
rect 387168 399922 387238 399978
rect 387294 399922 387362 399978
rect 387418 399922 387488 399978
rect 387168 399888 387488 399922
rect 377778 388294 377874 388350
rect 377930 388294 377998 388350
rect 378054 388294 378122 388350
rect 378178 388294 378246 388350
rect 378302 388294 378398 388350
rect 377778 388226 378398 388294
rect 377778 388170 377874 388226
rect 377930 388170 377998 388226
rect 378054 388170 378122 388226
rect 378178 388170 378246 388226
rect 378302 388170 378398 388226
rect 377778 388102 378398 388170
rect 377778 388046 377874 388102
rect 377930 388046 377998 388102
rect 378054 388046 378122 388102
rect 378178 388046 378246 388102
rect 378302 388046 378398 388102
rect 377778 387978 378398 388046
rect 377778 387922 377874 387978
rect 377930 387922 377998 387978
rect 378054 387922 378122 387978
rect 378178 387922 378246 387978
rect 378302 387922 378398 387978
rect 377778 370350 378398 387922
rect 377778 370294 377874 370350
rect 377930 370294 377998 370350
rect 378054 370294 378122 370350
rect 378178 370294 378246 370350
rect 378302 370294 378398 370350
rect 377778 370226 378398 370294
rect 377778 370170 377874 370226
rect 377930 370170 377998 370226
rect 378054 370170 378122 370226
rect 378178 370170 378246 370226
rect 378302 370170 378398 370226
rect 377778 370102 378398 370170
rect 377778 370046 377874 370102
rect 377930 370046 377998 370102
rect 378054 370046 378122 370102
rect 378178 370046 378246 370102
rect 378302 370046 378398 370102
rect 377778 369978 378398 370046
rect 377778 369922 377874 369978
rect 377930 369922 377998 369978
rect 378054 369922 378122 369978
rect 378178 369922 378246 369978
rect 378302 369922 378398 369978
rect 377778 352350 378398 369922
rect 392252 381332 392308 381342
rect 392252 361956 392308 381276
rect 393148 365428 393204 365438
rect 393148 364196 393204 365372
rect 393148 364130 393204 364140
rect 394828 362068 394884 410060
rect 394940 408100 394996 408110
rect 394940 368788 394996 408044
rect 395052 406084 395108 406094
rect 395052 378868 395108 406028
rect 395612 385588 395668 419916
rect 395612 385522 395668 385532
rect 396508 404740 396564 404750
rect 395052 378802 395108 378812
rect 394940 368722 394996 368732
rect 396508 365540 396564 404684
rect 396620 387716 396676 421484
rect 404778 418350 405398 435922
rect 404778 418294 404874 418350
rect 404930 418294 404998 418350
rect 405054 418294 405122 418350
rect 405178 418294 405246 418350
rect 405302 418294 405398 418350
rect 404778 418226 405398 418294
rect 404778 418170 404874 418226
rect 404930 418170 404998 418226
rect 405054 418170 405122 418226
rect 405178 418170 405246 418226
rect 405302 418170 405398 418226
rect 404778 418102 405398 418170
rect 404778 418046 404874 418102
rect 404930 418046 404998 418102
rect 405054 418046 405122 418102
rect 405178 418046 405246 418102
rect 405302 418046 405398 418102
rect 404778 417978 405398 418046
rect 404778 417922 404874 417978
rect 404930 417922 404998 417978
rect 405054 417922 405122 417978
rect 405178 417922 405246 417978
rect 405302 417922 405398 417978
rect 402332 410116 402388 410126
rect 401436 409978 401492 409988
rect 401436 408178 401492 409922
rect 401436 408112 401492 408122
rect 396620 387650 396676 387660
rect 396732 403396 396788 403406
rect 396732 381332 396788 403340
rect 401212 402724 401268 402734
rect 396732 381266 396788 381276
rect 398972 402388 399028 402398
rect 398972 366996 399028 402332
rect 401212 397918 401268 402668
rect 401212 397852 401268 397862
rect 401436 398998 401492 399008
rect 401324 397378 401380 397388
rect 401324 393058 401380 397322
rect 401436 396298 401492 398942
rect 401436 396232 401492 396242
rect 401324 392992 401380 393002
rect 400652 385588 400708 385598
rect 400652 374836 400708 385532
rect 400652 374770 400708 374780
rect 402332 367108 402388 410060
rect 402332 367042 402388 367052
rect 404778 400350 405398 417922
rect 408498 598172 409118 598268
rect 408498 598116 408594 598172
rect 408650 598116 408718 598172
rect 408774 598116 408842 598172
rect 408898 598116 408966 598172
rect 409022 598116 409118 598172
rect 408498 598048 409118 598116
rect 408498 597992 408594 598048
rect 408650 597992 408718 598048
rect 408774 597992 408842 598048
rect 408898 597992 408966 598048
rect 409022 597992 409118 598048
rect 408498 597924 409118 597992
rect 408498 597868 408594 597924
rect 408650 597868 408718 597924
rect 408774 597868 408842 597924
rect 408898 597868 408966 597924
rect 409022 597868 409118 597924
rect 408498 597800 409118 597868
rect 408498 597744 408594 597800
rect 408650 597744 408718 597800
rect 408774 597744 408842 597800
rect 408898 597744 408966 597800
rect 409022 597744 409118 597800
rect 408498 586350 409118 597744
rect 408498 586294 408594 586350
rect 408650 586294 408718 586350
rect 408774 586294 408842 586350
rect 408898 586294 408966 586350
rect 409022 586294 409118 586350
rect 408498 586226 409118 586294
rect 408498 586170 408594 586226
rect 408650 586170 408718 586226
rect 408774 586170 408842 586226
rect 408898 586170 408966 586226
rect 409022 586170 409118 586226
rect 408498 586102 409118 586170
rect 408498 586046 408594 586102
rect 408650 586046 408718 586102
rect 408774 586046 408842 586102
rect 408898 586046 408966 586102
rect 409022 586046 409118 586102
rect 408498 585978 409118 586046
rect 408498 585922 408594 585978
rect 408650 585922 408718 585978
rect 408774 585922 408842 585978
rect 408898 585922 408966 585978
rect 409022 585922 409118 585978
rect 408498 568350 409118 585922
rect 408498 568294 408594 568350
rect 408650 568294 408718 568350
rect 408774 568294 408842 568350
rect 408898 568294 408966 568350
rect 409022 568294 409118 568350
rect 408498 568226 409118 568294
rect 408498 568170 408594 568226
rect 408650 568170 408718 568226
rect 408774 568170 408842 568226
rect 408898 568170 408966 568226
rect 409022 568170 409118 568226
rect 408498 568102 409118 568170
rect 408498 568046 408594 568102
rect 408650 568046 408718 568102
rect 408774 568046 408842 568102
rect 408898 568046 408966 568102
rect 409022 568046 409118 568102
rect 408498 567978 409118 568046
rect 408498 567922 408594 567978
rect 408650 567922 408718 567978
rect 408774 567922 408842 567978
rect 408898 567922 408966 567978
rect 409022 567922 409118 567978
rect 408498 550350 409118 567922
rect 435498 597212 436118 598268
rect 435498 597156 435594 597212
rect 435650 597156 435718 597212
rect 435774 597156 435842 597212
rect 435898 597156 435966 597212
rect 436022 597156 436118 597212
rect 435498 597088 436118 597156
rect 435498 597032 435594 597088
rect 435650 597032 435718 597088
rect 435774 597032 435842 597088
rect 435898 597032 435966 597088
rect 436022 597032 436118 597088
rect 435498 596964 436118 597032
rect 435498 596908 435594 596964
rect 435650 596908 435718 596964
rect 435774 596908 435842 596964
rect 435898 596908 435966 596964
rect 436022 596908 436118 596964
rect 435498 596840 436118 596908
rect 435498 596784 435594 596840
rect 435650 596784 435718 596840
rect 435774 596784 435842 596840
rect 435898 596784 435966 596840
rect 436022 596784 436118 596840
rect 435498 580350 436118 596784
rect 435498 580294 435594 580350
rect 435650 580294 435718 580350
rect 435774 580294 435842 580350
rect 435898 580294 435966 580350
rect 436022 580294 436118 580350
rect 435498 580226 436118 580294
rect 435498 580170 435594 580226
rect 435650 580170 435718 580226
rect 435774 580170 435842 580226
rect 435898 580170 435966 580226
rect 436022 580170 436118 580226
rect 435498 580102 436118 580170
rect 435498 580046 435594 580102
rect 435650 580046 435718 580102
rect 435774 580046 435842 580102
rect 435898 580046 435966 580102
rect 436022 580046 436118 580102
rect 435498 579978 436118 580046
rect 435498 579922 435594 579978
rect 435650 579922 435718 579978
rect 435774 579922 435842 579978
rect 435898 579922 435966 579978
rect 436022 579922 436118 579978
rect 418448 562350 418768 562384
rect 418448 562294 418518 562350
rect 418574 562294 418642 562350
rect 418698 562294 418768 562350
rect 418448 562226 418768 562294
rect 418448 562170 418518 562226
rect 418574 562170 418642 562226
rect 418698 562170 418768 562226
rect 418448 562102 418768 562170
rect 418448 562046 418518 562102
rect 418574 562046 418642 562102
rect 418698 562046 418768 562102
rect 418448 561978 418768 562046
rect 418448 561922 418518 561978
rect 418574 561922 418642 561978
rect 418698 561922 418768 561978
rect 418448 561888 418768 561922
rect 435498 562350 436118 579922
rect 435498 562294 435594 562350
rect 435650 562294 435718 562350
rect 435774 562294 435842 562350
rect 435898 562294 435966 562350
rect 436022 562294 436118 562350
rect 435498 562226 436118 562294
rect 435498 562170 435594 562226
rect 435650 562170 435718 562226
rect 435774 562170 435842 562226
rect 435898 562170 435966 562226
rect 436022 562170 436118 562226
rect 435498 562102 436118 562170
rect 435498 562046 435594 562102
rect 435650 562046 435718 562102
rect 435774 562046 435842 562102
rect 435898 562046 435966 562102
rect 436022 562046 436118 562102
rect 435498 561978 436118 562046
rect 435498 561922 435594 561978
rect 435650 561922 435718 561978
rect 435774 561922 435842 561978
rect 435898 561922 435966 561978
rect 436022 561922 436118 561978
rect 414652 555238 414708 555248
rect 414652 555156 414708 555182
rect 414652 555090 414708 555100
rect 410956 553924 411012 553934
rect 408498 550294 408594 550350
rect 408650 550294 408718 550350
rect 408774 550294 408842 550350
rect 408898 550294 408966 550350
rect 409022 550294 409118 550350
rect 408498 550226 409118 550294
rect 408498 550170 408594 550226
rect 408650 550170 408718 550226
rect 408774 550170 408842 550226
rect 408898 550170 408966 550226
rect 409022 550170 409118 550226
rect 408498 550102 409118 550170
rect 408498 550046 408594 550102
rect 408650 550046 408718 550102
rect 408774 550046 408842 550102
rect 408898 550046 408966 550102
rect 409022 550046 409118 550102
rect 408498 549978 409118 550046
rect 408498 549922 408594 549978
rect 408650 549922 408718 549978
rect 408774 549922 408842 549978
rect 408898 549922 408966 549978
rect 409022 549922 409118 549978
rect 408498 532350 409118 549922
rect 408498 532294 408594 532350
rect 408650 532294 408718 532350
rect 408774 532294 408842 532350
rect 408898 532294 408966 532350
rect 409022 532294 409118 532350
rect 408498 532226 409118 532294
rect 408498 532170 408594 532226
rect 408650 532170 408718 532226
rect 408774 532170 408842 532226
rect 408898 532170 408966 532226
rect 409022 532170 409118 532226
rect 408498 532102 409118 532170
rect 408498 532046 408594 532102
rect 408650 532046 408718 532102
rect 408774 532046 408842 532102
rect 408898 532046 408966 532102
rect 409022 532046 409118 532102
rect 408498 531978 409118 532046
rect 408498 531922 408594 531978
rect 408650 531922 408718 531978
rect 408774 531922 408842 531978
rect 408898 531922 408966 531978
rect 409022 531922 409118 531978
rect 408498 514350 409118 531922
rect 408498 514294 408594 514350
rect 408650 514294 408718 514350
rect 408774 514294 408842 514350
rect 408898 514294 408966 514350
rect 409022 514294 409118 514350
rect 408498 514226 409118 514294
rect 408498 514170 408594 514226
rect 408650 514170 408718 514226
rect 408774 514170 408842 514226
rect 408898 514170 408966 514226
rect 409022 514170 409118 514226
rect 408498 514102 409118 514170
rect 408498 514046 408594 514102
rect 408650 514046 408718 514102
rect 408774 514046 408842 514102
rect 408898 514046 408966 514102
rect 409022 514046 409118 514102
rect 408498 513978 409118 514046
rect 408498 513922 408594 513978
rect 408650 513922 408718 513978
rect 408774 513922 408842 513978
rect 408898 513922 408966 513978
rect 409022 513922 409118 513978
rect 408498 496350 409118 513922
rect 410732 553252 410788 553262
rect 410732 505204 410788 553196
rect 410844 549892 410900 549902
rect 410844 508340 410900 549836
rect 410844 508274 410900 508284
rect 410956 506884 411012 553868
rect 435498 551870 436118 561922
rect 439218 598172 439838 598268
rect 439218 598116 439314 598172
rect 439370 598116 439438 598172
rect 439494 598116 439562 598172
rect 439618 598116 439686 598172
rect 439742 598116 439838 598172
rect 439218 598048 439838 598116
rect 439218 597992 439314 598048
rect 439370 597992 439438 598048
rect 439494 597992 439562 598048
rect 439618 597992 439686 598048
rect 439742 597992 439838 598048
rect 439218 597924 439838 597992
rect 439218 597868 439314 597924
rect 439370 597868 439438 597924
rect 439494 597868 439562 597924
rect 439618 597868 439686 597924
rect 439742 597868 439838 597924
rect 439218 597800 439838 597868
rect 439218 597744 439314 597800
rect 439370 597744 439438 597800
rect 439494 597744 439562 597800
rect 439618 597744 439686 597800
rect 439742 597744 439838 597800
rect 439218 586350 439838 597744
rect 439218 586294 439314 586350
rect 439370 586294 439438 586350
rect 439494 586294 439562 586350
rect 439618 586294 439686 586350
rect 439742 586294 439838 586350
rect 439218 586226 439838 586294
rect 439218 586170 439314 586226
rect 439370 586170 439438 586226
rect 439494 586170 439562 586226
rect 439618 586170 439686 586226
rect 439742 586170 439838 586226
rect 439218 586102 439838 586170
rect 439218 586046 439314 586102
rect 439370 586046 439438 586102
rect 439494 586046 439562 586102
rect 439618 586046 439686 586102
rect 439742 586046 439838 586102
rect 439218 585978 439838 586046
rect 439218 585922 439314 585978
rect 439370 585922 439438 585978
rect 439494 585922 439562 585978
rect 439618 585922 439686 585978
rect 439742 585922 439838 585978
rect 439218 568350 439838 585922
rect 439218 568294 439314 568350
rect 439370 568294 439438 568350
rect 439494 568294 439562 568350
rect 439618 568294 439686 568350
rect 439742 568294 439838 568350
rect 439218 568226 439838 568294
rect 439218 568170 439314 568226
rect 439370 568170 439438 568226
rect 439494 568170 439562 568226
rect 439618 568170 439686 568226
rect 439742 568170 439838 568226
rect 439218 568102 439838 568170
rect 439218 568046 439314 568102
rect 439370 568046 439438 568102
rect 439494 568046 439562 568102
rect 439618 568046 439686 568102
rect 439742 568046 439838 568102
rect 439218 567978 439838 568046
rect 439218 567922 439314 567978
rect 439370 567922 439438 567978
rect 439494 567922 439562 567978
rect 439618 567922 439686 567978
rect 439742 567922 439838 567978
rect 439218 551870 439838 567922
rect 466218 597212 466838 598268
rect 466218 597156 466314 597212
rect 466370 597156 466438 597212
rect 466494 597156 466562 597212
rect 466618 597156 466686 597212
rect 466742 597156 466838 597212
rect 466218 597088 466838 597156
rect 466218 597032 466314 597088
rect 466370 597032 466438 597088
rect 466494 597032 466562 597088
rect 466618 597032 466686 597088
rect 466742 597032 466838 597088
rect 466218 596964 466838 597032
rect 466218 596908 466314 596964
rect 466370 596908 466438 596964
rect 466494 596908 466562 596964
rect 466618 596908 466686 596964
rect 466742 596908 466838 596964
rect 466218 596840 466838 596908
rect 466218 596784 466314 596840
rect 466370 596784 466438 596840
rect 466494 596784 466562 596840
rect 466618 596784 466686 596840
rect 466742 596784 466838 596840
rect 466218 580350 466838 596784
rect 466218 580294 466314 580350
rect 466370 580294 466438 580350
rect 466494 580294 466562 580350
rect 466618 580294 466686 580350
rect 466742 580294 466838 580350
rect 466218 580226 466838 580294
rect 466218 580170 466314 580226
rect 466370 580170 466438 580226
rect 466494 580170 466562 580226
rect 466618 580170 466686 580226
rect 466742 580170 466838 580226
rect 466218 580102 466838 580170
rect 466218 580046 466314 580102
rect 466370 580046 466438 580102
rect 466494 580046 466562 580102
rect 466618 580046 466686 580102
rect 466742 580046 466838 580102
rect 466218 579978 466838 580046
rect 466218 579922 466314 579978
rect 466370 579922 466438 579978
rect 466494 579922 466562 579978
rect 466618 579922 466686 579978
rect 466742 579922 466838 579978
rect 449168 562350 449488 562384
rect 449168 562294 449238 562350
rect 449294 562294 449362 562350
rect 449418 562294 449488 562350
rect 449168 562226 449488 562294
rect 449168 562170 449238 562226
rect 449294 562170 449362 562226
rect 449418 562170 449488 562226
rect 449168 562102 449488 562170
rect 449168 562046 449238 562102
rect 449294 562046 449362 562102
rect 449418 562046 449488 562102
rect 449168 561978 449488 562046
rect 449168 561922 449238 561978
rect 449294 561922 449362 561978
rect 449418 561922 449488 561978
rect 449168 561888 449488 561922
rect 466218 562350 466838 579922
rect 466218 562294 466314 562350
rect 466370 562294 466438 562350
rect 466494 562294 466562 562350
rect 466618 562294 466686 562350
rect 466742 562294 466838 562350
rect 466218 562226 466838 562294
rect 466218 562170 466314 562226
rect 466370 562170 466438 562226
rect 466494 562170 466562 562226
rect 466618 562170 466686 562226
rect 466742 562170 466838 562226
rect 466218 562102 466838 562170
rect 466218 562046 466314 562102
rect 466370 562046 466438 562102
rect 466494 562046 466562 562102
rect 466618 562046 466686 562102
rect 466742 562046 466838 562102
rect 466218 561978 466838 562046
rect 466218 561922 466314 561978
rect 466370 561922 466438 561978
rect 466494 561922 466562 561978
rect 466618 561922 466686 561978
rect 466742 561922 466838 561978
rect 458780 553252 458836 553262
rect 458668 551908 458724 551918
rect 433808 550350 434128 550384
rect 433808 550294 433878 550350
rect 433934 550294 434002 550350
rect 434058 550294 434128 550350
rect 433808 550226 434128 550294
rect 433808 550170 433878 550226
rect 433934 550170 434002 550226
rect 434058 550170 434128 550226
rect 433808 550102 434128 550170
rect 433808 550046 433878 550102
rect 433934 550046 434002 550102
rect 434058 550046 434128 550102
rect 433808 549978 434128 550046
rect 433808 549922 433878 549978
rect 433934 549922 434002 549978
rect 434058 549922 434128 549978
rect 433808 549888 434128 549922
rect 456988 548548 457044 548558
rect 456092 547764 456148 547774
rect 411068 546532 411124 546542
rect 411068 520212 411124 546476
rect 418448 544350 418768 544384
rect 418448 544294 418518 544350
rect 418574 544294 418642 544350
rect 418698 544294 418768 544350
rect 418448 544226 418768 544294
rect 418448 544170 418518 544226
rect 418574 544170 418642 544226
rect 418698 544170 418768 544226
rect 418448 544102 418768 544170
rect 418448 544046 418518 544102
rect 418574 544046 418642 544102
rect 418698 544046 418768 544102
rect 418448 543978 418768 544046
rect 418448 543922 418518 543978
rect 418574 543922 418642 543978
rect 418698 543922 418768 543978
rect 418448 543888 418768 543922
rect 449168 544350 449488 544384
rect 449168 544294 449238 544350
rect 449294 544294 449362 544350
rect 449418 544294 449488 544350
rect 449168 544226 449488 544294
rect 449168 544170 449238 544226
rect 449294 544170 449362 544226
rect 449418 544170 449488 544226
rect 449168 544102 449488 544170
rect 449168 544046 449238 544102
rect 449294 544046 449362 544102
rect 449418 544046 449488 544102
rect 449168 543978 449488 544046
rect 449168 543922 449238 543978
rect 449294 543922 449362 543978
rect 449418 543922 449488 543978
rect 449168 543888 449488 543922
rect 455308 542500 455364 542510
rect 433808 532350 434128 532384
rect 433808 532294 433878 532350
rect 433934 532294 434002 532350
rect 434058 532294 434128 532350
rect 433808 532226 434128 532294
rect 433808 532170 433878 532226
rect 433934 532170 434002 532226
rect 434058 532170 434128 532226
rect 433808 532102 434128 532170
rect 433808 532046 433878 532102
rect 433934 532046 434002 532102
rect 434058 532046 434128 532102
rect 433808 531978 434128 532046
rect 433808 531922 433878 531978
rect 433934 531922 434002 531978
rect 434058 531922 434128 531978
rect 433808 531888 434128 531922
rect 411068 520146 411124 520156
rect 435498 526350 436118 540962
rect 435498 526294 435594 526350
rect 435650 526294 435718 526350
rect 435774 526294 435842 526350
rect 435898 526294 435966 526350
rect 436022 526294 436118 526350
rect 435498 526226 436118 526294
rect 435498 526170 435594 526226
rect 435650 526170 435718 526226
rect 435774 526170 435842 526226
rect 435898 526170 435966 526226
rect 436022 526170 436118 526226
rect 435498 526102 436118 526170
rect 435498 526046 435594 526102
rect 435650 526046 435718 526102
rect 435774 526046 435842 526102
rect 435898 526046 435966 526102
rect 436022 526046 436118 526102
rect 435498 525978 436118 526046
rect 435498 525922 435594 525978
rect 435650 525922 435718 525978
rect 435774 525922 435842 525978
rect 435898 525922 435966 525978
rect 436022 525922 436118 525978
rect 410956 506818 411012 506828
rect 435498 508350 436118 525922
rect 435498 508294 435594 508350
rect 435650 508294 435718 508350
rect 435774 508294 435842 508350
rect 435898 508294 435966 508350
rect 436022 508294 436118 508350
rect 435498 508226 436118 508294
rect 435498 508170 435594 508226
rect 435650 508170 435718 508226
rect 435774 508170 435842 508226
rect 435898 508170 435966 508226
rect 436022 508170 436118 508226
rect 435498 508102 436118 508170
rect 435498 508046 435594 508102
rect 435650 508046 435718 508102
rect 435774 508046 435842 508102
rect 435898 508046 435966 508102
rect 436022 508046 436118 508102
rect 435498 507978 436118 508046
rect 435498 507922 435594 507978
rect 435650 507922 435718 507978
rect 435774 507922 435842 507978
rect 435898 507922 435966 507978
rect 436022 507922 436118 507978
rect 410732 505138 410788 505148
rect 408498 496294 408594 496350
rect 408650 496294 408718 496350
rect 408774 496294 408842 496350
rect 408898 496294 408966 496350
rect 409022 496294 409118 496350
rect 408498 496226 409118 496294
rect 408498 496170 408594 496226
rect 408650 496170 408718 496226
rect 408774 496170 408842 496226
rect 408898 496170 408966 496226
rect 409022 496170 409118 496226
rect 408498 496102 409118 496170
rect 408498 496046 408594 496102
rect 408650 496046 408718 496102
rect 408774 496046 408842 496102
rect 408898 496046 408966 496102
rect 409022 496046 409118 496102
rect 408498 495978 409118 496046
rect 408498 495922 408594 495978
rect 408650 495922 408718 495978
rect 408774 495922 408842 495978
rect 408898 495922 408966 495978
rect 409022 495922 409118 495978
rect 408498 478350 409118 495922
rect 418448 490350 418768 490384
rect 418448 490294 418518 490350
rect 418574 490294 418642 490350
rect 418698 490294 418768 490350
rect 418448 490226 418768 490294
rect 418448 490170 418518 490226
rect 418574 490170 418642 490226
rect 418698 490170 418768 490226
rect 418448 490102 418768 490170
rect 418448 490046 418518 490102
rect 418574 490046 418642 490102
rect 418698 490046 418768 490102
rect 418448 489978 418768 490046
rect 418448 489922 418518 489978
rect 418574 489922 418642 489978
rect 418698 489922 418768 489978
rect 418448 489888 418768 489922
rect 435498 490350 436118 507922
rect 435498 490294 435594 490350
rect 435650 490294 435718 490350
rect 435774 490294 435842 490350
rect 435898 490294 435966 490350
rect 436022 490294 436118 490350
rect 435498 490226 436118 490294
rect 435498 490170 435594 490226
rect 435650 490170 435718 490226
rect 435774 490170 435842 490226
rect 435898 490170 435966 490226
rect 436022 490170 436118 490226
rect 435498 490102 436118 490170
rect 435498 490046 435594 490102
rect 435650 490046 435718 490102
rect 435774 490046 435842 490102
rect 435898 490046 435966 490102
rect 436022 490046 436118 490102
rect 435498 489978 436118 490046
rect 435498 489922 435594 489978
rect 435650 489922 435718 489978
rect 435774 489922 435842 489978
rect 435898 489922 435966 489978
rect 436022 489922 436118 489978
rect 414652 483958 414708 483968
rect 408498 478294 408594 478350
rect 408650 478294 408718 478350
rect 408774 478294 408842 478350
rect 408898 478294 408966 478350
rect 409022 478294 409118 478350
rect 408498 478226 409118 478294
rect 408498 478170 408594 478226
rect 408650 478170 408718 478226
rect 408774 478170 408842 478226
rect 408898 478170 408966 478226
rect 409022 478170 409118 478226
rect 408498 478102 409118 478170
rect 408498 478046 408594 478102
rect 408650 478046 408718 478102
rect 408774 478046 408842 478102
rect 408898 478046 408966 478102
rect 409022 478046 409118 478102
rect 408498 477978 409118 478046
rect 408498 477922 408594 477978
rect 408650 477922 408718 477978
rect 408774 477922 408842 477978
rect 408898 477922 408966 477978
rect 409022 477922 409118 477978
rect 408498 460350 409118 477922
rect 410844 482692 410900 482702
rect 408498 460294 408594 460350
rect 408650 460294 408718 460350
rect 408774 460294 408842 460350
rect 408898 460294 408966 460350
rect 409022 460294 409118 460350
rect 408498 460226 409118 460294
rect 408498 460170 408594 460226
rect 408650 460170 408718 460226
rect 408774 460170 408842 460226
rect 408898 460170 408966 460226
rect 409022 460170 409118 460226
rect 408498 460102 409118 460170
rect 408498 460046 408594 460102
rect 408650 460046 408718 460102
rect 408774 460046 408842 460102
rect 408898 460046 408966 460102
rect 409022 460046 409118 460102
rect 408498 459978 409118 460046
rect 408498 459922 408594 459978
rect 408650 459922 408718 459978
rect 408774 459922 408842 459978
rect 408898 459922 408966 459978
rect 409022 459922 409118 459978
rect 408498 442350 409118 459922
rect 410732 473284 410788 473294
rect 410732 446404 410788 473228
rect 410844 462868 410900 482636
rect 411180 482020 411236 482030
rect 410844 462802 410900 462812
rect 410956 481348 411012 481358
rect 410732 446338 410788 446348
rect 410956 446292 411012 481292
rect 411180 456372 411236 481964
rect 414652 481124 414708 483902
rect 414652 481058 414708 481068
rect 433808 478350 434128 478384
rect 433808 478294 433878 478350
rect 433934 478294 434002 478350
rect 434058 478294 434128 478350
rect 433808 478226 434128 478294
rect 433808 478170 433878 478226
rect 433934 478170 434002 478226
rect 434058 478170 434128 478226
rect 433808 478102 434128 478170
rect 433808 478046 433878 478102
rect 433934 478046 434002 478102
rect 434058 478046 434128 478102
rect 435498 478094 436118 489922
rect 439218 532350 439838 540962
rect 439218 532294 439314 532350
rect 439370 532294 439438 532350
rect 439494 532294 439562 532350
rect 439618 532294 439686 532350
rect 439742 532294 439838 532350
rect 439218 532226 439838 532294
rect 439218 532170 439314 532226
rect 439370 532170 439438 532226
rect 439494 532170 439562 532226
rect 439618 532170 439686 532226
rect 439742 532170 439838 532226
rect 439218 532102 439838 532170
rect 439218 532046 439314 532102
rect 439370 532046 439438 532102
rect 439494 532046 439562 532102
rect 439618 532046 439686 532102
rect 439742 532046 439838 532102
rect 439218 531978 439838 532046
rect 439218 531922 439314 531978
rect 439370 531922 439438 531978
rect 439494 531922 439562 531978
rect 439618 531922 439686 531978
rect 439742 531922 439838 531978
rect 439218 514350 439838 531922
rect 439218 514294 439314 514350
rect 439370 514294 439438 514350
rect 439494 514294 439562 514350
rect 439618 514294 439686 514350
rect 439742 514294 439838 514350
rect 439218 514226 439838 514294
rect 439218 514170 439314 514226
rect 439370 514170 439438 514226
rect 439494 514170 439562 514226
rect 439618 514170 439686 514226
rect 439742 514170 439838 514226
rect 439218 514102 439838 514170
rect 439218 514046 439314 514102
rect 439370 514046 439438 514102
rect 439494 514046 439562 514102
rect 439618 514046 439686 514102
rect 439742 514046 439838 514102
rect 439218 513978 439838 514046
rect 439218 513922 439314 513978
rect 439370 513922 439438 513978
rect 439494 513922 439562 513978
rect 439618 513922 439686 513978
rect 439742 513922 439838 513978
rect 439218 496350 439838 513922
rect 455308 510132 455364 542444
rect 456092 513156 456148 547708
rect 456876 530180 456932 530190
rect 456876 526596 456932 530124
rect 456876 526530 456932 526540
rect 456988 514836 457044 548492
rect 458668 547764 458724 551852
rect 458668 547698 458724 547708
rect 458668 546532 458724 546542
rect 456988 514770 457044 514780
rect 457772 546084 457828 546094
rect 456092 513090 456148 513100
rect 457772 512596 457828 546028
rect 457772 512530 457828 512540
rect 455308 510066 455364 510076
rect 458668 506772 458724 546476
rect 458780 546084 458836 553196
rect 459004 551236 459060 551246
rect 458780 546018 458836 546028
rect 458892 549220 458948 549230
rect 458668 506706 458724 506716
rect 458780 545188 458836 545198
rect 458780 505092 458836 545132
rect 458892 511700 458948 549164
rect 459004 520100 459060 551180
rect 459004 520034 459060 520044
rect 461132 548548 461188 548558
rect 461132 518756 461188 548492
rect 466218 544350 466838 561922
rect 466218 544294 466314 544350
rect 466370 544294 466438 544350
rect 466494 544294 466562 544350
rect 466618 544294 466686 544350
rect 466742 544294 466838 544350
rect 466218 544226 466838 544294
rect 466218 544170 466314 544226
rect 466370 544170 466438 544226
rect 466494 544170 466562 544226
rect 466618 544170 466686 544226
rect 466742 544170 466838 544226
rect 466218 544102 466838 544170
rect 466218 544046 466314 544102
rect 466370 544046 466438 544102
rect 466494 544046 466562 544102
rect 466618 544046 466686 544102
rect 466742 544046 466838 544102
rect 466218 543978 466838 544046
rect 466218 543922 466314 543978
rect 466370 543922 466438 543978
rect 466494 543922 466562 543978
rect 466618 543922 466686 543978
rect 466742 543922 466838 543978
rect 461132 518690 461188 518700
rect 464492 536788 464548 536798
rect 464492 517076 464548 536732
rect 464492 517010 464548 517020
rect 466218 526350 466838 543922
rect 466218 526294 466314 526350
rect 466370 526294 466438 526350
rect 466494 526294 466562 526350
rect 466618 526294 466686 526350
rect 466742 526294 466838 526350
rect 466218 526226 466838 526294
rect 466218 526170 466314 526226
rect 466370 526170 466438 526226
rect 466494 526170 466562 526226
rect 466618 526170 466686 526226
rect 466742 526170 466838 526226
rect 466218 526102 466838 526170
rect 466218 526046 466314 526102
rect 466370 526046 466438 526102
rect 466494 526046 466562 526102
rect 466618 526046 466686 526102
rect 466742 526046 466838 526102
rect 466218 525978 466838 526046
rect 466218 525922 466314 525978
rect 466370 525922 466438 525978
rect 466494 525922 466562 525978
rect 466618 525922 466686 525978
rect 466742 525922 466838 525978
rect 458892 511634 458948 511644
rect 458780 505026 458836 505036
rect 466218 508350 466838 525922
rect 466218 508294 466314 508350
rect 466370 508294 466438 508350
rect 466494 508294 466562 508350
rect 466618 508294 466686 508350
rect 466742 508294 466838 508350
rect 466218 508226 466838 508294
rect 466218 508170 466314 508226
rect 466370 508170 466438 508226
rect 466494 508170 466562 508226
rect 466618 508170 466686 508226
rect 466742 508170 466838 508226
rect 466218 508102 466838 508170
rect 466218 508046 466314 508102
rect 466370 508046 466438 508102
rect 466494 508046 466562 508102
rect 466618 508046 466686 508102
rect 466742 508046 466838 508102
rect 466218 507978 466838 508046
rect 466218 507922 466314 507978
rect 466370 507922 466438 507978
rect 466494 507922 466562 507978
rect 466618 507922 466686 507978
rect 466742 507922 466838 507978
rect 439218 496294 439314 496350
rect 439370 496294 439438 496350
rect 439494 496294 439562 496350
rect 439618 496294 439686 496350
rect 439742 496294 439838 496350
rect 439218 496226 439838 496294
rect 439218 496170 439314 496226
rect 439370 496170 439438 496226
rect 439494 496170 439562 496226
rect 439618 496170 439686 496226
rect 439742 496170 439838 496226
rect 439218 496102 439838 496170
rect 439218 496046 439314 496102
rect 439370 496046 439438 496102
rect 439494 496046 439562 496102
rect 439618 496046 439686 496102
rect 439742 496046 439838 496102
rect 439218 495978 439838 496046
rect 439218 495922 439314 495978
rect 439370 495922 439438 495978
rect 439494 495922 439562 495978
rect 439618 495922 439686 495978
rect 439742 495922 439838 495978
rect 439218 478350 439838 495922
rect 459228 493444 459284 493454
rect 449168 490350 449488 490384
rect 449168 490294 449238 490350
rect 449294 490294 449362 490350
rect 449418 490294 449488 490350
rect 449168 490226 449488 490294
rect 449168 490170 449238 490226
rect 449294 490170 449362 490226
rect 449418 490170 449488 490226
rect 449168 490102 449488 490170
rect 449168 490046 449238 490102
rect 449294 490046 449362 490102
rect 449418 490046 449488 490102
rect 449168 489978 449488 490046
rect 449168 489922 449238 489978
rect 449294 489922 449362 489978
rect 449418 489922 449488 489978
rect 449168 489888 449488 489922
rect 458668 483364 458724 483374
rect 456988 482020 457044 482030
rect 439218 478294 439314 478350
rect 439370 478294 439438 478350
rect 439494 478294 439562 478350
rect 439618 478294 439686 478350
rect 439742 478294 439838 478350
rect 439218 478226 439838 478294
rect 439218 478170 439314 478226
rect 439370 478170 439438 478226
rect 439494 478170 439562 478226
rect 439618 478170 439686 478226
rect 439742 478170 439838 478226
rect 439218 478102 439838 478170
rect 433808 477978 434128 478046
rect 433808 477922 433878 477978
rect 433934 477922 434002 477978
rect 434058 477922 434128 477978
rect 433808 477888 434128 477922
rect 439218 478046 439314 478102
rect 439370 478046 439438 478102
rect 439494 478046 439562 478102
rect 439618 478046 439686 478102
rect 439742 478046 439838 478102
rect 439218 477978 439838 478046
rect 439218 477922 439314 477978
rect 439370 477922 439438 477978
rect 439494 477922 439562 477978
rect 439618 477922 439686 477978
rect 439742 477922 439838 477978
rect 418448 472350 418768 472384
rect 418448 472294 418518 472350
rect 418574 472294 418642 472350
rect 418698 472294 418768 472350
rect 418448 472226 418768 472294
rect 418448 472170 418518 472226
rect 418574 472170 418642 472226
rect 418698 472170 418768 472226
rect 418448 472102 418768 472170
rect 418448 472046 418518 472102
rect 418574 472046 418642 472102
rect 418698 472046 418768 472102
rect 418448 471978 418768 472046
rect 418448 471922 418518 471978
rect 418574 471922 418642 471978
rect 418698 471922 418768 471978
rect 418448 471888 418768 471922
rect 435498 472060 436118 472114
rect 435498 472004 435594 472060
rect 435650 472004 435718 472060
rect 435774 472004 435842 472060
rect 435898 472004 435966 472060
rect 436022 472004 436118 472060
rect 435498 471936 436118 472004
rect 435498 471880 435594 471936
rect 435650 471880 435718 471936
rect 435774 471880 435842 471936
rect 435898 471880 435966 471936
rect 436022 471880 436118 471936
rect 433808 460350 434128 460384
rect 433808 460294 433878 460350
rect 433934 460294 434002 460350
rect 434058 460294 434128 460350
rect 433808 460226 434128 460294
rect 433808 460170 433878 460226
rect 433934 460170 434002 460226
rect 434058 460170 434128 460226
rect 433808 460102 434128 460170
rect 433808 460046 433878 460102
rect 433934 460046 434002 460102
rect 434058 460046 434128 460102
rect 433808 459978 434128 460046
rect 433808 459922 433878 459978
rect 433934 459922 434002 459978
rect 434058 459922 434128 459978
rect 433808 459888 434128 459922
rect 411180 456306 411236 456316
rect 410956 446226 411012 446236
rect 435498 454350 436118 471880
rect 435498 454294 435594 454350
rect 435650 454294 435718 454350
rect 435774 454294 435842 454350
rect 435898 454294 435966 454350
rect 436022 454294 436118 454350
rect 435498 454226 436118 454294
rect 435498 454170 435594 454226
rect 435650 454170 435718 454226
rect 435774 454170 435842 454226
rect 435898 454170 435966 454226
rect 436022 454170 436118 454226
rect 435498 454102 436118 454170
rect 435498 454046 435594 454102
rect 435650 454046 435718 454102
rect 435774 454046 435842 454102
rect 435898 454046 435966 454102
rect 436022 454046 436118 454102
rect 435498 453978 436118 454046
rect 435498 453922 435594 453978
rect 435650 453922 435718 453978
rect 435774 453922 435842 453978
rect 435898 453922 435966 453978
rect 436022 453922 436118 453978
rect 408498 442294 408594 442350
rect 408650 442294 408718 442350
rect 408774 442294 408842 442350
rect 408898 442294 408966 442350
rect 409022 442294 409118 442350
rect 408498 442226 409118 442294
rect 408498 442170 408594 442226
rect 408650 442170 408718 442226
rect 408774 442170 408842 442226
rect 408898 442170 408966 442226
rect 409022 442170 409118 442226
rect 408498 442102 409118 442170
rect 408498 442046 408594 442102
rect 408650 442046 408718 442102
rect 408774 442046 408842 442102
rect 408898 442046 408966 442102
rect 409022 442046 409118 442102
rect 408498 441978 409118 442046
rect 408498 441922 408594 441978
rect 408650 441922 408718 441978
rect 408774 441922 408842 441978
rect 408898 441922 408966 441978
rect 409022 441922 409118 441978
rect 408498 424350 409118 441922
rect 408498 424294 408594 424350
rect 408650 424294 408718 424350
rect 408774 424294 408842 424350
rect 408898 424294 408966 424350
rect 409022 424294 409118 424350
rect 408498 424226 409118 424294
rect 408498 424170 408594 424226
rect 408650 424170 408718 424226
rect 408774 424170 408842 424226
rect 408898 424170 408966 424226
rect 409022 424170 409118 424226
rect 408498 424102 409118 424170
rect 408498 424046 408594 424102
rect 408650 424046 408718 424102
rect 408774 424046 408842 424102
rect 408898 424046 408966 424102
rect 409022 424046 409118 424102
rect 408498 423978 409118 424046
rect 408498 423922 408594 423978
rect 408650 423922 408718 423978
rect 408774 423922 408842 423978
rect 408898 423922 408966 423978
rect 409022 423922 409118 423978
rect 408498 406350 409118 423922
rect 435498 436350 436118 453922
rect 435498 436294 435594 436350
rect 435650 436294 435718 436350
rect 435774 436294 435842 436350
rect 435898 436294 435966 436350
rect 436022 436294 436118 436350
rect 435498 436226 436118 436294
rect 435498 436170 435594 436226
rect 435650 436170 435718 436226
rect 435774 436170 435842 436226
rect 435898 436170 435966 436226
rect 436022 436170 436118 436226
rect 435498 436102 436118 436170
rect 435498 436046 435594 436102
rect 435650 436046 435718 436102
rect 435774 436046 435842 436102
rect 435898 436046 435966 436102
rect 436022 436046 436118 436102
rect 435498 435978 436118 436046
rect 435498 435922 435594 435978
rect 435650 435922 435718 435978
rect 435774 435922 435842 435978
rect 435898 435922 435966 435978
rect 436022 435922 436118 435978
rect 408498 406294 408594 406350
rect 408650 406294 408718 406350
rect 408774 406294 408842 406350
rect 408898 406294 408966 406350
rect 409022 406294 409118 406350
rect 408498 406226 409118 406294
rect 408498 406170 408594 406226
rect 408650 406170 408718 406226
rect 408774 406170 408842 406226
rect 408898 406170 408966 406226
rect 409022 406170 409118 406226
rect 408498 406102 409118 406170
rect 404778 400294 404874 400350
rect 404930 400294 404998 400350
rect 405054 400294 405122 400350
rect 405178 400294 405246 400350
rect 405302 400294 405398 400350
rect 404778 400226 405398 400294
rect 404778 400170 404874 400226
rect 404930 400170 404998 400226
rect 405054 400170 405122 400226
rect 405178 400170 405246 400226
rect 405302 400170 405398 400226
rect 404778 400102 405398 400170
rect 404778 400046 404874 400102
rect 404930 400046 404998 400102
rect 405054 400046 405122 400102
rect 405178 400046 405246 400102
rect 405302 400046 405398 400102
rect 404778 399978 405398 400046
rect 404778 399922 404874 399978
rect 404930 399922 404998 399978
rect 405054 399922 405122 399978
rect 405178 399922 405246 399978
rect 405302 399922 405398 399978
rect 404778 382350 405398 399922
rect 406588 406084 406644 406094
rect 406588 399718 406644 406028
rect 406588 399652 406644 399662
rect 408498 406046 408594 406102
rect 408650 406046 408718 406102
rect 408774 406046 408842 406102
rect 408898 406046 408966 406102
rect 409022 406046 409118 406102
rect 408498 405978 409118 406046
rect 408498 405922 408594 405978
rect 408650 405922 408718 405978
rect 408774 405922 408842 405978
rect 408898 405922 408966 405978
rect 409022 405922 409118 405978
rect 404778 382294 404874 382350
rect 404930 382294 404998 382350
rect 405054 382294 405122 382350
rect 405178 382294 405246 382350
rect 405302 382294 405398 382350
rect 404778 382226 405398 382294
rect 404778 382170 404874 382226
rect 404930 382170 404998 382226
rect 405054 382170 405122 382226
rect 405178 382170 405246 382226
rect 405302 382170 405398 382226
rect 404778 382102 405398 382170
rect 404778 382046 404874 382102
rect 404930 382046 404998 382102
rect 405054 382046 405122 382102
rect 405178 382046 405246 382102
rect 405302 382046 405398 382102
rect 404778 381978 405398 382046
rect 404778 381922 404874 381978
rect 404930 381922 404998 381978
rect 405054 381922 405122 381978
rect 405178 381922 405246 381978
rect 405302 381922 405398 381978
rect 398972 366930 399028 366940
rect 396508 365474 396564 365484
rect 394828 362002 394884 362012
rect 404778 364350 405398 381922
rect 404778 364294 404874 364350
rect 404930 364294 404998 364350
rect 405054 364294 405122 364350
rect 405178 364294 405246 364350
rect 405302 364294 405398 364350
rect 404778 364226 405398 364294
rect 404778 364170 404874 364226
rect 404930 364170 404998 364226
rect 405054 364170 405122 364226
rect 405178 364170 405246 364226
rect 405302 364170 405398 364226
rect 404778 364102 405398 364170
rect 404778 364046 404874 364102
rect 404930 364046 404998 364102
rect 405054 364046 405122 364102
rect 405178 364046 405246 364102
rect 405302 364046 405398 364102
rect 404778 363978 405398 364046
rect 404778 363922 404874 363978
rect 404930 363922 404998 363978
rect 405054 363922 405122 363978
rect 405178 363922 405246 363978
rect 405302 363922 405398 363978
rect 392252 361890 392308 361900
rect 377778 352294 377874 352350
rect 377930 352294 377998 352350
rect 378054 352294 378122 352350
rect 378178 352294 378246 352350
rect 378302 352294 378398 352350
rect 377778 352226 378398 352294
rect 377778 352170 377874 352226
rect 377930 352170 377998 352226
rect 378054 352170 378122 352226
rect 378178 352170 378246 352226
rect 378302 352170 378398 352226
rect 377778 352102 378398 352170
rect 377778 352046 377874 352102
rect 377930 352046 377998 352102
rect 378054 352046 378122 352102
rect 378178 352046 378246 352102
rect 378302 352046 378398 352102
rect 377778 351978 378398 352046
rect 377778 351922 377874 351978
rect 377930 351922 377998 351978
rect 378054 351922 378122 351978
rect 378178 351922 378246 351978
rect 378302 351922 378398 351978
rect 377778 334350 378398 351922
rect 393372 349972 393428 349982
rect 393372 349318 393428 349916
rect 393372 349252 393428 349262
rect 394828 348598 394884 348608
rect 387168 346350 387488 346384
rect 387168 346294 387238 346350
rect 387294 346294 387362 346350
rect 387418 346294 387488 346350
rect 387168 346226 387488 346294
rect 387168 346170 387238 346226
rect 387294 346170 387362 346226
rect 387418 346170 387488 346226
rect 387168 346102 387488 346170
rect 387168 346046 387238 346102
rect 387294 346046 387362 346102
rect 387418 346046 387488 346102
rect 387168 345978 387488 346046
rect 387168 345922 387238 345978
rect 387294 345922 387362 345978
rect 387418 345922 387488 345978
rect 387168 345888 387488 345922
rect 394828 344278 394884 348542
rect 394828 344212 394884 344222
rect 404778 346350 405398 363922
rect 404778 346294 404874 346350
rect 404930 346294 404998 346350
rect 405054 346294 405122 346350
rect 405178 346294 405246 346350
rect 405302 346294 405398 346350
rect 404778 346226 405398 346294
rect 404778 346170 404874 346226
rect 404930 346170 404998 346226
rect 405054 346170 405122 346226
rect 405178 346170 405246 346226
rect 405302 346170 405398 346226
rect 404778 346102 405398 346170
rect 404778 346046 404874 346102
rect 404930 346046 404998 346102
rect 405054 346046 405122 346102
rect 405178 346046 405246 346102
rect 405302 346046 405398 346102
rect 404778 345978 405398 346046
rect 404778 345922 404874 345978
rect 404930 345922 404998 345978
rect 405054 345922 405122 345978
rect 405178 345922 405246 345978
rect 405302 345922 405398 345978
rect 394044 340452 394100 340462
rect 393372 339780 393428 339790
rect 393372 339238 393428 339724
rect 393372 339172 393428 339182
rect 393484 337092 393540 337102
rect 377778 334294 377874 334350
rect 377930 334294 377998 334350
rect 378054 334294 378122 334350
rect 378178 334294 378246 334350
rect 378302 334294 378398 334350
rect 377778 334226 378398 334294
rect 377778 334170 377874 334226
rect 377930 334170 377998 334226
rect 378054 334170 378122 334226
rect 378178 334170 378246 334226
rect 378302 334170 378398 334226
rect 377778 334102 378398 334170
rect 377778 334046 377874 334102
rect 377930 334046 377998 334102
rect 378054 334046 378122 334102
rect 378178 334046 378246 334102
rect 378302 334046 378398 334102
rect 377778 333978 378398 334046
rect 377778 333922 377874 333978
rect 377930 333922 377998 333978
rect 378054 333922 378122 333978
rect 378178 333922 378246 333978
rect 378302 333922 378398 333978
rect 377778 316350 378398 333922
rect 393148 336358 393204 336368
rect 393148 331858 393204 336302
rect 393372 333732 393428 333742
rect 393372 332578 393428 333676
rect 393484 333658 393540 337036
rect 393484 333592 393540 333602
rect 393372 332512 393428 332522
rect 393148 331792 393204 331802
rect 393932 332276 393988 332286
rect 393260 329588 393316 329598
rect 393260 329518 393316 329532
rect 393260 329452 393316 329462
rect 387168 328350 387488 328384
rect 387168 328294 387238 328350
rect 387294 328294 387362 328350
rect 387418 328294 387488 328350
rect 387168 328226 387488 328294
rect 387168 328170 387238 328226
rect 387294 328170 387362 328226
rect 387418 328170 387488 328226
rect 387168 328102 387488 328170
rect 387168 328046 387238 328102
rect 387294 328046 387362 328102
rect 387418 328046 387488 328102
rect 387168 327978 387488 328046
rect 387168 327922 387238 327978
rect 387294 327922 387362 327978
rect 387418 327922 387488 327978
rect 387168 327888 387488 327922
rect 377778 316294 377874 316350
rect 377930 316294 377998 316350
rect 378054 316294 378122 316350
rect 378178 316294 378246 316350
rect 378302 316294 378398 316350
rect 377778 316226 378398 316294
rect 377778 316170 377874 316226
rect 377930 316170 377998 316226
rect 378054 316170 378122 316226
rect 378178 316170 378246 316226
rect 378302 316170 378398 316226
rect 377778 316102 378398 316170
rect 377778 316046 377874 316102
rect 377930 316046 377998 316102
rect 378054 316046 378122 316102
rect 378178 316046 378246 316102
rect 378302 316046 378398 316102
rect 377778 315978 378398 316046
rect 377778 315922 377874 315978
rect 377930 315922 377998 315978
rect 378054 315922 378122 315978
rect 378178 315922 378246 315978
rect 378302 315922 378398 315978
rect 377778 298350 378398 315922
rect 393932 307636 393988 332220
rect 394044 327358 394100 340396
rect 404460 339778 404516 339788
rect 394828 338518 394884 338528
rect 394828 337618 394884 338462
rect 394828 337552 394884 337562
rect 396508 337978 396564 337988
rect 396508 336898 396564 337922
rect 396508 336832 396564 336842
rect 396508 336420 396564 336430
rect 394828 336084 394884 336094
rect 394828 332578 394884 336028
rect 394828 332512 394884 332522
rect 394940 334292 394996 334302
rect 394940 330778 394996 334236
rect 394940 330712 394996 330722
rect 395612 330932 395668 330942
rect 394828 329700 394884 329710
rect 394828 327538 394884 329644
rect 394828 327472 394884 327482
rect 394044 327292 394100 327302
rect 393932 307570 393988 307580
rect 395612 299236 395668 330876
rect 396508 330932 396564 336364
rect 399756 336178 399812 336188
rect 399756 334292 399812 336122
rect 404460 335098 404516 339722
rect 404572 337798 404628 337808
rect 404572 335998 404628 337742
rect 404572 335932 404628 335942
rect 404460 335032 404516 335042
rect 399756 334226 399812 334236
rect 403228 334738 403284 334748
rect 396508 330866 396564 330876
rect 396844 332724 396900 332734
rect 396844 302596 396900 332668
rect 403228 330058 403284 334682
rect 403228 329992 403284 330002
rect 404778 328350 405398 345922
rect 408498 388350 409118 405922
rect 410732 421540 410788 421550
rect 410732 394498 410788 421484
rect 418448 418350 418768 418384
rect 418448 418294 418518 418350
rect 418574 418294 418642 418350
rect 418698 418294 418768 418350
rect 418448 418226 418768 418294
rect 418448 418170 418518 418226
rect 418574 418170 418642 418226
rect 418698 418170 418768 418226
rect 418448 418102 418768 418170
rect 418448 418046 418518 418102
rect 418574 418046 418642 418102
rect 418698 418046 418768 418102
rect 418448 417978 418768 418046
rect 418448 417922 418518 417978
rect 418574 417922 418642 417978
rect 418698 417922 418768 417978
rect 418448 417888 418768 417922
rect 435498 418350 436118 435922
rect 439218 460350 439838 477922
rect 455308 480004 455364 480014
rect 449168 472350 449488 472384
rect 449168 472294 449238 472350
rect 449294 472294 449362 472350
rect 449418 472294 449488 472350
rect 449168 472226 449488 472294
rect 449168 472170 449238 472226
rect 449294 472170 449362 472226
rect 449418 472170 449488 472226
rect 449168 472102 449488 472170
rect 449168 472046 449238 472102
rect 449294 472046 449362 472102
rect 449418 472046 449488 472102
rect 449168 471978 449488 472046
rect 449168 471922 449238 471978
rect 449294 471922 449362 471978
rect 449418 471922 449488 471978
rect 449168 471888 449488 471922
rect 439218 460294 439314 460350
rect 439370 460294 439438 460350
rect 439494 460294 439562 460350
rect 439618 460294 439686 460350
rect 439742 460294 439838 460350
rect 439218 460226 439838 460294
rect 439218 460170 439314 460226
rect 439370 460170 439438 460226
rect 439494 460170 439562 460226
rect 439618 460170 439686 460226
rect 439742 460170 439838 460226
rect 439218 460102 439838 460170
rect 439218 460046 439314 460102
rect 439370 460046 439438 460102
rect 439494 460046 439562 460102
rect 439618 460046 439686 460102
rect 439742 460046 439838 460102
rect 439218 459978 439838 460046
rect 439218 459922 439314 459978
rect 439370 459922 439438 459978
rect 439494 459922 439562 459978
rect 439618 459922 439686 459978
rect 439742 459922 439838 459978
rect 439218 442350 439838 459922
rect 439218 442294 439314 442350
rect 439370 442294 439438 442350
rect 439494 442294 439562 442350
rect 439618 442294 439686 442350
rect 439742 442294 439838 442350
rect 439218 442226 439838 442294
rect 439218 442170 439314 442226
rect 439370 442170 439438 442226
rect 439494 442170 439562 442226
rect 439618 442170 439686 442226
rect 439742 442170 439838 442226
rect 439218 442102 439838 442170
rect 439218 442046 439314 442102
rect 439370 442046 439438 442102
rect 439494 442046 439562 442102
rect 439618 442046 439686 442102
rect 439742 442046 439838 442102
rect 439218 441978 439838 442046
rect 439218 441922 439314 441978
rect 439370 441922 439438 441978
rect 439494 441922 439562 441978
rect 439618 441922 439686 441978
rect 439742 441922 439838 441978
rect 436828 427028 436884 427038
rect 436828 426244 436884 426972
rect 436828 426178 436884 426188
rect 438172 427028 438228 427038
rect 438172 426244 438228 426972
rect 438172 426178 438228 426188
rect 435498 418294 435594 418350
rect 435650 418294 435718 418350
rect 435774 418294 435842 418350
rect 435898 418294 435966 418350
rect 436022 418294 436118 418350
rect 435498 418226 436118 418294
rect 435498 418170 435594 418226
rect 435650 418170 435718 418226
rect 435774 418170 435842 418226
rect 435898 418170 435966 418226
rect 436022 418170 436118 418226
rect 435498 418102 436118 418170
rect 435498 418046 435594 418102
rect 435650 418046 435718 418102
rect 435774 418046 435842 418102
rect 435898 418046 435966 418102
rect 436022 418046 436118 418102
rect 435498 417978 436118 418046
rect 435498 417922 435594 417978
rect 435650 417922 435718 417978
rect 435774 417922 435842 417978
rect 435898 417922 435966 417978
rect 436022 417922 436118 417978
rect 414092 413758 414148 413768
rect 411516 411598 411572 411608
rect 411516 411460 411572 411542
rect 411516 411394 411572 411404
rect 411180 407428 411236 407438
rect 411068 406756 411124 406766
rect 411068 402418 411124 406700
rect 411180 406738 411236 407372
rect 411180 406672 411236 406682
rect 411068 402352 411124 402362
rect 411180 404740 411236 404750
rect 411180 402388 411236 404684
rect 414092 402958 414148 413702
rect 414652 413398 414708 413408
rect 414652 411460 414708 413342
rect 414652 411394 414708 411404
rect 428876 412138 428932 412148
rect 428876 407458 428932 412082
rect 435498 409918 436118 417922
rect 439218 424350 439838 441922
rect 455308 427588 455364 479948
rect 455420 479332 455476 479342
rect 455420 432628 455476 479276
rect 455532 475972 455588 475982
rect 455532 455476 455588 475916
rect 455532 455410 455588 455420
rect 456092 474516 456148 474526
rect 456092 454356 456148 474460
rect 456092 454290 456148 454300
rect 455420 432562 455476 432572
rect 455308 427522 455364 427532
rect 456988 424676 457044 481964
rect 457324 477988 457380 477998
rect 457212 474068 457268 474078
rect 457100 473956 457156 473966
rect 457100 427476 457156 473900
rect 457212 454916 457268 474012
rect 457324 457044 457380 477932
rect 457324 456978 457380 456988
rect 457772 475524 457828 475534
rect 457212 454850 457268 454860
rect 457772 451556 457828 475468
rect 458668 475524 458724 483308
rect 458668 475458 458724 475468
rect 458780 482692 458836 482702
rect 457772 451490 457828 451500
rect 458780 447860 458836 482636
rect 459004 481348 459060 481358
rect 458892 480676 458948 480686
rect 458892 456148 458948 480620
rect 459004 458052 459060 481292
rect 459116 478660 459172 478670
rect 459116 458164 459172 478604
rect 459116 458098 459172 458108
rect 459004 457986 459060 457996
rect 459228 456260 459284 493388
rect 466218 490350 466838 507922
rect 466218 490294 466314 490350
rect 466370 490294 466438 490350
rect 466494 490294 466562 490350
rect 466618 490294 466686 490350
rect 466742 490294 466838 490350
rect 466218 490226 466838 490294
rect 466218 490170 466314 490226
rect 466370 490170 466438 490226
rect 466494 490170 466562 490226
rect 466618 490170 466686 490226
rect 466742 490170 466838 490226
rect 466218 490102 466838 490170
rect 466218 490046 466314 490102
rect 466370 490046 466438 490102
rect 466494 490046 466562 490102
rect 466618 490046 466686 490102
rect 466742 490046 466838 490102
rect 466218 489978 466838 490046
rect 466218 489922 466314 489978
rect 466370 489922 466438 489978
rect 466494 489922 466562 489978
rect 466618 489922 466686 489978
rect 466742 489922 466838 489978
rect 459228 456194 459284 456204
rect 461132 481460 461188 481470
rect 458892 456082 458948 456092
rect 458780 447794 458836 447804
rect 461132 430836 461188 481404
rect 462812 481348 462868 481358
rect 462812 462898 462868 481292
rect 462812 462832 462868 462842
rect 466218 472350 466838 489922
rect 469938 598172 470558 598268
rect 469938 598116 470034 598172
rect 470090 598116 470158 598172
rect 470214 598116 470282 598172
rect 470338 598116 470406 598172
rect 470462 598116 470558 598172
rect 469938 598048 470558 598116
rect 469938 597992 470034 598048
rect 470090 597992 470158 598048
rect 470214 597992 470282 598048
rect 470338 597992 470406 598048
rect 470462 597992 470558 598048
rect 469938 597924 470558 597992
rect 469938 597868 470034 597924
rect 470090 597868 470158 597924
rect 470214 597868 470282 597924
rect 470338 597868 470406 597924
rect 470462 597868 470558 597924
rect 469938 597800 470558 597868
rect 469938 597744 470034 597800
rect 470090 597744 470158 597800
rect 470214 597744 470282 597800
rect 470338 597744 470406 597800
rect 470462 597744 470558 597800
rect 469938 586350 470558 597744
rect 469938 586294 470034 586350
rect 470090 586294 470158 586350
rect 470214 586294 470282 586350
rect 470338 586294 470406 586350
rect 470462 586294 470558 586350
rect 469938 586226 470558 586294
rect 469938 586170 470034 586226
rect 470090 586170 470158 586226
rect 470214 586170 470282 586226
rect 470338 586170 470406 586226
rect 470462 586170 470558 586226
rect 469938 586102 470558 586170
rect 469938 586046 470034 586102
rect 470090 586046 470158 586102
rect 470214 586046 470282 586102
rect 470338 586046 470406 586102
rect 470462 586046 470558 586102
rect 469938 585978 470558 586046
rect 469938 585922 470034 585978
rect 470090 585922 470158 585978
rect 470214 585922 470282 585978
rect 470338 585922 470406 585978
rect 470462 585922 470558 585978
rect 469938 568350 470558 585922
rect 469938 568294 470034 568350
rect 470090 568294 470158 568350
rect 470214 568294 470282 568350
rect 470338 568294 470406 568350
rect 470462 568294 470558 568350
rect 469938 568226 470558 568294
rect 469938 568170 470034 568226
rect 470090 568170 470158 568226
rect 470214 568170 470282 568226
rect 470338 568170 470406 568226
rect 470462 568170 470558 568226
rect 469938 568102 470558 568170
rect 469938 568046 470034 568102
rect 470090 568046 470158 568102
rect 470214 568046 470282 568102
rect 470338 568046 470406 568102
rect 470462 568046 470558 568102
rect 469938 567978 470558 568046
rect 469938 567922 470034 567978
rect 470090 567922 470158 567978
rect 470214 567922 470282 567978
rect 470338 567922 470406 567978
rect 470462 567922 470558 567978
rect 469938 550350 470558 567922
rect 496938 597212 497558 598268
rect 496938 597156 497034 597212
rect 497090 597156 497158 597212
rect 497214 597156 497282 597212
rect 497338 597156 497406 597212
rect 497462 597156 497558 597212
rect 496938 597088 497558 597156
rect 496938 597032 497034 597088
rect 497090 597032 497158 597088
rect 497214 597032 497282 597088
rect 497338 597032 497406 597088
rect 497462 597032 497558 597088
rect 496938 596964 497558 597032
rect 496938 596908 497034 596964
rect 497090 596908 497158 596964
rect 497214 596908 497282 596964
rect 497338 596908 497406 596964
rect 497462 596908 497558 596964
rect 496938 596840 497558 596908
rect 496938 596784 497034 596840
rect 497090 596784 497158 596840
rect 497214 596784 497282 596840
rect 497338 596784 497406 596840
rect 497462 596784 497558 596840
rect 496938 580350 497558 596784
rect 496938 580294 497034 580350
rect 497090 580294 497158 580350
rect 497214 580294 497282 580350
rect 497338 580294 497406 580350
rect 497462 580294 497558 580350
rect 496938 580226 497558 580294
rect 496938 580170 497034 580226
rect 497090 580170 497158 580226
rect 497214 580170 497282 580226
rect 497338 580170 497406 580226
rect 497462 580170 497558 580226
rect 496938 580102 497558 580170
rect 496938 580046 497034 580102
rect 497090 580046 497158 580102
rect 497214 580046 497282 580102
rect 497338 580046 497406 580102
rect 497462 580046 497558 580102
rect 496938 579978 497558 580046
rect 496938 579922 497034 579978
rect 497090 579922 497158 579978
rect 497214 579922 497282 579978
rect 497338 579922 497406 579978
rect 497462 579922 497558 579978
rect 480448 562350 480768 562384
rect 480448 562294 480518 562350
rect 480574 562294 480642 562350
rect 480698 562294 480768 562350
rect 480448 562226 480768 562294
rect 480448 562170 480518 562226
rect 480574 562170 480642 562226
rect 480698 562170 480768 562226
rect 480448 562102 480768 562170
rect 480448 562046 480518 562102
rect 480574 562046 480642 562102
rect 480698 562046 480768 562102
rect 480448 561978 480768 562046
rect 480448 561922 480518 561978
rect 480574 561922 480642 561978
rect 480698 561922 480768 561978
rect 480448 561888 480768 561922
rect 496938 562350 497558 579922
rect 496938 562294 497034 562350
rect 497090 562294 497158 562350
rect 497214 562294 497282 562350
rect 497338 562294 497406 562350
rect 497462 562294 497558 562350
rect 496938 562226 497558 562294
rect 496938 562170 497034 562226
rect 497090 562170 497158 562226
rect 497214 562170 497282 562226
rect 497338 562170 497406 562226
rect 497462 562170 497558 562226
rect 496938 562102 497558 562170
rect 496938 562046 497034 562102
rect 497090 562046 497158 562102
rect 497214 562046 497282 562102
rect 497338 562046 497406 562102
rect 497462 562046 497558 562102
rect 496938 561978 497558 562046
rect 496938 561922 497034 561978
rect 497090 561922 497158 561978
rect 497214 561922 497282 561978
rect 497338 561922 497406 561978
rect 497462 561922 497558 561978
rect 496938 557694 497558 561922
rect 500658 598172 501278 598268
rect 500658 598116 500754 598172
rect 500810 598116 500878 598172
rect 500934 598116 501002 598172
rect 501058 598116 501126 598172
rect 501182 598116 501278 598172
rect 500658 598048 501278 598116
rect 500658 597992 500754 598048
rect 500810 597992 500878 598048
rect 500934 597992 501002 598048
rect 501058 597992 501126 598048
rect 501182 597992 501278 598048
rect 500658 597924 501278 597992
rect 500658 597868 500754 597924
rect 500810 597868 500878 597924
rect 500934 597868 501002 597924
rect 501058 597868 501126 597924
rect 501182 597868 501278 597924
rect 500658 597800 501278 597868
rect 500658 597744 500754 597800
rect 500810 597744 500878 597800
rect 500934 597744 501002 597800
rect 501058 597744 501126 597800
rect 501182 597744 501278 597800
rect 500658 586350 501278 597744
rect 500658 586294 500754 586350
rect 500810 586294 500878 586350
rect 500934 586294 501002 586350
rect 501058 586294 501126 586350
rect 501182 586294 501278 586350
rect 500658 586226 501278 586294
rect 500658 586170 500754 586226
rect 500810 586170 500878 586226
rect 500934 586170 501002 586226
rect 501058 586170 501126 586226
rect 501182 586170 501278 586226
rect 500658 586102 501278 586170
rect 500658 586046 500754 586102
rect 500810 586046 500878 586102
rect 500934 586046 501002 586102
rect 501058 586046 501126 586102
rect 501182 586046 501278 586102
rect 500658 585978 501278 586046
rect 500658 585922 500754 585978
rect 500810 585922 500878 585978
rect 500934 585922 501002 585978
rect 501058 585922 501126 585978
rect 501182 585922 501278 585978
rect 500658 568350 501278 585922
rect 500658 568294 500754 568350
rect 500810 568294 500878 568350
rect 500934 568294 501002 568350
rect 501058 568294 501126 568350
rect 501182 568294 501278 568350
rect 500658 568226 501278 568294
rect 500658 568170 500754 568226
rect 500810 568170 500878 568226
rect 500934 568170 501002 568226
rect 501058 568170 501126 568226
rect 501182 568170 501278 568226
rect 500658 568102 501278 568170
rect 500658 568046 500754 568102
rect 500810 568046 500878 568102
rect 500934 568046 501002 568102
rect 501058 568046 501126 568102
rect 501182 568046 501278 568102
rect 500658 567978 501278 568046
rect 500658 567922 500754 567978
rect 500810 567922 500878 567978
rect 500934 567922 501002 567978
rect 501058 567922 501126 567978
rect 501182 567922 501278 567978
rect 500658 557694 501278 567922
rect 527658 597212 528278 598268
rect 527658 597156 527754 597212
rect 527810 597156 527878 597212
rect 527934 597156 528002 597212
rect 528058 597156 528126 597212
rect 528182 597156 528278 597212
rect 527658 597088 528278 597156
rect 527658 597032 527754 597088
rect 527810 597032 527878 597088
rect 527934 597032 528002 597088
rect 528058 597032 528126 597088
rect 528182 597032 528278 597088
rect 527658 596964 528278 597032
rect 527658 596908 527754 596964
rect 527810 596908 527878 596964
rect 527934 596908 528002 596964
rect 528058 596908 528126 596964
rect 528182 596908 528278 596964
rect 527658 596840 528278 596908
rect 527658 596784 527754 596840
rect 527810 596784 527878 596840
rect 527934 596784 528002 596840
rect 528058 596784 528126 596840
rect 528182 596784 528278 596840
rect 527658 580350 528278 596784
rect 527658 580294 527754 580350
rect 527810 580294 527878 580350
rect 527934 580294 528002 580350
rect 528058 580294 528126 580350
rect 528182 580294 528278 580350
rect 527658 580226 528278 580294
rect 527658 580170 527754 580226
rect 527810 580170 527878 580226
rect 527934 580170 528002 580226
rect 528058 580170 528126 580226
rect 528182 580170 528278 580226
rect 527658 580102 528278 580170
rect 527658 580046 527754 580102
rect 527810 580046 527878 580102
rect 527934 580046 528002 580102
rect 528058 580046 528126 580102
rect 528182 580046 528278 580102
rect 527658 579978 528278 580046
rect 527658 579922 527754 579978
rect 527810 579922 527878 579978
rect 527934 579922 528002 579978
rect 528058 579922 528126 579978
rect 528182 579922 528278 579978
rect 511168 562350 511488 562384
rect 511168 562294 511238 562350
rect 511294 562294 511362 562350
rect 511418 562294 511488 562350
rect 511168 562226 511488 562294
rect 511168 562170 511238 562226
rect 511294 562170 511362 562226
rect 511418 562170 511488 562226
rect 511168 562102 511488 562170
rect 511168 562046 511238 562102
rect 511294 562046 511362 562102
rect 511418 562046 511488 562102
rect 511168 561978 511488 562046
rect 511168 561922 511238 561978
rect 511294 561922 511362 561978
rect 511418 561922 511488 561978
rect 511168 561888 511488 561922
rect 527658 562350 528278 579922
rect 527658 562294 527754 562350
rect 527810 562294 527878 562350
rect 527934 562294 528002 562350
rect 528058 562294 528126 562350
rect 528182 562294 528278 562350
rect 527658 562226 528278 562294
rect 527658 562170 527754 562226
rect 527810 562170 527878 562226
rect 527934 562170 528002 562226
rect 528058 562170 528126 562226
rect 528182 562170 528278 562226
rect 527658 562102 528278 562170
rect 527658 562046 527754 562102
rect 527810 562046 527878 562102
rect 527934 562046 528002 562102
rect 528058 562046 528126 562102
rect 528182 562046 528278 562102
rect 527658 561978 528278 562046
rect 527658 561922 527754 561978
rect 527810 561922 527878 561978
rect 527934 561922 528002 561978
rect 528058 561922 528126 561978
rect 528182 561922 528278 561978
rect 473676 555268 473732 555278
rect 473676 555172 473732 555182
rect 476028 554820 476084 554830
rect 476028 554698 476084 554764
rect 476028 554632 476084 554642
rect 519036 554518 519092 554528
rect 473452 553924 473508 553934
rect 469938 550294 470034 550350
rect 470090 550294 470158 550350
rect 470214 550294 470282 550350
rect 470338 550294 470406 550350
rect 470462 550294 470558 550350
rect 469938 550226 470558 550294
rect 469938 550170 470034 550226
rect 470090 550170 470158 550226
rect 470214 550170 470282 550226
rect 470338 550170 470406 550226
rect 470462 550170 470558 550226
rect 469938 550102 470558 550170
rect 469938 550046 470034 550102
rect 470090 550046 470158 550102
rect 470214 550046 470282 550102
rect 470338 550046 470406 550102
rect 470462 550046 470558 550102
rect 469938 549978 470558 550046
rect 469938 549922 470034 549978
rect 470090 549922 470158 549978
rect 470214 549922 470282 549978
rect 470338 549922 470406 549978
rect 470462 549922 470558 549978
rect 469938 532350 470558 549922
rect 469938 532294 470034 532350
rect 470090 532294 470158 532350
rect 470214 532294 470282 532350
rect 470338 532294 470406 532350
rect 470462 532294 470558 532350
rect 469938 532226 470558 532294
rect 469938 532170 470034 532226
rect 470090 532170 470158 532226
rect 470214 532170 470282 532226
rect 470338 532170 470406 532226
rect 470462 532170 470558 532226
rect 469938 532102 470558 532170
rect 469938 532046 470034 532102
rect 470090 532046 470158 532102
rect 470214 532046 470282 532102
rect 470338 532046 470406 532102
rect 470462 532046 470558 532102
rect 469938 531978 470558 532046
rect 469938 531922 470034 531978
rect 470090 531922 470158 531978
rect 470214 531922 470282 531978
rect 470338 531922 470406 531978
rect 470462 531922 470558 531978
rect 469938 514350 470558 531922
rect 469938 514294 470034 514350
rect 470090 514294 470158 514350
rect 470214 514294 470282 514350
rect 470338 514294 470406 514350
rect 470462 514294 470558 514350
rect 469938 514226 470558 514294
rect 469938 514170 470034 514226
rect 470090 514170 470158 514226
rect 470214 514170 470282 514226
rect 470338 514170 470406 514226
rect 470462 514170 470558 514226
rect 469938 514102 470558 514170
rect 469938 514046 470034 514102
rect 470090 514046 470158 514102
rect 470214 514046 470282 514102
rect 470338 514046 470406 514102
rect 470462 514046 470558 514102
rect 469938 513978 470558 514046
rect 469938 513922 470034 513978
rect 470090 513922 470158 513978
rect 470214 513922 470282 513978
rect 470338 513922 470406 513978
rect 470462 513922 470558 513978
rect 469938 496350 470558 513922
rect 472892 553252 472948 553262
rect 472892 501508 472948 553196
rect 473228 552580 473284 552590
rect 473116 550564 473172 550574
rect 473004 546532 473060 546542
rect 473004 504980 473060 546476
rect 473116 510020 473172 550508
rect 473228 548548 473284 552524
rect 473228 548482 473284 548492
rect 473228 547876 473284 547886
rect 473228 513380 473284 547820
rect 473340 545860 473396 545870
rect 473340 523348 473396 545804
rect 473452 536788 473508 553868
rect 519036 553924 519092 554462
rect 519036 553858 519092 553868
rect 521276 551908 521332 551918
rect 495808 550350 496128 550384
rect 495808 550294 495878 550350
rect 495934 550294 496002 550350
rect 496058 550294 496128 550350
rect 495808 550226 496128 550294
rect 495808 550170 495878 550226
rect 495934 550170 496002 550226
rect 496058 550170 496128 550226
rect 495808 550102 496128 550170
rect 495808 550046 495878 550102
rect 495934 550046 496002 550102
rect 496058 550046 496128 550102
rect 495808 549978 496128 550046
rect 495808 549922 495878 549978
rect 495934 549922 496002 549978
rect 496058 549922 496128 549978
rect 495808 549888 496128 549922
rect 480448 544350 480768 544384
rect 480448 544294 480518 544350
rect 480574 544294 480642 544350
rect 480698 544294 480768 544350
rect 480448 544226 480768 544294
rect 480448 544170 480518 544226
rect 480574 544170 480642 544226
rect 480698 544170 480768 544226
rect 480448 544102 480768 544170
rect 480448 544046 480518 544102
rect 480574 544046 480642 544102
rect 480698 544046 480768 544102
rect 480448 543978 480768 544046
rect 480448 543922 480518 543978
rect 480574 543922 480642 543978
rect 480698 543922 480768 543978
rect 480448 543888 480768 543922
rect 496938 544350 497558 551602
rect 496938 544294 497034 544350
rect 497090 544294 497158 544350
rect 497214 544294 497282 544350
rect 497338 544294 497406 544350
rect 497462 544294 497558 544350
rect 496938 544226 497558 544294
rect 496938 544170 497034 544226
rect 497090 544170 497158 544226
rect 497214 544170 497282 544226
rect 497338 544170 497406 544226
rect 497462 544170 497558 544226
rect 496938 544102 497558 544170
rect 496938 544046 497034 544102
rect 497090 544046 497158 544102
rect 497214 544046 497282 544102
rect 497338 544046 497406 544102
rect 497462 544046 497558 544102
rect 496938 543978 497558 544046
rect 496938 543922 497034 543978
rect 497090 543922 497158 543978
rect 497214 543922 497282 543978
rect 497338 543922 497406 543978
rect 497462 543922 497558 543978
rect 473452 536722 473508 536732
rect 495808 532350 496128 532384
rect 495808 532294 495878 532350
rect 495934 532294 496002 532350
rect 496058 532294 496128 532350
rect 495808 532226 496128 532294
rect 495808 532170 495878 532226
rect 495934 532170 496002 532226
rect 496058 532170 496128 532226
rect 495808 532102 496128 532170
rect 495808 532046 495878 532102
rect 495934 532046 496002 532102
rect 496058 532046 496128 532102
rect 495808 531978 496128 532046
rect 495808 531922 495878 531978
rect 495934 531922 496002 531978
rect 496058 531922 496128 531978
rect 495808 531888 496128 531922
rect 473340 523282 473396 523292
rect 496938 526350 497558 543922
rect 496938 526294 497034 526350
rect 497090 526294 497158 526350
rect 497214 526294 497282 526350
rect 497338 526294 497406 526350
rect 497462 526294 497558 526350
rect 496938 526226 497558 526294
rect 496938 526170 497034 526226
rect 497090 526170 497158 526226
rect 497214 526170 497282 526226
rect 497338 526170 497406 526226
rect 497462 526170 497558 526226
rect 496938 526102 497558 526170
rect 496938 526046 497034 526102
rect 497090 526046 497158 526102
rect 497214 526046 497282 526102
rect 497338 526046 497406 526102
rect 497462 526046 497558 526102
rect 496938 525978 497558 526046
rect 496938 525922 497034 525978
rect 497090 525922 497158 525978
rect 497214 525922 497282 525978
rect 497338 525922 497406 525978
rect 497462 525922 497558 525978
rect 473228 513314 473284 513324
rect 473116 509954 473172 509964
rect 473004 504914 473060 504924
rect 496938 508350 497558 525922
rect 496938 508294 497034 508350
rect 497090 508294 497158 508350
rect 497214 508294 497282 508350
rect 497338 508294 497406 508350
rect 497462 508294 497558 508350
rect 496938 508226 497558 508294
rect 496938 508170 497034 508226
rect 497090 508170 497158 508226
rect 497214 508170 497282 508226
rect 497338 508170 497406 508226
rect 497462 508170 497558 508226
rect 496938 508102 497558 508170
rect 496938 508046 497034 508102
rect 497090 508046 497158 508102
rect 497214 508046 497282 508102
rect 497338 508046 497406 508102
rect 497462 508046 497558 508102
rect 496938 507978 497558 508046
rect 496938 507922 497034 507978
rect 497090 507922 497158 507978
rect 497214 507922 497282 507978
rect 497338 507922 497406 507978
rect 497462 507922 497558 507978
rect 472892 501442 472948 501452
rect 469938 496294 470034 496350
rect 470090 496294 470158 496350
rect 470214 496294 470282 496350
rect 470338 496294 470406 496350
rect 470462 496294 470558 496350
rect 469938 496226 470558 496294
rect 469938 496170 470034 496226
rect 470090 496170 470158 496226
rect 470214 496170 470282 496226
rect 470338 496170 470406 496226
rect 470462 496170 470558 496226
rect 469938 496102 470558 496170
rect 469938 496046 470034 496102
rect 470090 496046 470158 496102
rect 470214 496046 470282 496102
rect 470338 496046 470406 496102
rect 470462 496046 470558 496102
rect 469938 495978 470558 496046
rect 469938 495922 470034 495978
rect 470090 495922 470158 495978
rect 470214 495922 470282 495978
rect 470338 495922 470406 495978
rect 470462 495922 470558 495978
rect 469938 478350 470558 495922
rect 480448 490350 480768 490384
rect 480448 490294 480518 490350
rect 480574 490294 480642 490350
rect 480698 490294 480768 490350
rect 480448 490226 480768 490294
rect 480448 490170 480518 490226
rect 480574 490170 480642 490226
rect 480698 490170 480768 490226
rect 480448 490102 480768 490170
rect 480448 490046 480518 490102
rect 480574 490046 480642 490102
rect 480698 490046 480768 490102
rect 480448 489978 480768 490046
rect 480448 489922 480518 489978
rect 480574 489922 480642 489978
rect 480698 489922 480768 489978
rect 480448 489888 480768 489922
rect 496938 490350 497558 507922
rect 496938 490294 497034 490350
rect 497090 490294 497158 490350
rect 497214 490294 497282 490350
rect 497338 490294 497406 490350
rect 497462 490294 497558 490350
rect 496938 490226 497558 490294
rect 496938 490170 497034 490226
rect 497090 490170 497158 490226
rect 497214 490170 497282 490226
rect 497338 490170 497406 490226
rect 497462 490170 497558 490226
rect 496938 490102 497558 490170
rect 496938 490046 497034 490102
rect 497090 490046 497158 490102
rect 497214 490046 497282 490102
rect 497338 490046 497406 490102
rect 497462 490046 497558 490102
rect 496938 489978 497558 490046
rect 496938 489922 497034 489978
rect 497090 489922 497158 489978
rect 497214 489922 497282 489978
rect 497338 489922 497406 489978
rect 497462 489922 497558 489978
rect 476028 484678 476084 484688
rect 476028 484372 476084 484622
rect 476028 484306 476084 484316
rect 473676 484036 473732 484046
rect 473676 483958 473732 483980
rect 473676 483892 473732 483902
rect 472108 482692 472164 482702
rect 472108 481460 472164 482636
rect 472108 481394 472164 481404
rect 472220 482020 472276 482030
rect 472220 480538 472276 481964
rect 472220 480472 472276 480482
rect 469938 478294 470034 478350
rect 470090 478294 470158 478350
rect 470214 478294 470282 478350
rect 470338 478294 470406 478350
rect 470462 478294 470558 478350
rect 469938 478226 470558 478294
rect 469938 478170 470034 478226
rect 470090 478170 470158 478226
rect 470214 478170 470282 478226
rect 470338 478170 470406 478226
rect 470462 478170 470558 478226
rect 469938 478102 470558 478170
rect 469938 478046 470034 478102
rect 470090 478046 470158 478102
rect 470214 478046 470282 478102
rect 470338 478046 470406 478102
rect 470462 478046 470558 478102
rect 466218 472294 466314 472350
rect 466370 472294 466438 472350
rect 466494 472294 466562 472350
rect 466618 472294 466686 472350
rect 466742 472294 466838 472350
rect 466218 472226 466838 472294
rect 466218 472170 466314 472226
rect 466370 472170 466438 472226
rect 466494 472170 466562 472226
rect 466618 472170 466686 472226
rect 466742 472170 466838 472226
rect 466218 472102 466838 472170
rect 466218 472046 466314 472102
rect 466370 472046 466438 472102
rect 466494 472046 466562 472102
rect 466618 472046 466686 472102
rect 466742 472046 466838 472102
rect 466218 471978 466838 472046
rect 466218 471922 466314 471978
rect 466370 471922 466438 471978
rect 466494 471922 466562 471978
rect 466618 471922 466686 471978
rect 466742 471922 466838 471978
rect 461132 430770 461188 430780
rect 466218 454350 466838 471922
rect 466218 454294 466314 454350
rect 466370 454294 466438 454350
rect 466494 454294 466562 454350
rect 466618 454294 466686 454350
rect 466742 454294 466838 454350
rect 466218 454226 466838 454294
rect 466218 454170 466314 454226
rect 466370 454170 466438 454226
rect 466494 454170 466562 454226
rect 466618 454170 466686 454226
rect 466742 454170 466838 454226
rect 466218 454102 466838 454170
rect 466218 454046 466314 454102
rect 466370 454046 466438 454102
rect 466494 454046 466562 454102
rect 466618 454046 466686 454102
rect 466742 454046 466838 454102
rect 466218 453978 466838 454046
rect 466218 453922 466314 453978
rect 466370 453922 466438 453978
rect 466494 453922 466562 453978
rect 466618 453922 466686 453978
rect 466742 453922 466838 453978
rect 466218 436350 466838 453922
rect 466218 436294 466314 436350
rect 466370 436294 466438 436350
rect 466494 436294 466562 436350
rect 466618 436294 466686 436350
rect 466742 436294 466838 436350
rect 466218 436226 466838 436294
rect 466218 436170 466314 436226
rect 466370 436170 466438 436226
rect 466494 436170 466562 436226
rect 466618 436170 466686 436226
rect 466742 436170 466838 436226
rect 466218 436102 466838 436170
rect 466218 436046 466314 436102
rect 466370 436046 466438 436102
rect 466494 436046 466562 436102
rect 466618 436046 466686 436102
rect 466742 436046 466838 436102
rect 466218 435978 466838 436046
rect 466218 435922 466314 435978
rect 466370 435922 466438 435978
rect 466494 435922 466562 435978
rect 466618 435922 466686 435978
rect 466742 435922 466838 435978
rect 457100 427410 457156 427420
rect 456988 424610 457044 424620
rect 439218 424294 439314 424350
rect 439370 424294 439438 424350
rect 439494 424294 439562 424350
rect 439618 424294 439686 424350
rect 439742 424294 439838 424350
rect 439218 424226 439838 424294
rect 439218 424170 439314 424226
rect 439370 424170 439438 424226
rect 439494 424170 439562 424226
rect 439618 424170 439686 424226
rect 439742 424170 439838 424226
rect 439218 424102 439838 424170
rect 439218 424046 439314 424102
rect 439370 424046 439438 424102
rect 439494 424046 439562 424102
rect 439618 424046 439686 424102
rect 439742 424046 439838 424102
rect 439218 423978 439838 424046
rect 439218 423922 439314 423978
rect 439370 423922 439438 423978
rect 439494 423922 439562 423978
rect 439618 423922 439686 423978
rect 439742 423922 439838 423978
rect 439218 409918 439838 423922
rect 449168 418350 449488 418384
rect 449168 418294 449238 418350
rect 449294 418294 449362 418350
rect 449418 418294 449488 418350
rect 449168 418226 449488 418294
rect 449168 418170 449238 418226
rect 449294 418170 449362 418226
rect 449418 418170 449488 418226
rect 449168 418102 449488 418170
rect 449168 418046 449238 418102
rect 449294 418046 449362 418102
rect 449418 418046 449488 418102
rect 449168 417978 449488 418046
rect 449168 417922 449238 417978
rect 449294 417922 449362 417978
rect 449418 417922 449488 417978
rect 449168 417888 449488 417922
rect 466218 418350 466838 435922
rect 467852 477988 467908 477998
rect 467852 431956 467908 477932
rect 467852 431890 467908 431900
rect 469938 477978 470558 478046
rect 469938 477922 470034 477978
rect 470090 477922 470158 477978
rect 470214 477922 470282 477978
rect 470338 477922 470406 477978
rect 470462 477922 470558 477978
rect 469938 460350 470558 477922
rect 469938 460294 470034 460350
rect 470090 460294 470158 460350
rect 470214 460294 470282 460350
rect 470338 460294 470406 460350
rect 470462 460294 470558 460350
rect 469938 460226 470558 460294
rect 469938 460170 470034 460226
rect 470090 460170 470158 460226
rect 470214 460170 470282 460226
rect 470338 460170 470406 460226
rect 470462 460170 470558 460226
rect 469938 460102 470558 460170
rect 469938 460046 470034 460102
rect 470090 460046 470158 460102
rect 470214 460046 470282 460102
rect 470338 460046 470406 460102
rect 470462 460046 470558 460102
rect 469938 459978 470558 460046
rect 469938 459922 470034 459978
rect 470090 459922 470158 459978
rect 470214 459922 470282 459978
rect 470338 459922 470406 459978
rect 470462 459922 470558 459978
rect 469938 442350 470558 459922
rect 472892 480004 472948 480014
rect 472892 444612 472948 479948
rect 473116 479332 473172 479342
rect 473116 465238 473172 479276
rect 495808 478350 496128 478384
rect 495808 478294 495878 478350
rect 495934 478294 496002 478350
rect 496058 478294 496128 478350
rect 495808 478226 496128 478294
rect 495808 478170 495878 478226
rect 495934 478170 496002 478226
rect 496058 478170 496128 478226
rect 495808 478102 496128 478170
rect 495808 478046 495878 478102
rect 495934 478046 496002 478102
rect 496058 478046 496128 478102
rect 495808 477978 496128 478046
rect 495808 477922 495878 477978
rect 495934 477922 496002 477978
rect 496058 477922 496128 477978
rect 495808 477888 496128 477922
rect 496938 476414 497558 489922
rect 500658 550350 501278 551602
rect 500658 550294 500754 550350
rect 500810 550294 500878 550350
rect 500934 550294 501002 550350
rect 501058 550294 501126 550350
rect 501182 550294 501278 550350
rect 500658 550226 501278 550294
rect 500658 550170 500754 550226
rect 500810 550170 500878 550226
rect 500934 550170 501002 550226
rect 501058 550170 501126 550226
rect 501182 550170 501278 550226
rect 500658 550102 501278 550170
rect 500658 550046 500754 550102
rect 500810 550046 500878 550102
rect 500934 550046 501002 550102
rect 501058 550046 501126 550102
rect 501182 550046 501278 550102
rect 500658 549978 501278 550046
rect 500658 549922 500754 549978
rect 500810 549922 500878 549978
rect 500934 549922 501002 549978
rect 501058 549922 501126 549978
rect 501182 549922 501278 549978
rect 500658 532350 501278 549922
rect 518252 551124 518308 551134
rect 511168 544350 511488 544384
rect 511168 544294 511238 544350
rect 511294 544294 511362 544350
rect 511418 544294 511488 544350
rect 511168 544226 511488 544294
rect 511168 544170 511238 544226
rect 511294 544170 511362 544226
rect 511418 544170 511488 544226
rect 511168 544102 511488 544170
rect 511168 544046 511238 544102
rect 511294 544046 511362 544102
rect 511418 544046 511488 544102
rect 511168 543978 511488 544046
rect 511168 543922 511238 543978
rect 511294 543922 511362 543978
rect 511418 543922 511488 543978
rect 511168 543888 511488 543922
rect 500658 532294 500754 532350
rect 500810 532294 500878 532350
rect 500934 532294 501002 532350
rect 501058 532294 501126 532350
rect 501182 532294 501278 532350
rect 500658 532226 501278 532294
rect 500658 532170 500754 532226
rect 500810 532170 500878 532226
rect 500934 532170 501002 532226
rect 501058 532170 501126 532226
rect 501182 532170 501278 532226
rect 500658 532102 501278 532170
rect 500658 532046 500754 532102
rect 500810 532046 500878 532102
rect 500934 532046 501002 532102
rect 501058 532046 501126 532102
rect 501182 532046 501278 532102
rect 500658 531978 501278 532046
rect 500658 531922 500754 531978
rect 500810 531922 500878 531978
rect 500934 531922 501002 531978
rect 501058 531922 501126 531978
rect 501182 531922 501278 531978
rect 500658 514350 501278 531922
rect 518252 522676 518308 551068
rect 520940 549892 520996 549902
rect 519260 546532 519316 546542
rect 519148 544516 519204 544526
rect 519036 533428 519092 533438
rect 519036 528276 519092 533372
rect 519036 528210 519092 528220
rect 518252 522610 518308 522620
rect 519148 516628 519204 544460
rect 519260 519316 519316 546476
rect 519260 519250 519316 519260
rect 519932 544852 519988 544862
rect 519932 518196 519988 544796
rect 520828 543172 520884 543182
rect 520828 527940 520884 543116
rect 520828 527874 520884 527884
rect 519932 518130 519988 518140
rect 519148 516562 519204 516572
rect 500658 514294 500754 514350
rect 500810 514294 500878 514350
rect 500934 514294 501002 514350
rect 501058 514294 501126 514350
rect 501182 514294 501278 514350
rect 500658 514226 501278 514294
rect 500658 514170 500754 514226
rect 500810 514170 500878 514226
rect 500934 514170 501002 514226
rect 501058 514170 501126 514226
rect 501182 514170 501278 514226
rect 500658 514102 501278 514170
rect 500658 514046 500754 514102
rect 500810 514046 500878 514102
rect 500934 514046 501002 514102
rect 501058 514046 501126 514102
rect 501182 514046 501278 514102
rect 500658 513978 501278 514046
rect 500658 513922 500754 513978
rect 500810 513922 500878 513978
rect 500934 513922 501002 513978
rect 501058 513922 501126 513978
rect 501182 513922 501278 513978
rect 500658 496350 501278 513922
rect 520940 511588 520996 549836
rect 521052 547204 521108 547214
rect 521052 519988 521108 547148
rect 521164 541828 521220 541838
rect 521164 523796 521220 541772
rect 521164 523730 521220 523740
rect 521052 519922 521108 519932
rect 520940 511522 520996 511532
rect 521276 506548 521332 551852
rect 523292 548548 523348 548558
rect 523292 530516 523348 548492
rect 523292 530450 523348 530460
rect 527658 544350 528278 561922
rect 527658 544294 527754 544350
rect 527810 544294 527878 544350
rect 527934 544294 528002 544350
rect 528058 544294 528126 544350
rect 528182 544294 528278 544350
rect 527658 544226 528278 544294
rect 527658 544170 527754 544226
rect 527810 544170 527878 544226
rect 527934 544170 528002 544226
rect 528058 544170 528126 544226
rect 528182 544170 528278 544226
rect 527658 544102 528278 544170
rect 527658 544046 527754 544102
rect 527810 544046 527878 544102
rect 527934 544046 528002 544102
rect 528058 544046 528126 544102
rect 528182 544046 528278 544102
rect 527658 543978 528278 544046
rect 527658 543922 527754 543978
rect 527810 543922 527878 543978
rect 527934 543922 528002 543978
rect 528058 543922 528126 543978
rect 528182 543922 528278 543978
rect 521276 506482 521332 506492
rect 527658 526350 528278 543922
rect 527658 526294 527754 526350
rect 527810 526294 527878 526350
rect 527934 526294 528002 526350
rect 528058 526294 528126 526350
rect 528182 526294 528278 526350
rect 527658 526226 528278 526294
rect 527658 526170 527754 526226
rect 527810 526170 527878 526226
rect 527934 526170 528002 526226
rect 528058 526170 528126 526226
rect 528182 526170 528278 526226
rect 527658 526102 528278 526170
rect 527658 526046 527754 526102
rect 527810 526046 527878 526102
rect 527934 526046 528002 526102
rect 528058 526046 528126 526102
rect 528182 526046 528278 526102
rect 527658 525978 528278 526046
rect 527658 525922 527754 525978
rect 527810 525922 527878 525978
rect 527934 525922 528002 525978
rect 528058 525922 528126 525978
rect 528182 525922 528278 525978
rect 527658 508350 528278 525922
rect 527658 508294 527754 508350
rect 527810 508294 527878 508350
rect 527934 508294 528002 508350
rect 528058 508294 528126 508350
rect 528182 508294 528278 508350
rect 527658 508226 528278 508294
rect 527658 508170 527754 508226
rect 527810 508170 527878 508226
rect 527934 508170 528002 508226
rect 528058 508170 528126 508226
rect 528182 508170 528278 508226
rect 527658 508102 528278 508170
rect 527658 508046 527754 508102
rect 527810 508046 527878 508102
rect 527934 508046 528002 508102
rect 528058 508046 528126 508102
rect 528182 508046 528278 508102
rect 527658 507978 528278 508046
rect 527658 507922 527754 507978
rect 527810 507922 527878 507978
rect 527934 507922 528002 507978
rect 528058 507922 528126 507978
rect 528182 507922 528278 507978
rect 500658 496294 500754 496350
rect 500810 496294 500878 496350
rect 500934 496294 501002 496350
rect 501058 496294 501126 496350
rect 501182 496294 501278 496350
rect 500658 496226 501278 496294
rect 500658 496170 500754 496226
rect 500810 496170 500878 496226
rect 500934 496170 501002 496226
rect 501058 496170 501126 496226
rect 501182 496170 501278 496226
rect 500658 496102 501278 496170
rect 500658 496046 500754 496102
rect 500810 496046 500878 496102
rect 500934 496046 501002 496102
rect 501058 496046 501126 496102
rect 501182 496046 501278 496102
rect 500658 495978 501278 496046
rect 500658 495922 500754 495978
rect 500810 495922 500878 495978
rect 500934 495922 501002 495978
rect 501058 495922 501126 495978
rect 501182 495922 501278 495978
rect 500658 478350 501278 495922
rect 511168 490350 511488 490384
rect 511168 490294 511238 490350
rect 511294 490294 511362 490350
rect 511418 490294 511488 490350
rect 511168 490226 511488 490294
rect 511168 490170 511238 490226
rect 511294 490170 511362 490226
rect 511418 490170 511488 490226
rect 511168 490102 511488 490170
rect 511168 490046 511238 490102
rect 511294 490046 511362 490102
rect 511418 490046 511488 490102
rect 511168 489978 511488 490046
rect 511168 489922 511238 489978
rect 511294 489922 511362 489978
rect 511418 489922 511488 489978
rect 511168 489888 511488 489922
rect 527658 490350 528278 507922
rect 527658 490294 527754 490350
rect 527810 490294 527878 490350
rect 527934 490294 528002 490350
rect 528058 490294 528126 490350
rect 528182 490294 528278 490350
rect 527658 490226 528278 490294
rect 527658 490170 527754 490226
rect 527810 490170 527878 490226
rect 527934 490170 528002 490226
rect 528058 490170 528126 490226
rect 528182 490170 528278 490226
rect 527658 490102 528278 490170
rect 527658 490046 527754 490102
rect 527810 490046 527878 490102
rect 527934 490046 528002 490102
rect 528058 490046 528126 490102
rect 528182 490046 528278 490102
rect 527658 489978 528278 490046
rect 527658 489922 527754 489978
rect 527810 489922 527878 489978
rect 527934 489922 528002 489978
rect 528058 489922 528126 489978
rect 528182 489922 528278 489978
rect 519148 483364 519204 483374
rect 518252 481908 518308 481918
rect 500658 478294 500754 478350
rect 500810 478294 500878 478350
rect 500934 478294 501002 478350
rect 501058 478294 501126 478350
rect 501182 478294 501278 478350
rect 500658 478226 501278 478294
rect 500658 478170 500754 478226
rect 500810 478170 500878 478226
rect 500934 478170 501002 478226
rect 501058 478170 501126 478226
rect 501182 478170 501278 478226
rect 500658 478102 501278 478170
rect 500658 478046 500754 478102
rect 500810 478046 500878 478102
rect 500934 478046 501002 478102
rect 501058 478046 501126 478102
rect 501182 478046 501278 478102
rect 500658 477978 501278 478046
rect 500658 477922 500754 477978
rect 500810 477922 500878 477978
rect 500934 477922 501002 477978
rect 501058 477922 501126 477978
rect 501182 477922 501278 477978
rect 480448 472350 480768 472384
rect 480448 472294 480518 472350
rect 480574 472294 480642 472350
rect 480698 472294 480768 472350
rect 480448 472226 480768 472294
rect 480448 472170 480518 472226
rect 480574 472170 480642 472226
rect 480698 472170 480768 472226
rect 480448 472102 480768 472170
rect 480448 472046 480518 472102
rect 480574 472046 480642 472102
rect 480698 472046 480768 472102
rect 480448 471978 480768 472046
rect 480448 471922 480518 471978
rect 480574 471922 480642 471978
rect 480698 471922 480768 471978
rect 480448 471888 480768 471922
rect 473116 465172 473172 465182
rect 495808 460350 496128 460384
rect 495808 460294 495878 460350
rect 495934 460294 496002 460350
rect 496058 460294 496128 460350
rect 495808 460226 496128 460294
rect 495808 460170 495878 460226
rect 495934 460170 496002 460226
rect 496058 460170 496128 460226
rect 495808 460102 496128 460170
rect 495808 460046 495878 460102
rect 495934 460046 496002 460102
rect 496058 460046 496128 460102
rect 495808 459978 496128 460046
rect 495808 459922 495878 459978
rect 495934 459922 496002 459978
rect 496058 459922 496128 459978
rect 495808 459888 496128 459922
rect 493724 457940 493780 457950
rect 493724 457156 493780 457884
rect 493724 457090 493780 457100
rect 472892 444546 472948 444556
rect 496938 454350 497558 470322
rect 496938 454294 497034 454350
rect 497090 454294 497158 454350
rect 497214 454294 497282 454350
rect 497338 454294 497406 454350
rect 497462 454294 497558 454350
rect 496938 454226 497558 454294
rect 496938 454170 497034 454226
rect 497090 454170 497158 454226
rect 497214 454170 497282 454226
rect 497338 454170 497406 454226
rect 497462 454170 497558 454226
rect 496938 454102 497558 454170
rect 496938 454046 497034 454102
rect 497090 454046 497158 454102
rect 497214 454046 497282 454102
rect 497338 454046 497406 454102
rect 497462 454046 497558 454102
rect 496938 453978 497558 454046
rect 496938 453922 497034 453978
rect 497090 453922 497158 453978
rect 497214 453922 497282 453978
rect 497338 453922 497406 453978
rect 497462 453922 497558 453978
rect 469938 442294 470034 442350
rect 470090 442294 470158 442350
rect 470214 442294 470282 442350
rect 470338 442294 470406 442350
rect 470462 442294 470558 442350
rect 469938 442226 470558 442294
rect 469938 442170 470034 442226
rect 470090 442170 470158 442226
rect 470214 442170 470282 442226
rect 470338 442170 470406 442226
rect 470462 442170 470558 442226
rect 469938 442102 470558 442170
rect 469938 442046 470034 442102
rect 470090 442046 470158 442102
rect 470214 442046 470282 442102
rect 470338 442046 470406 442102
rect 470462 442046 470558 442102
rect 469938 441978 470558 442046
rect 469938 441922 470034 441978
rect 470090 441922 470158 441978
rect 470214 441922 470282 441978
rect 470338 441922 470406 441978
rect 470462 441922 470558 441978
rect 466218 418294 466314 418350
rect 466370 418294 466438 418350
rect 466494 418294 466562 418350
rect 466618 418294 466686 418350
rect 466742 418294 466838 418350
rect 466218 418226 466838 418294
rect 466218 418170 466314 418226
rect 466370 418170 466438 418226
rect 466494 418170 466562 418226
rect 466618 418170 466686 418226
rect 466742 418170 466838 418226
rect 466218 418102 466838 418170
rect 466218 418046 466314 418102
rect 466370 418046 466438 418102
rect 466494 418046 466562 418102
rect 466618 418046 466686 418102
rect 466742 418046 466838 418102
rect 466218 417978 466838 418046
rect 466218 417922 466314 417978
rect 466370 417922 466438 417978
rect 466494 417922 466562 417978
rect 466618 417922 466686 417978
rect 466742 417922 466838 417978
rect 440972 411958 441028 411968
rect 428876 407392 428932 407402
rect 440972 407458 441028 411902
rect 464492 411460 464548 411470
rect 457324 410788 457380 410798
rect 456092 409444 456148 409454
rect 440972 407392 441028 407402
rect 455532 407428 455588 407438
rect 433808 406350 434128 406384
rect 433808 406294 433878 406350
rect 433934 406294 434002 406350
rect 434058 406294 434128 406350
rect 433808 406226 434128 406294
rect 433808 406170 433878 406226
rect 433934 406170 434002 406226
rect 434058 406170 434128 406226
rect 433808 406102 434128 406170
rect 433808 406046 433878 406102
rect 433934 406046 434002 406102
rect 434058 406046 434128 406102
rect 433808 405978 434128 406046
rect 433808 405922 433878 405978
rect 433934 405922 434002 405978
rect 434058 405922 434128 405978
rect 433808 405888 434128 405922
rect 414092 402892 414148 402902
rect 411180 402322 411236 402332
rect 411180 402052 411236 402062
rect 411180 398098 411236 401996
rect 418448 400350 418768 400384
rect 418448 400294 418518 400350
rect 418574 400294 418642 400350
rect 418698 400294 418768 400350
rect 418448 400226 418768 400294
rect 418448 400170 418518 400226
rect 418574 400170 418642 400226
rect 418698 400170 418768 400226
rect 418448 400102 418768 400170
rect 418448 400046 418518 400102
rect 418574 400046 418642 400102
rect 418698 400046 418768 400102
rect 418448 399978 418768 400046
rect 418448 399922 418518 399978
rect 418574 399922 418642 399978
rect 418698 399922 418768 399978
rect 418448 399888 418768 399922
rect 435498 400350 436118 404498
rect 435498 400294 435594 400350
rect 435650 400294 435718 400350
rect 435774 400294 435842 400350
rect 435898 400294 435966 400350
rect 436022 400294 436118 400350
rect 435498 400226 436118 400294
rect 435498 400170 435594 400226
rect 435650 400170 435718 400226
rect 435774 400170 435842 400226
rect 435898 400170 435966 400226
rect 436022 400170 436118 400226
rect 435498 400102 436118 400170
rect 435498 400046 435594 400102
rect 435650 400046 435718 400102
rect 435774 400046 435842 400102
rect 435898 400046 435966 400102
rect 436022 400046 436118 400102
rect 435498 399978 436118 400046
rect 435498 399922 435594 399978
rect 435650 399922 435718 399978
rect 435774 399922 435842 399978
rect 435898 399922 435966 399978
rect 436022 399922 436118 399978
rect 411180 398032 411236 398042
rect 410732 394432 410788 394442
rect 408498 388294 408594 388350
rect 408650 388294 408718 388350
rect 408774 388294 408842 388350
rect 408898 388294 408966 388350
rect 409022 388294 409118 388350
rect 408498 388226 409118 388294
rect 433808 388389 434128 388446
rect 433808 388333 433836 388389
rect 433892 388333 433940 388389
rect 433996 388333 434044 388389
rect 434100 388333 434128 388389
rect 433808 388276 434128 388333
rect 408498 388170 408594 388226
rect 408650 388170 408718 388226
rect 408774 388170 408842 388226
rect 408898 388170 408966 388226
rect 409022 388170 409118 388226
rect 408498 388102 409118 388170
rect 408498 388046 408594 388102
rect 408650 388046 408718 388102
rect 408774 388046 408842 388102
rect 408898 388046 408966 388102
rect 409022 388046 409118 388102
rect 408498 387978 409118 388046
rect 408498 387922 408594 387978
rect 408650 387922 408718 387978
rect 408774 387922 408842 387978
rect 408898 387922 408966 387978
rect 409022 387922 409118 387978
rect 408498 370350 409118 387922
rect 408498 370294 408594 370350
rect 408650 370294 408718 370350
rect 408774 370294 408842 370350
rect 408898 370294 408966 370350
rect 409022 370294 409118 370350
rect 408498 370226 409118 370294
rect 408498 370170 408594 370226
rect 408650 370170 408718 370226
rect 408774 370170 408842 370226
rect 408898 370170 408966 370226
rect 409022 370170 409118 370226
rect 408498 370102 409118 370170
rect 408498 370046 408594 370102
rect 408650 370046 408718 370102
rect 408774 370046 408842 370102
rect 408898 370046 408966 370102
rect 409022 370046 409118 370102
rect 408498 369978 409118 370046
rect 408498 369922 408594 369978
rect 408650 369922 408718 369978
rect 408774 369922 408842 369978
rect 408898 369922 408966 369978
rect 409022 369922 409118 369978
rect 408498 352350 409118 369922
rect 435498 382350 436118 399922
rect 435498 382294 435594 382350
rect 435650 382294 435718 382350
rect 435774 382294 435842 382350
rect 435898 382294 435966 382350
rect 436022 382294 436118 382350
rect 435498 382226 436118 382294
rect 435498 382170 435594 382226
rect 435650 382170 435718 382226
rect 435774 382170 435842 382226
rect 435898 382170 435966 382226
rect 436022 382170 436118 382226
rect 435498 382102 436118 382170
rect 435498 382046 435594 382102
rect 435650 382046 435718 382102
rect 435774 382046 435842 382102
rect 435898 382046 435966 382102
rect 436022 382046 436118 382102
rect 435498 381978 436118 382046
rect 435498 381922 435594 381978
rect 435650 381922 435718 381978
rect 435774 381922 435842 381978
rect 435898 381922 435966 381978
rect 436022 381922 436118 381978
rect 435498 364350 436118 381922
rect 435498 364294 435594 364350
rect 435650 364294 435718 364350
rect 435774 364294 435842 364350
rect 435898 364294 435966 364350
rect 436022 364294 436118 364350
rect 435498 364226 436118 364294
rect 435498 364170 435594 364226
rect 435650 364170 435718 364226
rect 435774 364170 435842 364226
rect 435898 364170 435966 364226
rect 436022 364170 436118 364226
rect 435498 364102 436118 364170
rect 435498 364046 435594 364102
rect 435650 364046 435718 364102
rect 435774 364046 435842 364102
rect 435898 364046 435966 364102
rect 436022 364046 436118 364102
rect 435498 363978 436118 364046
rect 435498 363922 435594 363978
rect 435650 363922 435718 363978
rect 435774 363922 435842 363978
rect 435898 363922 435966 363978
rect 436022 363922 436118 363978
rect 408498 352294 408594 352350
rect 408650 352294 408718 352350
rect 408774 352294 408842 352350
rect 408898 352294 408966 352350
rect 409022 352294 409118 352350
rect 408498 352226 409118 352294
rect 408498 352170 408594 352226
rect 408650 352170 408718 352226
rect 408774 352170 408842 352226
rect 408898 352170 408966 352226
rect 409022 352170 409118 352226
rect 408498 352102 409118 352170
rect 408498 352046 408594 352102
rect 408650 352046 408718 352102
rect 408774 352046 408842 352102
rect 408898 352046 408966 352102
rect 409022 352046 409118 352102
rect 408498 351978 409118 352046
rect 408498 351922 408594 351978
rect 408650 351922 408718 351978
rect 408774 351922 408842 351978
rect 408898 351922 408966 351978
rect 409022 351922 409118 351978
rect 407372 341578 407428 341588
rect 407372 330260 407428 341522
rect 407372 330194 407428 330204
rect 408498 334350 409118 351922
rect 433808 352350 434128 352384
rect 433808 352294 433878 352350
rect 433934 352294 434002 352350
rect 434058 352294 434128 352350
rect 433808 352226 434128 352294
rect 433808 352170 433878 352226
rect 433934 352170 434002 352226
rect 434058 352170 434128 352226
rect 433808 352102 434128 352170
rect 433808 352046 433878 352102
rect 433934 352046 434002 352102
rect 434058 352046 434128 352102
rect 433808 351978 434128 352046
rect 433808 351922 433878 351978
rect 433934 351922 434002 351978
rect 434058 351922 434128 351978
rect 433808 351888 434128 351922
rect 418448 346350 418768 346384
rect 418448 346294 418518 346350
rect 418574 346294 418642 346350
rect 418698 346294 418768 346350
rect 418448 346226 418768 346294
rect 418448 346170 418518 346226
rect 418574 346170 418642 346226
rect 418698 346170 418768 346226
rect 418448 346102 418768 346170
rect 418448 346046 418518 346102
rect 418574 346046 418642 346102
rect 418698 346046 418768 346102
rect 418448 345978 418768 346046
rect 418448 345922 418518 345978
rect 418574 345922 418642 345978
rect 418698 345922 418768 345978
rect 418448 345888 418768 345922
rect 435498 346350 436118 363922
rect 435498 346294 435594 346350
rect 435650 346294 435718 346350
rect 435774 346294 435842 346350
rect 435898 346294 435966 346350
rect 436022 346294 436118 346350
rect 435498 346226 436118 346294
rect 435498 346170 435594 346226
rect 435650 346170 435718 346226
rect 435774 346170 435842 346226
rect 435898 346170 435966 346226
rect 436022 346170 436118 346226
rect 435498 346102 436118 346170
rect 435498 346046 435594 346102
rect 435650 346046 435718 346102
rect 435774 346046 435842 346102
rect 435898 346046 435966 346102
rect 436022 346046 436118 346102
rect 435498 345978 436118 346046
rect 435498 345922 435594 345978
rect 435650 345922 435718 345978
rect 435774 345922 435842 345978
rect 435898 345922 435966 345978
rect 436022 345922 436118 345978
rect 414652 341218 414708 341228
rect 414652 341012 414708 341162
rect 414652 340946 414708 340956
rect 408498 334294 408594 334350
rect 408650 334294 408718 334350
rect 408774 334294 408842 334350
rect 408898 334294 408966 334350
rect 409022 334294 409118 334350
rect 408498 334226 409118 334294
rect 408498 334170 408594 334226
rect 408650 334170 408718 334226
rect 408774 334170 408842 334226
rect 408898 334170 408966 334226
rect 409022 334170 409118 334226
rect 408498 334102 409118 334170
rect 408498 334046 408594 334102
rect 408650 334046 408718 334102
rect 408774 334046 408842 334102
rect 408898 334046 408966 334102
rect 409022 334046 409118 334102
rect 408498 333978 409118 334046
rect 408498 333922 408594 333978
rect 408650 333922 408718 333978
rect 408774 333922 408842 333978
rect 408898 333922 408966 333978
rect 409022 333922 409118 333978
rect 404778 328294 404874 328350
rect 404930 328294 404998 328350
rect 405054 328294 405122 328350
rect 405178 328294 405246 328350
rect 405302 328294 405398 328350
rect 404778 328226 405398 328294
rect 404778 328170 404874 328226
rect 404930 328170 404998 328226
rect 405054 328170 405122 328226
rect 405178 328170 405246 328226
rect 405302 328170 405398 328226
rect 404778 328102 405398 328170
rect 404778 328046 404874 328102
rect 404930 328046 404998 328102
rect 405054 328046 405122 328102
rect 405178 328046 405246 328102
rect 405302 328046 405398 328102
rect 404778 327978 405398 328046
rect 404778 327922 404874 327978
rect 404930 327922 404998 327978
rect 405054 327922 405122 327978
rect 405178 327922 405246 327978
rect 405302 327922 405398 327978
rect 404572 326818 404628 326828
rect 404572 320878 404628 326762
rect 404572 320812 404628 320822
rect 396844 302530 396900 302540
rect 404778 310350 405398 327922
rect 404778 310294 404874 310350
rect 404930 310294 404998 310350
rect 405054 310294 405122 310350
rect 405178 310294 405246 310350
rect 405302 310294 405398 310350
rect 404778 310226 405398 310294
rect 404778 310170 404874 310226
rect 404930 310170 404998 310226
rect 405054 310170 405122 310226
rect 405178 310170 405246 310226
rect 405302 310170 405398 310226
rect 404778 310102 405398 310170
rect 404778 310046 404874 310102
rect 404930 310046 404998 310102
rect 405054 310046 405122 310102
rect 405178 310046 405246 310102
rect 405302 310046 405398 310102
rect 404778 309978 405398 310046
rect 404778 309922 404874 309978
rect 404930 309922 404998 309978
rect 405054 309922 405122 309978
rect 405178 309922 405246 309978
rect 405302 309922 405398 309978
rect 395612 299170 395668 299180
rect 377778 298294 377874 298350
rect 377930 298294 377998 298350
rect 378054 298294 378122 298350
rect 378178 298294 378246 298350
rect 378302 298294 378398 298350
rect 377778 298226 378398 298294
rect 377778 298170 377874 298226
rect 377930 298170 377998 298226
rect 378054 298170 378122 298226
rect 378178 298170 378246 298226
rect 378302 298170 378398 298226
rect 377778 298102 378398 298170
rect 377778 298046 377874 298102
rect 377930 298046 377998 298102
rect 378054 298046 378122 298102
rect 378178 298046 378246 298102
rect 378302 298046 378398 298102
rect 377778 297978 378398 298046
rect 377778 297922 377874 297978
rect 377930 297922 377998 297978
rect 378054 297922 378122 297978
rect 378178 297922 378246 297978
rect 378302 297922 378398 297978
rect 377778 280350 378398 297922
rect 377778 280294 377874 280350
rect 377930 280294 377998 280350
rect 378054 280294 378122 280350
rect 378178 280294 378246 280350
rect 378302 280294 378398 280350
rect 377778 280226 378398 280294
rect 377778 280170 377874 280226
rect 377930 280170 377998 280226
rect 378054 280170 378122 280226
rect 378178 280170 378246 280226
rect 378302 280170 378398 280226
rect 377778 280102 378398 280170
rect 377778 280046 377874 280102
rect 377930 280046 377998 280102
rect 378054 280046 378122 280102
rect 378178 280046 378246 280102
rect 378302 280046 378398 280102
rect 377778 279978 378398 280046
rect 377778 279922 377874 279978
rect 377930 279922 377998 279978
rect 378054 279922 378122 279978
rect 378178 279922 378246 279978
rect 378302 279922 378398 279978
rect 377778 262350 378398 279922
rect 404778 292350 405398 309922
rect 404778 292294 404874 292350
rect 404930 292294 404998 292350
rect 405054 292294 405122 292350
rect 405178 292294 405246 292350
rect 405302 292294 405398 292350
rect 404778 292226 405398 292294
rect 404778 292170 404874 292226
rect 404930 292170 404998 292226
rect 405054 292170 405122 292226
rect 405178 292170 405246 292226
rect 405302 292170 405398 292226
rect 404778 292102 405398 292170
rect 404778 292046 404874 292102
rect 404930 292046 404998 292102
rect 405054 292046 405122 292102
rect 405178 292046 405246 292102
rect 405302 292046 405398 292102
rect 404778 291978 405398 292046
rect 404778 291922 404874 291978
rect 404930 291922 404998 291978
rect 405054 291922 405122 291978
rect 405178 291922 405246 291978
rect 405302 291922 405398 291978
rect 394828 275698 394884 275708
rect 387168 274350 387488 274384
rect 387168 274294 387238 274350
rect 387294 274294 387362 274350
rect 387418 274294 387488 274350
rect 387168 274226 387488 274294
rect 387168 274170 387238 274226
rect 387294 274170 387362 274226
rect 387418 274170 387488 274226
rect 387168 274102 387488 274170
rect 387168 274046 387238 274102
rect 387294 274046 387362 274102
rect 387418 274046 387488 274102
rect 387168 273978 387488 274046
rect 387168 273922 387238 273978
rect 387294 273922 387362 273978
rect 387418 273922 387488 273978
rect 387168 273888 387488 273922
rect 394828 271378 394884 275642
rect 404778 274350 405398 291922
rect 404778 274294 404874 274350
rect 404930 274294 404998 274350
rect 405054 274294 405122 274350
rect 405178 274294 405246 274350
rect 405302 274294 405398 274350
rect 404778 274226 405398 274294
rect 404778 274170 404874 274226
rect 404930 274170 404998 274226
rect 405054 274170 405122 274226
rect 405178 274170 405246 274226
rect 405302 274170 405398 274226
rect 404778 274102 405398 274170
rect 404778 274046 404874 274102
rect 404930 274046 404998 274102
rect 405054 274046 405122 274102
rect 405178 274046 405246 274102
rect 405302 274046 405398 274102
rect 404778 273978 405398 274046
rect 404778 273922 404874 273978
rect 404930 273922 404998 273978
rect 405054 273922 405122 273978
rect 405178 273922 405246 273978
rect 405302 273922 405398 273978
rect 396620 272998 396676 273008
rect 394828 271312 394884 271322
rect 395612 272278 395668 272288
rect 394828 269758 394884 269768
rect 393820 269038 393876 269048
rect 393484 268858 393540 268868
rect 377778 262294 377874 262350
rect 377930 262294 377998 262350
rect 378054 262294 378122 262350
rect 378178 262294 378246 262350
rect 378302 262294 378398 262350
rect 377778 262226 378398 262294
rect 377778 262170 377874 262226
rect 377930 262170 377998 262226
rect 378054 262170 378122 262226
rect 378178 262170 378246 262226
rect 378302 262170 378398 262226
rect 377778 262102 378398 262170
rect 377778 262046 377874 262102
rect 377930 262046 377998 262102
rect 378054 262046 378122 262102
rect 378178 262046 378246 262102
rect 378302 262046 378398 262102
rect 377778 261978 378398 262046
rect 377778 261922 377874 261978
rect 377930 261922 377998 261978
rect 378054 261922 378122 261978
rect 378178 261922 378246 261978
rect 378302 261922 378398 261978
rect 377778 244350 378398 261922
rect 393260 267418 393316 267428
rect 393260 260372 393316 267362
rect 393372 266698 393428 266708
rect 393372 266308 393428 266642
rect 393372 266242 393428 266252
rect 393372 264898 393428 264908
rect 393372 264786 393428 264796
rect 393484 261492 393540 268802
rect 393596 266698 393652 266708
rect 393596 263638 393652 266642
rect 393596 263572 393652 263582
rect 393484 261426 393540 261436
rect 393820 260398 393876 268982
rect 394828 263060 394884 269702
rect 395052 267092 395108 267102
rect 394828 262994 394884 263004
rect 394940 265076 394996 265086
rect 393820 260332 393876 260342
rect 393260 260306 393316 260316
rect 393148 258958 393204 258968
rect 393148 258418 393204 258902
rect 393148 258352 393204 258362
rect 387168 256350 387488 256384
rect 387168 256294 387238 256350
rect 387294 256294 387362 256350
rect 387418 256294 387488 256350
rect 387168 256226 387488 256294
rect 387168 256170 387238 256226
rect 387294 256170 387362 256226
rect 387418 256170 387488 256226
rect 387168 256102 387488 256170
rect 387168 256046 387238 256102
rect 387294 256046 387362 256102
rect 387418 256046 387488 256102
rect 387168 255978 387488 256046
rect 387168 255922 387238 255978
rect 387294 255922 387362 255978
rect 387418 255922 387488 255978
rect 387168 255888 387488 255922
rect 377778 244294 377874 244350
rect 377930 244294 377998 244350
rect 378054 244294 378122 244350
rect 378178 244294 378246 244350
rect 378302 244294 378398 244350
rect 377778 244226 378398 244294
rect 377778 244170 377874 244226
rect 377930 244170 377998 244226
rect 378054 244170 378122 244226
rect 378178 244170 378246 244226
rect 378302 244170 378398 244226
rect 377778 244102 378398 244170
rect 377778 244046 377874 244102
rect 377930 244046 377998 244102
rect 378054 244046 378122 244102
rect 378178 244046 378246 244102
rect 378302 244046 378398 244102
rect 377778 243978 378398 244046
rect 377778 243922 377874 243978
rect 377930 243922 377998 243978
rect 378054 243922 378122 243978
rect 378178 243922 378246 243978
rect 378302 243922 378398 243978
rect 377778 226350 378398 243922
rect 394940 241556 394996 265020
rect 395052 242676 395108 267036
rect 395612 259588 395668 272222
rect 396620 263732 396676 272942
rect 396620 263666 396676 263676
rect 396844 271738 396900 271748
rect 396844 261716 396900 271682
rect 396956 271558 397012 271568
rect 396956 262388 397012 271502
rect 404012 269108 404068 269118
rect 396956 262322 397012 262332
rect 402332 265076 402388 265086
rect 396844 261650 396900 261660
rect 398972 261716 399028 261726
rect 395612 259522 395668 259532
rect 396620 259700 396676 259710
rect 396620 244468 396676 259644
rect 398972 254998 399028 261660
rect 398972 254932 399028 254942
rect 402332 248518 402388 265020
rect 404012 250138 404068 269052
rect 404012 250072 404068 250082
rect 404778 256350 405398 273922
rect 408498 316350 409118 333922
rect 433808 334350 434128 334384
rect 433808 334294 433878 334350
rect 433934 334294 434002 334350
rect 434058 334294 434128 334350
rect 433808 334226 434128 334294
rect 433808 334170 433878 334226
rect 433934 334170 434002 334226
rect 434058 334170 434128 334226
rect 433808 334102 434128 334170
rect 433808 334046 433878 334102
rect 433934 334046 434002 334102
rect 434058 334046 434128 334102
rect 433808 333978 434128 334046
rect 433808 333922 433878 333978
rect 433934 333922 434002 333978
rect 434058 333922 434128 333978
rect 433808 333888 434128 333922
rect 418448 328350 418768 328384
rect 418448 328294 418518 328350
rect 418574 328294 418642 328350
rect 418698 328294 418768 328350
rect 418448 328226 418768 328294
rect 418448 328170 418518 328226
rect 418574 328170 418642 328226
rect 418698 328170 418768 328226
rect 418448 328102 418768 328170
rect 418448 328046 418518 328102
rect 418574 328046 418642 328102
rect 418698 328046 418768 328102
rect 418448 327978 418768 328046
rect 418448 327922 418518 327978
rect 418574 327922 418642 327978
rect 418698 327922 418768 327978
rect 418448 327888 418768 327922
rect 435498 328350 436118 345922
rect 435498 328294 435594 328350
rect 435650 328294 435718 328350
rect 435774 328294 435842 328350
rect 435898 328294 435966 328350
rect 436022 328294 436118 328350
rect 435498 328226 436118 328294
rect 435498 328170 435594 328226
rect 435650 328170 435718 328226
rect 435774 328170 435842 328226
rect 435898 328170 435966 328226
rect 436022 328170 436118 328226
rect 435498 328102 436118 328170
rect 435498 328046 435594 328102
rect 435650 328046 435718 328102
rect 435774 328046 435842 328102
rect 435898 328046 435966 328102
rect 436022 328046 436118 328102
rect 435498 327978 436118 328046
rect 435498 327922 435594 327978
rect 435650 327922 435718 327978
rect 435774 327922 435842 327978
rect 435898 327922 435966 327978
rect 436022 327922 436118 327978
rect 408498 316294 408594 316350
rect 408650 316294 408718 316350
rect 408774 316294 408842 316350
rect 408898 316294 408966 316350
rect 409022 316294 409118 316350
rect 408498 316226 409118 316294
rect 408498 316170 408594 316226
rect 408650 316170 408718 316226
rect 408774 316170 408842 316226
rect 408898 316170 408966 316226
rect 409022 316170 409118 316226
rect 408498 316102 409118 316170
rect 408498 316046 408594 316102
rect 408650 316046 408718 316102
rect 408774 316046 408842 316102
rect 408898 316046 408966 316102
rect 409022 316046 409118 316102
rect 408498 315978 409118 316046
rect 408498 315922 408594 315978
rect 408650 315922 408718 315978
rect 408774 315922 408842 315978
rect 408898 315922 408966 315978
rect 409022 315922 409118 315978
rect 408498 298350 409118 315922
rect 408498 298294 408594 298350
rect 408650 298294 408718 298350
rect 408774 298294 408842 298350
rect 408898 298294 408966 298350
rect 409022 298294 409118 298350
rect 408498 298226 409118 298294
rect 408498 298170 408594 298226
rect 408650 298170 408718 298226
rect 408774 298170 408842 298226
rect 408898 298170 408966 298226
rect 409022 298170 409118 298226
rect 408498 298102 409118 298170
rect 408498 298046 408594 298102
rect 408650 298046 408718 298102
rect 408774 298046 408842 298102
rect 408898 298046 408966 298102
rect 409022 298046 409118 298102
rect 408498 297978 409118 298046
rect 408498 297922 408594 297978
rect 408650 297922 408718 297978
rect 408774 297922 408842 297978
rect 408898 297922 408966 297978
rect 409022 297922 409118 297978
rect 408498 280350 409118 297922
rect 435498 310350 436118 327922
rect 435498 310294 435594 310350
rect 435650 310294 435718 310350
rect 435774 310294 435842 310350
rect 435898 310294 435966 310350
rect 436022 310294 436118 310350
rect 435498 310226 436118 310294
rect 435498 310170 435594 310226
rect 435650 310170 435718 310226
rect 435774 310170 435842 310226
rect 435898 310170 435966 310226
rect 436022 310170 436118 310226
rect 435498 310102 436118 310170
rect 435498 310046 435594 310102
rect 435650 310046 435718 310102
rect 435774 310046 435842 310102
rect 435898 310046 435966 310102
rect 436022 310046 436118 310102
rect 435498 309978 436118 310046
rect 435498 309922 435594 309978
rect 435650 309922 435718 309978
rect 435774 309922 435842 309978
rect 435898 309922 435966 309978
rect 436022 309922 436118 309978
rect 435498 292350 436118 309922
rect 435498 292294 435594 292350
rect 435650 292294 435718 292350
rect 435774 292294 435842 292350
rect 435898 292294 435966 292350
rect 436022 292294 436118 292350
rect 435498 292226 436118 292294
rect 435498 292170 435594 292226
rect 435650 292170 435718 292226
rect 435774 292170 435842 292226
rect 435898 292170 435966 292226
rect 436022 292170 436118 292226
rect 435498 292102 436118 292170
rect 435498 292046 435594 292102
rect 435650 292046 435718 292102
rect 435774 292046 435842 292102
rect 435898 292046 435966 292102
rect 436022 292046 436118 292102
rect 435498 291978 436118 292046
rect 430108 291956 430164 291966
rect 430108 284788 430164 291900
rect 430108 284722 430164 284732
rect 435498 291922 435594 291978
rect 435650 291922 435718 291978
rect 435774 291922 435842 291978
rect 435898 291922 435966 291978
rect 436022 291922 436118 291978
rect 408498 280294 408594 280350
rect 408650 280294 408718 280350
rect 408774 280294 408842 280350
rect 408898 280294 408966 280350
rect 409022 280294 409118 280350
rect 408498 280226 409118 280294
rect 408498 280170 408594 280226
rect 408650 280170 408718 280226
rect 408774 280170 408842 280226
rect 408898 280170 408966 280226
rect 409022 280170 409118 280226
rect 408498 280102 409118 280170
rect 408498 280046 408594 280102
rect 408650 280046 408718 280102
rect 408774 280046 408842 280102
rect 408898 280046 408966 280102
rect 409022 280046 409118 280102
rect 408498 279978 409118 280046
rect 408498 279922 408594 279978
rect 408650 279922 408718 279978
rect 408774 279922 408842 279978
rect 408898 279922 408966 279978
rect 409022 279922 409118 279978
rect 404778 256294 404874 256350
rect 404930 256294 404998 256350
rect 405054 256294 405122 256350
rect 405178 256294 405246 256350
rect 405302 256294 405398 256350
rect 404778 256226 405398 256294
rect 404778 256170 404874 256226
rect 404930 256170 404998 256226
rect 405054 256170 405122 256226
rect 405178 256170 405246 256226
rect 405302 256170 405398 256226
rect 404778 256102 405398 256170
rect 404778 256046 404874 256102
rect 404930 256046 404998 256102
rect 405054 256046 405122 256102
rect 405178 256046 405246 256102
rect 405302 256046 405398 256102
rect 404778 255978 405398 256046
rect 404778 255922 404874 255978
rect 404930 255922 404998 255978
rect 405054 255922 405122 255978
rect 405178 255922 405246 255978
rect 405302 255922 405398 255978
rect 402332 248452 402388 248462
rect 396620 244402 396676 244412
rect 395052 242610 395108 242620
rect 394940 241490 394996 241500
rect 404778 238350 405398 255922
rect 407372 266420 407428 266430
rect 407372 251758 407428 266364
rect 407372 251692 407428 251702
rect 408498 262350 409118 279922
rect 433808 280350 434128 280384
rect 433808 280294 433878 280350
rect 433934 280294 434002 280350
rect 434058 280294 434128 280350
rect 433808 280226 434128 280294
rect 433808 280170 433878 280226
rect 433934 280170 434002 280226
rect 434058 280170 434128 280226
rect 433808 280102 434128 280170
rect 433808 280046 433878 280102
rect 433934 280046 434002 280102
rect 434058 280046 434128 280102
rect 433808 279978 434128 280046
rect 433808 279922 433878 279978
rect 433934 279922 434002 279978
rect 434058 279922 434128 279978
rect 433808 279888 434128 279922
rect 418448 274350 418768 274384
rect 418448 274294 418518 274350
rect 418574 274294 418642 274350
rect 418698 274294 418768 274350
rect 418448 274226 418768 274294
rect 418448 274170 418518 274226
rect 418574 274170 418642 274226
rect 418698 274170 418768 274226
rect 418448 274102 418768 274170
rect 418448 274046 418518 274102
rect 418574 274046 418642 274102
rect 418698 274046 418768 274102
rect 418448 273978 418768 274046
rect 418448 273922 418518 273978
rect 418574 273922 418642 273978
rect 418698 273922 418768 273978
rect 418448 273888 418768 273922
rect 435498 274350 436118 291922
rect 435498 274294 435594 274350
rect 435650 274294 435718 274350
rect 435774 274294 435842 274350
rect 435898 274294 435966 274350
rect 436022 274294 436118 274350
rect 435498 274226 436118 274294
rect 435498 274170 435594 274226
rect 435650 274170 435718 274226
rect 435774 274170 435842 274226
rect 435898 274170 435966 274226
rect 436022 274170 436118 274226
rect 435498 274102 436118 274170
rect 435498 274046 435594 274102
rect 435650 274046 435718 274102
rect 435774 274046 435842 274102
rect 435898 274046 435966 274102
rect 436022 274046 436118 274102
rect 435498 273978 436118 274046
rect 435498 273922 435594 273978
rect 435650 273922 435718 273978
rect 435774 273922 435842 273978
rect 435898 273922 435966 273978
rect 436022 273922 436118 273978
rect 414652 269578 414708 269588
rect 414652 269484 414708 269500
rect 428316 268858 428372 268868
rect 408498 262294 408594 262350
rect 408650 262294 408718 262350
rect 408774 262294 408842 262350
rect 408898 262294 408966 262350
rect 409022 262294 409118 262350
rect 408498 262226 409118 262294
rect 408498 262170 408594 262226
rect 408650 262170 408718 262226
rect 408774 262170 408842 262226
rect 408898 262170 408966 262226
rect 409022 262170 409118 262226
rect 408498 262102 409118 262170
rect 408498 262046 408594 262102
rect 408650 262046 408718 262102
rect 408774 262046 408842 262102
rect 408898 262046 408966 262102
rect 409022 262046 409118 262102
rect 408498 261978 409118 262046
rect 408498 261922 408594 261978
rect 408650 261922 408718 261978
rect 408774 261922 408842 261978
rect 408898 261922 408966 261978
rect 409022 261922 409118 261978
rect 404778 238294 404874 238350
rect 404930 238294 404998 238350
rect 405054 238294 405122 238350
rect 405178 238294 405246 238350
rect 405302 238294 405398 238350
rect 404778 238226 405398 238294
rect 404778 238170 404874 238226
rect 404930 238170 404998 238226
rect 405054 238170 405122 238226
rect 405178 238170 405246 238226
rect 405302 238170 405398 238226
rect 404778 238102 405398 238170
rect 404778 238046 404874 238102
rect 404930 238046 404998 238102
rect 405054 238046 405122 238102
rect 405178 238046 405246 238102
rect 405302 238046 405398 238102
rect 404778 237978 405398 238046
rect 404778 237922 404874 237978
rect 404930 237922 404998 237978
rect 405054 237922 405122 237978
rect 405178 237922 405246 237978
rect 405302 237922 405398 237978
rect 400652 236516 400708 236526
rect 377778 226294 377874 226350
rect 377930 226294 377998 226350
rect 378054 226294 378122 226350
rect 378178 226294 378246 226350
rect 378302 226294 378398 226350
rect 377778 226226 378398 226294
rect 377778 226170 377874 226226
rect 377930 226170 377998 226226
rect 378054 226170 378122 226226
rect 378178 226170 378246 226226
rect 378302 226170 378398 226226
rect 377778 226102 378398 226170
rect 377778 226046 377874 226102
rect 377930 226046 377998 226102
rect 378054 226046 378122 226102
rect 378178 226046 378246 226102
rect 378302 226046 378398 226102
rect 377778 225978 378398 226046
rect 377778 225922 377874 225978
rect 377930 225922 377998 225978
rect 378054 225922 378122 225978
rect 378178 225922 378246 225978
rect 378302 225922 378398 225978
rect 375788 212884 375844 212894
rect 375788 212660 375844 212828
rect 375788 212594 375844 212604
rect 374058 202294 374154 202350
rect 374210 202294 374278 202350
rect 374334 202294 374402 202350
rect 374458 202294 374526 202350
rect 374582 202294 374678 202350
rect 374058 202226 374678 202294
rect 374058 202170 374154 202226
rect 374210 202170 374278 202226
rect 374334 202170 374402 202226
rect 374458 202170 374526 202226
rect 374582 202170 374678 202226
rect 374058 202102 374678 202170
rect 374058 202046 374154 202102
rect 374210 202046 374278 202102
rect 374334 202046 374402 202102
rect 374458 202046 374526 202102
rect 374582 202046 374678 202102
rect 374058 201978 374678 202046
rect 374058 201922 374154 201978
rect 374210 201922 374278 201978
rect 374334 201922 374402 201978
rect 374458 201922 374526 201978
rect 374582 201922 374678 201978
rect 352716 199018 352772 199028
rect 352716 198548 352772 198962
rect 352716 198482 352772 198492
rect 351820 195238 351876 195248
rect 351820 192724 351876 195182
rect 351820 192658 351876 192668
rect 347058 190294 347154 190350
rect 347210 190294 347278 190350
rect 347334 190294 347402 190350
rect 347458 190294 347526 190350
rect 347582 190294 347678 190350
rect 347058 190226 347678 190294
rect 347058 190170 347154 190226
rect 347210 190170 347278 190226
rect 347334 190170 347402 190226
rect 347458 190170 347526 190226
rect 347582 190170 347678 190226
rect 347058 190102 347678 190170
rect 347058 190046 347154 190102
rect 347210 190046 347278 190102
rect 347334 190046 347402 190102
rect 347458 190046 347526 190102
rect 347582 190046 347678 190102
rect 347058 189978 347678 190046
rect 347058 189922 347154 189978
rect 347210 189922 347278 189978
rect 347334 189922 347402 189978
rect 347458 189922 347526 189978
rect 347582 189922 347678 189978
rect 346108 188468 346164 188478
rect 346108 185556 346164 188412
rect 346108 185490 346164 185500
rect 343338 184294 343434 184350
rect 343490 184294 343558 184350
rect 343614 184294 343682 184350
rect 343738 184294 343806 184350
rect 343862 184294 343958 184350
rect 343338 184226 343958 184294
rect 343338 184170 343434 184226
rect 343490 184170 343558 184226
rect 343614 184170 343682 184226
rect 343738 184170 343806 184226
rect 343862 184170 343958 184226
rect 343338 184102 343958 184170
rect 343338 184046 343434 184102
rect 343490 184046 343558 184102
rect 343614 184046 343682 184102
rect 343738 184046 343806 184102
rect 343862 184046 343958 184102
rect 343338 183978 343958 184046
rect 343338 183922 343434 183978
rect 343490 183922 343558 183978
rect 343614 183922 343682 183978
rect 343738 183922 343806 183978
rect 343862 183922 343958 183978
rect 338492 181076 338548 181086
rect 335356 177716 335412 177726
rect 334460 176596 334516 176606
rect 334460 173908 334516 176540
rect 334460 173842 334516 173852
rect 335356 158788 335412 177660
rect 336028 171556 336084 171566
rect 336028 170548 336084 171500
rect 336028 170482 336084 170492
rect 335356 158722 335412 158732
rect 338492 155540 338548 181020
rect 341852 175476 341908 175486
rect 338940 169316 338996 169326
rect 338604 164836 338660 164846
rect 338604 157220 338660 164780
rect 338940 160580 338996 169260
rect 341852 163828 341908 175420
rect 341852 163762 341908 163772
rect 343338 166350 343958 183922
rect 343338 166294 343434 166350
rect 343490 166294 343558 166350
rect 343614 166294 343682 166350
rect 343738 166294 343806 166350
rect 343862 166294 343958 166350
rect 343338 166226 343958 166294
rect 343338 166170 343434 166226
rect 343490 166170 343558 166226
rect 343614 166170 343682 166226
rect 343738 166170 343806 166226
rect 343862 166170 343958 166226
rect 343338 166102 343958 166170
rect 343338 166046 343434 166102
rect 343490 166046 343558 166102
rect 343614 166046 343682 166102
rect 343738 166046 343806 166102
rect 343862 166046 343958 166102
rect 343338 165978 343958 166046
rect 343338 165922 343434 165978
rect 343490 165922 343558 165978
rect 343614 165922 343682 165978
rect 343738 165922 343806 165978
rect 343862 165922 343958 165978
rect 338940 160514 338996 160524
rect 338604 157154 338660 157164
rect 338492 155474 338548 155484
rect 341852 156436 341908 156446
rect 334348 142996 334404 143006
rect 334348 140644 334404 142940
rect 334460 142548 334516 142558
rect 334460 141764 334516 142492
rect 334460 141698 334516 141708
rect 334348 140578 334404 140588
rect 334460 134596 334516 134606
rect 334460 133498 334516 134540
rect 334460 133432 334516 133442
rect 334460 132356 334516 132366
rect 334348 131796 334404 131806
rect 334348 131158 334404 131740
rect 334460 131338 334516 132300
rect 334460 131272 334516 131282
rect 338492 131236 338548 131246
rect 334460 131158 334516 131168
rect 334348 131102 334460 131158
rect 334460 131092 334516 131102
rect 334460 126838 334516 126848
rect 334460 126756 334516 126782
rect 334460 126690 334516 126700
rect 334460 125636 334516 125646
rect 334460 125218 334516 125580
rect 334460 125152 334516 125162
rect 338492 124318 338548 131180
rect 341852 129332 341908 156380
rect 343338 148350 343958 165922
rect 343338 148294 343434 148350
rect 343490 148294 343558 148350
rect 343614 148294 343682 148350
rect 343738 148294 343806 148350
rect 343862 148294 343958 148350
rect 343338 148226 343958 148294
rect 343338 148170 343434 148226
rect 343490 148170 343558 148226
rect 343614 148170 343682 148226
rect 343738 148170 343806 148226
rect 343862 148170 343958 148226
rect 343338 148102 343958 148170
rect 343338 148046 343434 148102
rect 343490 148046 343558 148102
rect 343614 148046 343682 148102
rect 343738 148046 343806 148102
rect 343862 148046 343958 148102
rect 343338 147978 343958 148046
rect 343338 147922 343434 147978
rect 343490 147922 343558 147978
rect 343614 147922 343682 147978
rect 343738 147922 343806 147978
rect 343862 147922 343958 147978
rect 343338 130350 343958 147922
rect 345212 179956 345268 179966
rect 345212 140308 345268 179900
rect 347058 172350 347678 189922
rect 347788 192538 347844 192548
rect 347788 189476 347844 192482
rect 371808 190350 372128 190384
rect 371808 190294 371878 190350
rect 371934 190294 372002 190350
rect 372058 190294 372128 190350
rect 371808 190226 372128 190294
rect 371808 190170 371878 190226
rect 371934 190170 372002 190226
rect 372058 190170 372128 190226
rect 371808 190102 372128 190170
rect 371808 190046 371878 190102
rect 371934 190046 372002 190102
rect 372058 190046 372128 190102
rect 371808 189978 372128 190046
rect 371808 189922 371878 189978
rect 371934 189922 372002 189978
rect 372058 189922 372128 189978
rect 371808 189888 372128 189922
rect 347788 189410 347844 189420
rect 356448 184350 356768 184384
rect 356448 184294 356518 184350
rect 356574 184294 356642 184350
rect 356698 184294 356768 184350
rect 356448 184226 356768 184294
rect 356448 184170 356518 184226
rect 356574 184170 356642 184226
rect 356698 184170 356768 184226
rect 356448 184102 356768 184170
rect 356448 184046 356518 184102
rect 356574 184046 356642 184102
rect 356698 184046 356768 184102
rect 356448 183978 356768 184046
rect 356448 183922 356518 183978
rect 356574 183922 356642 183978
rect 356698 183922 356768 183978
rect 356448 183888 356768 183922
rect 374058 184350 374678 201922
rect 374058 184294 374154 184350
rect 374210 184294 374278 184350
rect 374334 184294 374402 184350
rect 374458 184294 374526 184350
rect 374582 184294 374678 184350
rect 374058 184226 374678 184294
rect 374058 184170 374154 184226
rect 374210 184170 374278 184226
rect 374334 184170 374402 184226
rect 374458 184170 374526 184226
rect 374582 184170 374678 184226
rect 374058 184102 374678 184170
rect 374058 184046 374154 184102
rect 374210 184046 374278 184102
rect 374334 184046 374402 184102
rect 374458 184046 374526 184102
rect 374582 184046 374678 184102
rect 374058 183978 374678 184046
rect 374058 183922 374154 183978
rect 374210 183922 374278 183978
rect 374334 183922 374402 183978
rect 374458 183922 374526 183978
rect 374582 183922 374678 183978
rect 350252 177156 350308 177166
rect 347058 172294 347154 172350
rect 347210 172294 347278 172350
rect 347334 172294 347402 172350
rect 347458 172294 347526 172350
rect 347582 172294 347678 172350
rect 347058 172226 347678 172294
rect 347058 172170 347154 172226
rect 347210 172170 347278 172226
rect 347334 172170 347402 172226
rect 347458 172170 347526 172226
rect 347582 172170 347678 172226
rect 345436 172116 345492 172126
rect 345436 140420 345492 172060
rect 345436 140354 345492 140364
rect 347058 172102 347678 172170
rect 347058 172046 347154 172102
rect 347210 172046 347278 172102
rect 347334 172046 347402 172102
rect 347458 172046 347526 172102
rect 347582 172046 347678 172102
rect 347058 171978 347678 172046
rect 347058 171922 347154 171978
rect 347210 171922 347278 171978
rect 347334 171922 347402 171978
rect 347458 171922 347526 171978
rect 347582 171922 347678 171978
rect 347058 154350 347678 171922
rect 348572 176036 348628 176046
rect 348572 157108 348628 175980
rect 348572 157042 348628 157052
rect 347058 154294 347154 154350
rect 347210 154294 347278 154350
rect 347334 154294 347402 154350
rect 347458 154294 347526 154350
rect 347582 154294 347678 154350
rect 347058 154226 347678 154294
rect 347058 154170 347154 154226
rect 347210 154170 347278 154226
rect 347334 154170 347402 154226
rect 347458 154170 347526 154226
rect 347582 154170 347678 154226
rect 347058 154102 347678 154170
rect 347058 154046 347154 154102
rect 347210 154046 347278 154102
rect 347334 154046 347402 154102
rect 347458 154046 347526 154102
rect 347582 154046 347678 154102
rect 347058 153978 347678 154046
rect 347058 153922 347154 153978
rect 347210 153922 347278 153978
rect 347334 153922 347402 153978
rect 347458 153922 347526 153978
rect 347582 153922 347678 153978
rect 345212 140242 345268 140252
rect 347058 136350 347678 153922
rect 350252 141988 350308 177100
rect 351932 174916 351988 174926
rect 350364 172676 350420 172686
rect 350364 143668 350420 172620
rect 351932 155428 351988 174860
rect 356972 166516 357028 166526
rect 351932 155362 351988 155372
rect 352044 158676 352100 158686
rect 350364 143602 350420 143612
rect 350252 141922 350308 141932
rect 352044 140868 352100 158620
rect 356972 155652 357028 166460
rect 374058 166350 374678 183922
rect 374058 166294 374154 166350
rect 374210 166294 374278 166350
rect 374334 166294 374402 166350
rect 374458 166294 374526 166350
rect 374582 166294 374678 166350
rect 374058 166226 374678 166294
rect 374058 166170 374154 166226
rect 374210 166170 374278 166226
rect 374334 166170 374402 166226
rect 374458 166170 374526 166226
rect 374582 166170 374678 166226
rect 374058 166102 374678 166170
rect 374058 166046 374154 166102
rect 374210 166046 374278 166102
rect 374334 166046 374402 166102
rect 374458 166046 374526 166102
rect 374582 166046 374678 166102
rect 374058 165978 374678 166046
rect 374058 165922 374154 165978
rect 374210 165922 374278 165978
rect 374334 165922 374402 165978
rect 374458 165922 374526 165978
rect 374582 165922 374678 165978
rect 356972 155586 357028 155596
rect 357196 155876 357252 155886
rect 357196 143780 357252 155820
rect 357196 143714 357252 143724
rect 374058 148350 374678 165922
rect 374058 148294 374154 148350
rect 374210 148294 374278 148350
rect 374334 148294 374402 148350
rect 374458 148294 374526 148350
rect 374582 148294 374678 148350
rect 374058 148226 374678 148294
rect 374058 148170 374154 148226
rect 374210 148170 374278 148226
rect 374334 148170 374402 148226
rect 374458 148170 374526 148226
rect 374582 148170 374678 148226
rect 374058 148102 374678 148170
rect 374058 148046 374154 148102
rect 374210 148046 374278 148102
rect 374334 148046 374402 148102
rect 374458 148046 374526 148102
rect 374582 148046 374678 148102
rect 374058 147978 374678 148046
rect 374058 147922 374154 147978
rect 374210 147922 374278 147978
rect 374334 147922 374402 147978
rect 374458 147922 374526 147978
rect 374582 147922 374678 147978
rect 352044 140802 352100 140812
rect 347058 136294 347154 136350
rect 347210 136294 347278 136350
rect 347334 136294 347402 136350
rect 347458 136294 347526 136350
rect 347582 136294 347678 136350
rect 347058 136226 347678 136294
rect 347058 136170 347154 136226
rect 347210 136170 347278 136226
rect 347334 136170 347402 136226
rect 347458 136170 347526 136226
rect 347582 136170 347678 136226
rect 347058 136102 347678 136170
rect 347058 136046 347154 136102
rect 347210 136046 347278 136102
rect 347334 136046 347402 136102
rect 347458 136046 347526 136102
rect 347582 136046 347678 136102
rect 347058 135978 347678 136046
rect 347058 135922 347154 135978
rect 347210 135922 347278 135978
rect 347334 135922 347402 135978
rect 347458 135922 347526 135978
rect 347582 135922 347678 135978
rect 343338 130294 343434 130350
rect 343490 130294 343558 130350
rect 343614 130294 343682 130350
rect 343738 130294 343806 130350
rect 343862 130294 343958 130350
rect 343338 130226 343958 130294
rect 343338 130170 343434 130226
rect 343490 130170 343558 130226
rect 343614 130170 343682 130226
rect 343738 130170 343806 130226
rect 343862 130170 343958 130226
rect 341852 129266 341908 129276
rect 342188 130116 342244 130126
rect 338492 124252 338548 124262
rect 341964 127316 342020 127326
rect 336812 123396 336868 123406
rect 335244 117236 335300 117246
rect 335132 112756 335188 112766
rect 334460 102116 334516 102126
rect 334460 99988 334516 102060
rect 334460 99922 334516 99932
rect 334572 101556 334628 101566
rect 334348 99876 334404 99886
rect 334348 98308 334404 99820
rect 334348 98242 334404 98252
rect 334460 98196 334516 98206
rect 334460 97188 334516 98140
rect 334460 97122 334516 97132
rect 334572 95060 334628 101500
rect 334572 94994 334628 95004
rect 334684 99316 334740 99326
rect 334684 91700 334740 99260
rect 334684 91634 334740 91644
rect 334460 75796 334516 75806
rect 334348 75236 334404 75246
rect 334348 73444 334404 75180
rect 334460 74788 334516 75740
rect 334460 74722 334516 74732
rect 334572 74116 334628 74126
rect 334348 73378 334404 73388
rect 334460 73556 334516 73566
rect 333452 73154 333508 73164
rect 263788 73042 263844 73052
rect 334460 71652 334516 73500
rect 334460 71586 334516 71596
rect 262892 69794 262948 69804
rect 261324 69682 261380 69692
rect 334572 68180 334628 74060
rect 335132 73332 335188 112700
rect 335244 103348 335300 117180
rect 335468 112196 335524 112206
rect 335244 103282 335300 103292
rect 335356 110516 335412 110526
rect 335244 100996 335300 101006
rect 335244 84980 335300 100940
rect 335356 91588 335412 110460
rect 335468 101108 335524 112140
rect 335468 101042 335524 101052
rect 335916 106596 335972 106606
rect 335916 100884 335972 106540
rect 335916 100818 335972 100828
rect 335356 91522 335412 91532
rect 335244 84914 335300 84924
rect 335132 73266 335188 73276
rect 336812 69748 336868 123340
rect 337036 122276 337092 122286
rect 336924 120036 336980 120046
rect 336924 71428 336980 119980
rect 337036 73108 337092 122220
rect 341852 120596 341908 120606
rect 338716 118356 338772 118366
rect 338604 116676 338660 116686
rect 337036 73042 337092 73052
rect 338492 111636 338548 111646
rect 336924 71362 336980 71372
rect 338492 69972 338548 111580
rect 338604 79828 338660 116620
rect 338716 96628 338772 118300
rect 338716 96562 338772 96572
rect 338940 109396 338996 109406
rect 338940 93380 338996 109340
rect 340396 106036 340452 106046
rect 338940 93314 338996 93324
rect 340172 97636 340228 97646
rect 338604 79762 338660 79772
rect 338492 69906 338548 69916
rect 336812 69682 336868 69692
rect 334572 68114 334628 68124
rect 272448 58350 272768 58384
rect 272448 58294 272518 58350
rect 272574 58294 272642 58350
rect 272698 58294 272768 58350
rect 272448 58226 272768 58294
rect 272448 58170 272518 58226
rect 272574 58170 272642 58226
rect 272698 58170 272768 58226
rect 272448 58102 272768 58170
rect 272448 58046 272518 58102
rect 272574 58046 272642 58102
rect 272698 58046 272768 58102
rect 272448 57978 272768 58046
rect 272448 57922 272518 57978
rect 272574 57922 272642 57978
rect 272698 57922 272768 57978
rect 272448 57888 272768 57922
rect 281898 58350 282518 68098
rect 281898 58294 281994 58350
rect 282050 58294 282118 58350
rect 282174 58294 282242 58350
rect 282298 58294 282366 58350
rect 282422 58294 282518 58350
rect 281898 58226 282518 58294
rect 281898 58170 281994 58226
rect 282050 58170 282118 58226
rect 282174 58170 282242 58226
rect 282298 58170 282366 58226
rect 282422 58170 282518 58226
rect 281898 58102 282518 58170
rect 281898 58046 281994 58102
rect 282050 58046 282118 58102
rect 282174 58046 282242 58102
rect 282298 58046 282366 58102
rect 282422 58046 282518 58102
rect 281898 57978 282518 58046
rect 281898 57922 281994 57978
rect 282050 57922 282118 57978
rect 282174 57922 282242 57978
rect 282298 57922 282366 57978
rect 282422 57922 282518 57978
rect 261212 52098 261268 52108
rect 270060 55558 270116 55568
rect 258188 47394 258244 47404
rect 254898 46294 254994 46350
rect 255050 46294 255118 46350
rect 255174 46294 255242 46350
rect 255298 46294 255366 46350
rect 255422 46294 255518 46350
rect 254898 46226 255518 46294
rect 254898 46170 254994 46226
rect 255050 46170 255118 46226
rect 255174 46170 255242 46226
rect 255298 46170 255366 46226
rect 255422 46170 255518 46226
rect 254898 46102 255518 46170
rect 254898 46046 254994 46102
rect 255050 46046 255118 46102
rect 255174 46046 255242 46102
rect 255298 46046 255366 46102
rect 255422 46046 255518 46102
rect 254898 45978 255518 46046
rect 254898 45922 254994 45978
rect 255050 45922 255118 45978
rect 255174 45922 255242 45978
rect 255298 45922 255366 45978
rect 255422 45922 255518 45978
rect 251178 40294 251274 40350
rect 251330 40294 251398 40350
rect 251454 40294 251522 40350
rect 251578 40294 251646 40350
rect 251702 40294 251798 40350
rect 251178 40226 251798 40294
rect 251178 40170 251274 40226
rect 251330 40170 251398 40226
rect 251454 40170 251522 40226
rect 251578 40170 251646 40226
rect 251702 40170 251798 40226
rect 251178 40102 251798 40170
rect 251178 40046 251274 40102
rect 251330 40046 251398 40102
rect 251454 40046 251522 40102
rect 251578 40046 251646 40102
rect 251702 40046 251798 40102
rect 251178 39978 251798 40046
rect 251178 39922 251274 39978
rect 251330 39922 251398 39978
rect 251454 39922 251522 39978
rect 251578 39922 251646 39978
rect 251702 39922 251798 39978
rect 224178 28294 224274 28350
rect 224330 28294 224398 28350
rect 224454 28294 224522 28350
rect 224578 28294 224646 28350
rect 224702 28294 224798 28350
rect 224178 28226 224798 28294
rect 224178 28170 224274 28226
rect 224330 28170 224398 28226
rect 224454 28170 224522 28226
rect 224578 28170 224646 28226
rect 224702 28170 224798 28226
rect 224178 28102 224798 28170
rect 224178 28046 224274 28102
rect 224330 28046 224398 28102
rect 224454 28046 224522 28102
rect 224578 28046 224646 28102
rect 224702 28046 224798 28102
rect 224178 27978 224798 28046
rect 224178 27922 224274 27978
rect 224330 27922 224398 27978
rect 224454 27922 224522 27978
rect 224578 27922 224646 27978
rect 224702 27922 224798 27978
rect 224178 10350 224798 27922
rect 224178 10294 224274 10350
rect 224330 10294 224398 10350
rect 224454 10294 224522 10350
rect 224578 10294 224646 10350
rect 224702 10294 224798 10350
rect 224178 10226 224798 10294
rect 224178 10170 224274 10226
rect 224330 10170 224398 10226
rect 224454 10170 224522 10226
rect 224578 10170 224646 10226
rect 224702 10170 224798 10226
rect 224178 10102 224798 10170
rect 224178 10046 224274 10102
rect 224330 10046 224398 10102
rect 224454 10046 224522 10102
rect 224578 10046 224646 10102
rect 224702 10046 224798 10102
rect 224178 9978 224798 10046
rect 224178 9922 224274 9978
rect 224330 9922 224398 9978
rect 224454 9922 224522 9978
rect 224578 9922 224646 9978
rect 224702 9922 224798 9978
rect 224178 -1120 224798 9922
rect 224178 -1176 224274 -1120
rect 224330 -1176 224398 -1120
rect 224454 -1176 224522 -1120
rect 224578 -1176 224646 -1120
rect 224702 -1176 224798 -1120
rect 224178 -1244 224798 -1176
rect 224178 -1300 224274 -1244
rect 224330 -1300 224398 -1244
rect 224454 -1300 224522 -1244
rect 224578 -1300 224646 -1244
rect 224702 -1300 224798 -1244
rect 224178 -1368 224798 -1300
rect 224178 -1424 224274 -1368
rect 224330 -1424 224398 -1368
rect 224454 -1424 224522 -1368
rect 224578 -1424 224646 -1368
rect 224702 -1424 224798 -1368
rect 224178 -1492 224798 -1424
rect 224178 -1548 224274 -1492
rect 224330 -1548 224398 -1492
rect 224454 -1548 224522 -1492
rect 224578 -1548 224646 -1492
rect 224702 -1548 224798 -1492
rect 224178 -1644 224798 -1548
rect 251178 22350 251798 39922
rect 251178 22294 251274 22350
rect 251330 22294 251398 22350
rect 251454 22294 251522 22350
rect 251578 22294 251646 22350
rect 251702 22294 251798 22350
rect 251178 22226 251798 22294
rect 251178 22170 251274 22226
rect 251330 22170 251398 22226
rect 251454 22170 251522 22226
rect 251578 22170 251646 22226
rect 251702 22170 251798 22226
rect 251178 22102 251798 22170
rect 251178 22046 251274 22102
rect 251330 22046 251398 22102
rect 251454 22046 251522 22102
rect 251578 22046 251646 22102
rect 251702 22046 251798 22102
rect 251178 21978 251798 22046
rect 251178 21922 251274 21978
rect 251330 21922 251398 21978
rect 251454 21922 251522 21978
rect 251578 21922 251646 21978
rect 251702 21922 251798 21978
rect 251178 4350 251798 21922
rect 251178 4294 251274 4350
rect 251330 4294 251398 4350
rect 251454 4294 251522 4350
rect 251578 4294 251646 4350
rect 251702 4294 251798 4350
rect 251178 4226 251798 4294
rect 251178 4170 251274 4226
rect 251330 4170 251398 4226
rect 251454 4170 251522 4226
rect 251578 4170 251646 4226
rect 251702 4170 251798 4226
rect 251178 4102 251798 4170
rect 251178 4046 251274 4102
rect 251330 4046 251398 4102
rect 251454 4046 251522 4102
rect 251578 4046 251646 4102
rect 251702 4046 251798 4102
rect 251178 3978 251798 4046
rect 251178 3922 251274 3978
rect 251330 3922 251398 3978
rect 251454 3922 251522 3978
rect 251578 3922 251646 3978
rect 251702 3922 251798 3978
rect 251178 -160 251798 3922
rect 251178 -216 251274 -160
rect 251330 -216 251398 -160
rect 251454 -216 251522 -160
rect 251578 -216 251646 -160
rect 251702 -216 251798 -160
rect 251178 -284 251798 -216
rect 251178 -340 251274 -284
rect 251330 -340 251398 -284
rect 251454 -340 251522 -284
rect 251578 -340 251646 -284
rect 251702 -340 251798 -284
rect 251178 -408 251798 -340
rect 251178 -464 251274 -408
rect 251330 -464 251398 -408
rect 251454 -464 251522 -408
rect 251578 -464 251646 -408
rect 251702 -464 251798 -408
rect 251178 -532 251798 -464
rect 251178 -588 251274 -532
rect 251330 -588 251398 -532
rect 251454 -588 251522 -532
rect 251578 -588 251646 -532
rect 251702 -588 251798 -532
rect 251178 -1644 251798 -588
rect 254898 28350 255518 45922
rect 270060 29988 270116 55502
rect 272448 40350 272768 40384
rect 272448 40294 272518 40350
rect 272574 40294 272642 40350
rect 272698 40294 272768 40350
rect 272448 40226 272768 40294
rect 272448 40170 272518 40226
rect 272574 40170 272642 40226
rect 272698 40170 272768 40226
rect 272448 40102 272768 40170
rect 272448 40046 272518 40102
rect 272574 40046 272642 40102
rect 272698 40046 272768 40102
rect 272448 39978 272768 40046
rect 272448 39922 272518 39978
rect 272574 39922 272642 39978
rect 272698 39922 272768 39978
rect 272448 39888 272768 39922
rect 281898 40350 282518 57922
rect 281898 40294 281994 40350
rect 282050 40294 282118 40350
rect 282174 40294 282242 40350
rect 282298 40294 282366 40350
rect 282422 40294 282518 40350
rect 281898 40226 282518 40294
rect 281898 40170 281994 40226
rect 282050 40170 282118 40226
rect 282174 40170 282242 40226
rect 282298 40170 282366 40226
rect 282422 40170 282518 40226
rect 281898 40102 282518 40170
rect 281898 40046 281994 40102
rect 282050 40046 282118 40102
rect 282174 40046 282242 40102
rect 282298 40046 282366 40102
rect 282422 40046 282518 40102
rect 281898 39978 282518 40046
rect 281898 39922 281994 39978
rect 282050 39922 282118 39978
rect 282174 39922 282242 39978
rect 282298 39922 282366 39978
rect 282422 39922 282518 39978
rect 270060 29922 270116 29932
rect 254898 28294 254994 28350
rect 255050 28294 255118 28350
rect 255174 28294 255242 28350
rect 255298 28294 255366 28350
rect 255422 28294 255518 28350
rect 254898 28226 255518 28294
rect 254898 28170 254994 28226
rect 255050 28170 255118 28226
rect 255174 28170 255242 28226
rect 255298 28170 255366 28226
rect 255422 28170 255518 28226
rect 254898 28102 255518 28170
rect 254898 28046 254994 28102
rect 255050 28046 255118 28102
rect 255174 28046 255242 28102
rect 255298 28046 255366 28102
rect 255422 28046 255518 28102
rect 254898 27978 255518 28046
rect 254898 27922 254994 27978
rect 255050 27922 255118 27978
rect 255174 27922 255242 27978
rect 255298 27922 255366 27978
rect 255422 27922 255518 27978
rect 254898 10350 255518 27922
rect 254898 10294 254994 10350
rect 255050 10294 255118 10350
rect 255174 10294 255242 10350
rect 255298 10294 255366 10350
rect 255422 10294 255518 10350
rect 254898 10226 255518 10294
rect 254898 10170 254994 10226
rect 255050 10170 255118 10226
rect 255174 10170 255242 10226
rect 255298 10170 255366 10226
rect 255422 10170 255518 10226
rect 254898 10102 255518 10170
rect 254898 10046 254994 10102
rect 255050 10046 255118 10102
rect 255174 10046 255242 10102
rect 255298 10046 255366 10102
rect 255422 10046 255518 10102
rect 254898 9978 255518 10046
rect 254898 9922 254994 9978
rect 255050 9922 255118 9978
rect 255174 9922 255242 9978
rect 255298 9922 255366 9978
rect 255422 9922 255518 9978
rect 254898 -1120 255518 9922
rect 254898 -1176 254994 -1120
rect 255050 -1176 255118 -1120
rect 255174 -1176 255242 -1120
rect 255298 -1176 255366 -1120
rect 255422 -1176 255518 -1120
rect 254898 -1244 255518 -1176
rect 254898 -1300 254994 -1244
rect 255050 -1300 255118 -1244
rect 255174 -1300 255242 -1244
rect 255298 -1300 255366 -1244
rect 255422 -1300 255518 -1244
rect 254898 -1368 255518 -1300
rect 254898 -1424 254994 -1368
rect 255050 -1424 255118 -1368
rect 255174 -1424 255242 -1368
rect 255298 -1424 255366 -1368
rect 255422 -1424 255518 -1368
rect 254898 -1492 255518 -1424
rect 254898 -1548 254994 -1492
rect 255050 -1548 255118 -1492
rect 255174 -1548 255242 -1492
rect 255298 -1548 255366 -1492
rect 255422 -1548 255518 -1492
rect 254898 -1644 255518 -1548
rect 281898 22350 282518 39922
rect 281898 22294 281994 22350
rect 282050 22294 282118 22350
rect 282174 22294 282242 22350
rect 282298 22294 282366 22350
rect 282422 22294 282518 22350
rect 281898 22226 282518 22294
rect 281898 22170 281994 22226
rect 282050 22170 282118 22226
rect 282174 22170 282242 22226
rect 282298 22170 282366 22226
rect 282422 22170 282518 22226
rect 281898 22102 282518 22170
rect 281898 22046 281994 22102
rect 282050 22046 282118 22102
rect 282174 22046 282242 22102
rect 282298 22046 282366 22102
rect 282422 22046 282518 22102
rect 281898 21978 282518 22046
rect 281898 21922 281994 21978
rect 282050 21922 282118 21978
rect 282174 21922 282242 21978
rect 282298 21922 282366 21978
rect 282422 21922 282518 21978
rect 281898 4350 282518 21922
rect 281898 4294 281994 4350
rect 282050 4294 282118 4350
rect 282174 4294 282242 4350
rect 282298 4294 282366 4350
rect 282422 4294 282518 4350
rect 281898 4226 282518 4294
rect 281898 4170 281994 4226
rect 282050 4170 282118 4226
rect 282174 4170 282242 4226
rect 282298 4170 282366 4226
rect 282422 4170 282518 4226
rect 281898 4102 282518 4170
rect 281898 4046 281994 4102
rect 282050 4046 282118 4102
rect 282174 4046 282242 4102
rect 282298 4046 282366 4102
rect 282422 4046 282518 4102
rect 281898 3978 282518 4046
rect 281898 3922 281994 3978
rect 282050 3922 282118 3978
rect 282174 3922 282242 3978
rect 282298 3922 282366 3978
rect 282422 3922 282518 3978
rect 281898 -160 282518 3922
rect 281898 -216 281994 -160
rect 282050 -216 282118 -160
rect 282174 -216 282242 -160
rect 282298 -216 282366 -160
rect 282422 -216 282518 -160
rect 281898 -284 282518 -216
rect 281898 -340 281994 -284
rect 282050 -340 282118 -284
rect 282174 -340 282242 -284
rect 282298 -340 282366 -284
rect 282422 -340 282518 -284
rect 281898 -408 282518 -340
rect 281898 -464 281994 -408
rect 282050 -464 282118 -408
rect 282174 -464 282242 -408
rect 282298 -464 282366 -408
rect 282422 -464 282518 -408
rect 281898 -532 282518 -464
rect 281898 -588 281994 -532
rect 282050 -588 282118 -532
rect 282174 -588 282242 -532
rect 282298 -588 282366 -532
rect 282422 -588 282518 -532
rect 281898 -1644 282518 -588
rect 285618 64350 286238 68098
rect 285618 64294 285714 64350
rect 285770 64294 285838 64350
rect 285894 64294 285962 64350
rect 286018 64294 286086 64350
rect 286142 64294 286238 64350
rect 285618 64226 286238 64294
rect 285618 64170 285714 64226
rect 285770 64170 285838 64226
rect 285894 64170 285962 64226
rect 286018 64170 286086 64226
rect 286142 64170 286238 64226
rect 285618 64102 286238 64170
rect 285618 64046 285714 64102
rect 285770 64046 285838 64102
rect 285894 64046 285962 64102
rect 286018 64046 286086 64102
rect 286142 64046 286238 64102
rect 285618 63978 286238 64046
rect 285618 63922 285714 63978
rect 285770 63922 285838 63978
rect 285894 63922 285962 63978
rect 286018 63922 286086 63978
rect 286142 63922 286238 63978
rect 285618 46350 286238 63922
rect 287808 64350 288128 64384
rect 287808 64294 287878 64350
rect 287934 64294 288002 64350
rect 288058 64294 288128 64350
rect 287808 64226 288128 64294
rect 287808 64170 287878 64226
rect 287934 64170 288002 64226
rect 288058 64170 288128 64226
rect 287808 64102 288128 64170
rect 287808 64046 287878 64102
rect 287934 64046 288002 64102
rect 288058 64046 288128 64102
rect 287808 63978 288128 64046
rect 287808 63922 287878 63978
rect 287934 63922 288002 63978
rect 288058 63922 288128 63978
rect 287808 63888 288128 63922
rect 303168 58350 303488 58384
rect 303168 58294 303238 58350
rect 303294 58294 303362 58350
rect 303418 58294 303488 58350
rect 303168 58226 303488 58294
rect 303168 58170 303238 58226
rect 303294 58170 303362 58226
rect 303418 58170 303488 58226
rect 303168 58102 303488 58170
rect 303168 58046 303238 58102
rect 303294 58046 303362 58102
rect 303418 58046 303488 58102
rect 303168 57978 303488 58046
rect 303168 57922 303238 57978
rect 303294 57922 303362 57978
rect 303418 57922 303488 57978
rect 303168 57888 303488 57922
rect 312618 58350 313238 68098
rect 312618 58294 312714 58350
rect 312770 58294 312838 58350
rect 312894 58294 312962 58350
rect 313018 58294 313086 58350
rect 313142 58294 313238 58350
rect 312618 58226 313238 58294
rect 312618 58170 312714 58226
rect 312770 58170 312838 58226
rect 312894 58170 312962 58226
rect 313018 58170 313086 58226
rect 313142 58170 313238 58226
rect 312618 58102 313238 58170
rect 312618 58046 312714 58102
rect 312770 58046 312838 58102
rect 312894 58046 312962 58102
rect 313018 58046 313086 58102
rect 313142 58046 313238 58102
rect 312618 57978 313238 58046
rect 312618 57922 312714 57978
rect 312770 57922 312838 57978
rect 312894 57922 312962 57978
rect 313018 57922 313086 57978
rect 313142 57922 313238 57978
rect 285618 46294 285714 46350
rect 285770 46294 285838 46350
rect 285894 46294 285962 46350
rect 286018 46294 286086 46350
rect 286142 46294 286238 46350
rect 285618 46226 286238 46294
rect 285618 46170 285714 46226
rect 285770 46170 285838 46226
rect 285894 46170 285962 46226
rect 286018 46170 286086 46226
rect 286142 46170 286238 46226
rect 285618 46102 286238 46170
rect 285618 46046 285714 46102
rect 285770 46046 285838 46102
rect 285894 46046 285962 46102
rect 286018 46046 286086 46102
rect 286142 46046 286238 46102
rect 285618 45978 286238 46046
rect 285618 45922 285714 45978
rect 285770 45922 285838 45978
rect 285894 45922 285962 45978
rect 286018 45922 286086 45978
rect 286142 45922 286238 45978
rect 285618 28350 286238 45922
rect 287808 46350 288128 46384
rect 287808 46294 287878 46350
rect 287934 46294 288002 46350
rect 288058 46294 288128 46350
rect 287808 46226 288128 46294
rect 287808 46170 287878 46226
rect 287934 46170 288002 46226
rect 288058 46170 288128 46226
rect 287808 46102 288128 46170
rect 287808 46046 287878 46102
rect 287934 46046 288002 46102
rect 288058 46046 288128 46102
rect 287808 45978 288128 46046
rect 287808 45922 287878 45978
rect 287934 45922 288002 45978
rect 288058 45922 288128 45978
rect 287808 45888 288128 45922
rect 303168 40350 303488 40384
rect 303168 40294 303238 40350
rect 303294 40294 303362 40350
rect 303418 40294 303488 40350
rect 303168 40226 303488 40294
rect 303168 40170 303238 40226
rect 303294 40170 303362 40226
rect 303418 40170 303488 40226
rect 303168 40102 303488 40170
rect 303168 40046 303238 40102
rect 303294 40046 303362 40102
rect 303418 40046 303488 40102
rect 303168 39978 303488 40046
rect 303168 39922 303238 39978
rect 303294 39922 303362 39978
rect 303418 39922 303488 39978
rect 303168 39888 303488 39922
rect 312618 40350 313238 57922
rect 312618 40294 312714 40350
rect 312770 40294 312838 40350
rect 312894 40294 312962 40350
rect 313018 40294 313086 40350
rect 313142 40294 313238 40350
rect 312618 40226 313238 40294
rect 312618 40170 312714 40226
rect 312770 40170 312838 40226
rect 312894 40170 312962 40226
rect 313018 40170 313086 40226
rect 313142 40170 313238 40226
rect 312618 40102 313238 40170
rect 312618 40046 312714 40102
rect 312770 40046 312838 40102
rect 312894 40046 312962 40102
rect 313018 40046 313086 40102
rect 313142 40046 313238 40102
rect 312618 39978 313238 40046
rect 312618 39922 312714 39978
rect 312770 39922 312838 39978
rect 312894 39922 312962 39978
rect 313018 39922 313086 39978
rect 313142 39922 313238 39978
rect 285618 28294 285714 28350
rect 285770 28294 285838 28350
rect 285894 28294 285962 28350
rect 286018 28294 286086 28350
rect 286142 28294 286238 28350
rect 285618 28226 286238 28294
rect 285618 28170 285714 28226
rect 285770 28170 285838 28226
rect 285894 28170 285962 28226
rect 286018 28170 286086 28226
rect 286142 28170 286238 28226
rect 285618 28102 286238 28170
rect 285618 28046 285714 28102
rect 285770 28046 285838 28102
rect 285894 28046 285962 28102
rect 286018 28046 286086 28102
rect 286142 28046 286238 28102
rect 285618 27978 286238 28046
rect 285618 27922 285714 27978
rect 285770 27922 285838 27978
rect 285894 27922 285962 27978
rect 286018 27922 286086 27978
rect 286142 27922 286238 27978
rect 285618 10350 286238 27922
rect 285618 10294 285714 10350
rect 285770 10294 285838 10350
rect 285894 10294 285962 10350
rect 286018 10294 286086 10350
rect 286142 10294 286238 10350
rect 285618 10226 286238 10294
rect 285618 10170 285714 10226
rect 285770 10170 285838 10226
rect 285894 10170 285962 10226
rect 286018 10170 286086 10226
rect 286142 10170 286238 10226
rect 285618 10102 286238 10170
rect 285618 10046 285714 10102
rect 285770 10046 285838 10102
rect 285894 10046 285962 10102
rect 286018 10046 286086 10102
rect 286142 10046 286238 10102
rect 285618 9978 286238 10046
rect 285618 9922 285714 9978
rect 285770 9922 285838 9978
rect 285894 9922 285962 9978
rect 286018 9922 286086 9978
rect 286142 9922 286238 9978
rect 285618 -1120 286238 9922
rect 285618 -1176 285714 -1120
rect 285770 -1176 285838 -1120
rect 285894 -1176 285962 -1120
rect 286018 -1176 286086 -1120
rect 286142 -1176 286238 -1120
rect 285618 -1244 286238 -1176
rect 285618 -1300 285714 -1244
rect 285770 -1300 285838 -1244
rect 285894 -1300 285962 -1244
rect 286018 -1300 286086 -1244
rect 286142 -1300 286238 -1244
rect 285618 -1368 286238 -1300
rect 285618 -1424 285714 -1368
rect 285770 -1424 285838 -1368
rect 285894 -1424 285962 -1368
rect 286018 -1424 286086 -1368
rect 286142 -1424 286238 -1368
rect 285618 -1492 286238 -1424
rect 285618 -1548 285714 -1492
rect 285770 -1548 285838 -1492
rect 285894 -1548 285962 -1492
rect 286018 -1548 286086 -1492
rect 286142 -1548 286238 -1492
rect 285618 -1644 286238 -1548
rect 312618 22350 313238 39922
rect 312618 22294 312714 22350
rect 312770 22294 312838 22350
rect 312894 22294 312962 22350
rect 313018 22294 313086 22350
rect 313142 22294 313238 22350
rect 312618 22226 313238 22294
rect 312618 22170 312714 22226
rect 312770 22170 312838 22226
rect 312894 22170 312962 22226
rect 313018 22170 313086 22226
rect 313142 22170 313238 22226
rect 312618 22102 313238 22170
rect 312618 22046 312714 22102
rect 312770 22046 312838 22102
rect 312894 22046 312962 22102
rect 313018 22046 313086 22102
rect 313142 22046 313238 22102
rect 312618 21978 313238 22046
rect 312618 21922 312714 21978
rect 312770 21922 312838 21978
rect 312894 21922 312962 21978
rect 313018 21922 313086 21978
rect 313142 21922 313238 21978
rect 312618 4350 313238 21922
rect 312618 4294 312714 4350
rect 312770 4294 312838 4350
rect 312894 4294 312962 4350
rect 313018 4294 313086 4350
rect 313142 4294 313238 4350
rect 312618 4226 313238 4294
rect 312618 4170 312714 4226
rect 312770 4170 312838 4226
rect 312894 4170 312962 4226
rect 313018 4170 313086 4226
rect 313142 4170 313238 4226
rect 312618 4102 313238 4170
rect 312618 4046 312714 4102
rect 312770 4046 312838 4102
rect 312894 4046 312962 4102
rect 313018 4046 313086 4102
rect 313142 4046 313238 4102
rect 312618 3978 313238 4046
rect 312618 3922 312714 3978
rect 312770 3922 312838 3978
rect 312894 3922 312962 3978
rect 313018 3922 313086 3978
rect 313142 3922 313238 3978
rect 312618 -160 313238 3922
rect 312618 -216 312714 -160
rect 312770 -216 312838 -160
rect 312894 -216 312962 -160
rect 313018 -216 313086 -160
rect 313142 -216 313238 -160
rect 312618 -284 313238 -216
rect 312618 -340 312714 -284
rect 312770 -340 312838 -284
rect 312894 -340 312962 -284
rect 313018 -340 313086 -284
rect 313142 -340 313238 -284
rect 312618 -408 313238 -340
rect 312618 -464 312714 -408
rect 312770 -464 312838 -408
rect 312894 -464 312962 -408
rect 313018 -464 313086 -408
rect 313142 -464 313238 -408
rect 312618 -532 313238 -464
rect 312618 -588 312714 -532
rect 312770 -588 312838 -532
rect 312894 -588 312962 -532
rect 313018 -588 313086 -532
rect 313142 -588 313238 -532
rect 312618 -1644 313238 -588
rect 316338 64350 316958 68098
rect 316338 64294 316434 64350
rect 316490 64294 316558 64350
rect 316614 64294 316682 64350
rect 316738 64294 316806 64350
rect 316862 64294 316958 64350
rect 316338 64226 316958 64294
rect 316338 64170 316434 64226
rect 316490 64170 316558 64226
rect 316614 64170 316682 64226
rect 316738 64170 316806 64226
rect 316862 64170 316958 64226
rect 316338 64102 316958 64170
rect 316338 64046 316434 64102
rect 316490 64046 316558 64102
rect 316614 64046 316682 64102
rect 316738 64046 316806 64102
rect 316862 64046 316958 64102
rect 316338 63978 316958 64046
rect 316338 63922 316434 63978
rect 316490 63922 316558 63978
rect 316614 63922 316682 63978
rect 316738 63922 316806 63978
rect 316862 63922 316958 63978
rect 316338 46350 316958 63922
rect 318528 64350 318848 64384
rect 318528 64294 318598 64350
rect 318654 64294 318722 64350
rect 318778 64294 318848 64350
rect 318528 64226 318848 64294
rect 318528 64170 318598 64226
rect 318654 64170 318722 64226
rect 318778 64170 318848 64226
rect 318528 64102 318848 64170
rect 318528 64046 318598 64102
rect 318654 64046 318722 64102
rect 318778 64046 318848 64102
rect 318528 63978 318848 64046
rect 318528 63922 318598 63978
rect 318654 63922 318722 63978
rect 318778 63922 318848 63978
rect 318528 63888 318848 63922
rect 340172 49476 340228 97580
rect 340284 95956 340340 95966
rect 340284 66276 340340 95900
rect 340396 86660 340452 105980
rect 340396 86594 340452 86604
rect 341852 70532 341908 120540
rect 341964 117236 342020 127260
rect 342188 119924 342244 130060
rect 343338 130102 343958 130170
rect 343338 130046 343434 130102
rect 343490 130046 343558 130102
rect 343614 130046 343682 130102
rect 343738 130046 343806 130102
rect 343862 130046 343958 130102
rect 343338 129978 343958 130046
rect 343338 129922 343434 129978
rect 343490 129922 343558 129978
rect 343614 129922 343682 129978
rect 343738 129922 343806 129978
rect 343862 129922 343958 129978
rect 342188 119858 342244 119868
rect 342636 127876 342692 127886
rect 342636 117908 342692 127820
rect 342636 117842 342692 117852
rect 341964 117170 342020 117180
rect 343338 112350 343958 129922
rect 345212 133476 345268 133486
rect 345212 122518 345268 133420
rect 345212 122452 345268 122462
rect 343338 112294 343434 112350
rect 343490 112294 343558 112350
rect 343614 112294 343682 112350
rect 343738 112294 343806 112350
rect 343862 112294 343958 112350
rect 343338 112226 343958 112294
rect 343338 112170 343434 112226
rect 343490 112170 343558 112226
rect 343614 112170 343682 112226
rect 343738 112170 343806 112226
rect 343862 112170 343958 112226
rect 343338 112102 343958 112170
rect 343338 112046 343434 112102
rect 343490 112046 343558 112102
rect 343614 112046 343682 112102
rect 343738 112046 343806 112102
rect 343862 112046 343958 112102
rect 343338 111978 343958 112046
rect 343338 111922 343434 111978
rect 343490 111922 343558 111978
rect 343614 111922 343682 111978
rect 343738 111922 343806 111978
rect 343862 111922 343958 111978
rect 341852 70466 341908 70476
rect 341964 98756 342020 98766
rect 340284 66210 340340 66220
rect 341964 52164 342020 98700
rect 341964 52098 342020 52108
rect 343338 94350 343958 111922
rect 345324 118916 345380 118926
rect 343338 94294 343434 94350
rect 343490 94294 343558 94350
rect 343614 94294 343682 94350
rect 343738 94294 343806 94350
rect 343862 94294 343958 94350
rect 343338 94226 343958 94294
rect 343338 94170 343434 94226
rect 343490 94170 343558 94226
rect 343614 94170 343682 94226
rect 343738 94170 343806 94226
rect 343862 94170 343958 94226
rect 343338 94102 343958 94170
rect 343338 94046 343434 94102
rect 343490 94046 343558 94102
rect 343614 94046 343682 94102
rect 343738 94046 343806 94102
rect 343862 94046 343958 94102
rect 343338 93978 343958 94046
rect 343338 93922 343434 93978
rect 343490 93922 343558 93978
rect 343614 93922 343682 93978
rect 343738 93922 343806 93978
rect 343862 93922 343958 93978
rect 343338 76350 343958 93922
rect 343338 76294 343434 76350
rect 343490 76294 343558 76350
rect 343614 76294 343682 76350
rect 343738 76294 343806 76350
rect 343862 76294 343958 76350
rect 343338 76226 343958 76294
rect 343338 76170 343434 76226
rect 343490 76170 343558 76226
rect 343614 76170 343682 76226
rect 343738 76170 343806 76226
rect 343862 76170 343958 76226
rect 343338 76102 343958 76170
rect 343338 76046 343434 76102
rect 343490 76046 343558 76102
rect 343614 76046 343682 76102
rect 343738 76046 343806 76102
rect 343862 76046 343958 76102
rect 343338 75978 343958 76046
rect 343338 75922 343434 75978
rect 343490 75922 343558 75978
rect 343614 75922 343682 75978
rect 343738 75922 343806 75978
rect 343862 75922 343958 75978
rect 343338 58350 343958 75922
rect 343338 58294 343434 58350
rect 343490 58294 343558 58350
rect 343614 58294 343682 58350
rect 343738 58294 343806 58350
rect 343862 58294 343958 58350
rect 343338 58226 343958 58294
rect 343338 58170 343434 58226
rect 343490 58170 343558 58226
rect 343614 58170 343682 58226
rect 343738 58170 343806 58226
rect 343862 58170 343958 58226
rect 343338 58102 343958 58170
rect 343338 58046 343434 58102
rect 343490 58046 343558 58102
rect 343614 58046 343682 58102
rect 343738 58046 343806 58102
rect 343862 58046 343958 58102
rect 343338 57978 343958 58046
rect 343338 57922 343434 57978
rect 343490 57922 343558 57978
rect 343614 57922 343682 57978
rect 343738 57922 343806 57978
rect 343862 57922 343958 57978
rect 340172 49410 340228 49420
rect 316338 46294 316434 46350
rect 316490 46294 316558 46350
rect 316614 46294 316682 46350
rect 316738 46294 316806 46350
rect 316862 46294 316958 46350
rect 316338 46226 316958 46294
rect 316338 46170 316434 46226
rect 316490 46170 316558 46226
rect 316614 46170 316682 46226
rect 316738 46170 316806 46226
rect 316862 46170 316958 46226
rect 316338 46102 316958 46170
rect 316338 46046 316434 46102
rect 316490 46046 316558 46102
rect 316614 46046 316682 46102
rect 316738 46046 316806 46102
rect 316862 46046 316958 46102
rect 316338 45978 316958 46046
rect 316338 45922 316434 45978
rect 316490 45922 316558 45978
rect 316614 45922 316682 45978
rect 316738 45922 316806 45978
rect 316862 45922 316958 45978
rect 316338 28350 316958 45922
rect 318528 46350 318848 46384
rect 318528 46294 318598 46350
rect 318654 46294 318722 46350
rect 318778 46294 318848 46350
rect 318528 46226 318848 46294
rect 318528 46170 318598 46226
rect 318654 46170 318722 46226
rect 318778 46170 318848 46226
rect 318528 46102 318848 46170
rect 318528 46046 318598 46102
rect 318654 46046 318722 46102
rect 318778 46046 318848 46102
rect 318528 45978 318848 46046
rect 318528 45922 318598 45978
rect 318654 45922 318722 45978
rect 318778 45922 318848 45978
rect 318528 45888 318848 45922
rect 316338 28294 316434 28350
rect 316490 28294 316558 28350
rect 316614 28294 316682 28350
rect 316738 28294 316806 28350
rect 316862 28294 316958 28350
rect 316338 28226 316958 28294
rect 316338 28170 316434 28226
rect 316490 28170 316558 28226
rect 316614 28170 316682 28226
rect 316738 28170 316806 28226
rect 316862 28170 316958 28226
rect 316338 28102 316958 28170
rect 316338 28046 316434 28102
rect 316490 28046 316558 28102
rect 316614 28046 316682 28102
rect 316738 28046 316806 28102
rect 316862 28046 316958 28102
rect 316338 27978 316958 28046
rect 316338 27922 316434 27978
rect 316490 27922 316558 27978
rect 316614 27922 316682 27978
rect 316738 27922 316806 27978
rect 316862 27922 316958 27978
rect 316338 10350 316958 27922
rect 316338 10294 316434 10350
rect 316490 10294 316558 10350
rect 316614 10294 316682 10350
rect 316738 10294 316806 10350
rect 316862 10294 316958 10350
rect 316338 10226 316958 10294
rect 316338 10170 316434 10226
rect 316490 10170 316558 10226
rect 316614 10170 316682 10226
rect 316738 10170 316806 10226
rect 316862 10170 316958 10226
rect 316338 10102 316958 10170
rect 316338 10046 316434 10102
rect 316490 10046 316558 10102
rect 316614 10046 316682 10102
rect 316738 10046 316806 10102
rect 316862 10046 316958 10102
rect 316338 9978 316958 10046
rect 316338 9922 316434 9978
rect 316490 9922 316558 9978
rect 316614 9922 316682 9978
rect 316738 9922 316806 9978
rect 316862 9922 316958 9978
rect 316338 -1120 316958 9922
rect 316338 -1176 316434 -1120
rect 316490 -1176 316558 -1120
rect 316614 -1176 316682 -1120
rect 316738 -1176 316806 -1120
rect 316862 -1176 316958 -1120
rect 316338 -1244 316958 -1176
rect 316338 -1300 316434 -1244
rect 316490 -1300 316558 -1244
rect 316614 -1300 316682 -1244
rect 316738 -1300 316806 -1244
rect 316862 -1300 316958 -1244
rect 316338 -1368 316958 -1300
rect 316338 -1424 316434 -1368
rect 316490 -1424 316558 -1368
rect 316614 -1424 316682 -1368
rect 316738 -1424 316806 -1368
rect 316862 -1424 316958 -1368
rect 316338 -1492 316958 -1424
rect 316338 -1548 316434 -1492
rect 316490 -1548 316558 -1492
rect 316614 -1548 316682 -1492
rect 316738 -1548 316806 -1492
rect 316862 -1548 316958 -1492
rect 316338 -1644 316958 -1548
rect 343338 40350 343958 57922
rect 345212 97076 345268 97086
rect 345212 47460 345268 97020
rect 345324 69860 345380 118860
rect 347058 118350 347678 135922
rect 371808 136350 372128 136384
rect 371808 136294 371878 136350
rect 371934 136294 372002 136350
rect 372058 136294 372128 136350
rect 371808 136226 372128 136294
rect 371808 136170 371878 136226
rect 371934 136170 372002 136226
rect 372058 136170 372128 136226
rect 371808 136102 372128 136170
rect 371808 136046 371878 136102
rect 371934 136046 372002 136102
rect 372058 136046 372128 136102
rect 371808 135978 372128 136046
rect 371808 135922 371878 135978
rect 371934 135922 372002 135978
rect 372058 135922 372128 135978
rect 371808 135888 372128 135922
rect 351932 132916 351988 132926
rect 347788 129332 347844 129342
rect 347788 120596 347844 129276
rect 351820 121716 351876 121726
rect 347788 120530 347844 120540
rect 350252 121156 350308 121166
rect 347058 118294 347154 118350
rect 347210 118294 347278 118350
rect 347334 118294 347402 118350
rect 347458 118294 347526 118350
rect 347582 118294 347678 118350
rect 347058 118226 347678 118294
rect 347058 118170 347154 118226
rect 347210 118170 347278 118226
rect 347334 118170 347402 118226
rect 347458 118170 347526 118226
rect 347582 118170 347678 118226
rect 347058 118102 347678 118170
rect 347058 118046 347154 118102
rect 347210 118046 347278 118102
rect 347334 118046 347402 118102
rect 347458 118046 347526 118102
rect 347582 118046 347678 118102
rect 347058 117978 347678 118046
rect 347058 117922 347154 117978
rect 347210 117922 347278 117978
rect 347334 117922 347402 117978
rect 347458 117922 347526 117978
rect 347582 117922 347678 117978
rect 345436 108836 345492 108846
rect 345436 89908 345492 108780
rect 345436 89842 345492 89852
rect 345548 105476 345604 105486
rect 345548 88340 345604 105420
rect 345548 88274 345604 88284
rect 347058 100350 347678 117922
rect 348684 113316 348740 113326
rect 347058 100294 347154 100350
rect 347210 100294 347278 100350
rect 347334 100294 347402 100350
rect 347458 100294 347526 100350
rect 347582 100294 347678 100350
rect 347058 100226 347678 100294
rect 347058 100170 347154 100226
rect 347210 100170 347278 100226
rect 347334 100170 347402 100226
rect 347458 100170 347526 100226
rect 347582 100170 347678 100226
rect 347058 100102 347678 100170
rect 347058 100046 347154 100102
rect 347210 100046 347278 100102
rect 347334 100046 347402 100102
rect 347458 100046 347526 100102
rect 347582 100046 347678 100102
rect 347058 99978 347678 100046
rect 347058 99922 347154 99978
rect 347210 99922 347278 99978
rect 347334 99922 347402 99978
rect 347458 99922 347526 99978
rect 347582 99922 347678 99978
rect 347058 82350 347678 99922
rect 347058 82294 347154 82350
rect 347210 82294 347278 82350
rect 347334 82294 347402 82350
rect 347458 82294 347526 82350
rect 347582 82294 347678 82350
rect 347058 82226 347678 82294
rect 347058 82170 347154 82226
rect 347210 82170 347278 82226
rect 347334 82170 347402 82226
rect 347458 82170 347526 82226
rect 347582 82170 347678 82226
rect 347058 82102 347678 82170
rect 347058 82046 347154 82102
rect 347210 82046 347278 82102
rect 347334 82046 347402 82102
rect 347458 82046 347526 82102
rect 347582 82046 347678 82102
rect 347058 81978 347678 82046
rect 347058 81922 347154 81978
rect 347210 81922 347278 81978
rect 347334 81922 347402 81978
rect 347458 81922 347526 81978
rect 347582 81922 347678 81978
rect 345324 69794 345380 69804
rect 346892 71876 346948 71886
rect 346780 67956 346836 67966
rect 346780 54180 346836 67900
rect 346780 54114 346836 54124
rect 346892 52836 346948 71820
rect 346892 52770 346948 52780
rect 347058 64350 347678 81922
rect 348572 104916 348628 104926
rect 348572 73556 348628 104860
rect 348684 84868 348740 113260
rect 348684 84802 348740 84812
rect 348572 73490 348628 73500
rect 350252 71540 350308 121100
rect 351820 114268 351876 121660
rect 351932 120898 351988 132860
rect 356448 130350 356768 130384
rect 356448 130294 356518 130350
rect 356574 130294 356642 130350
rect 356698 130294 356768 130350
rect 356448 130226 356768 130294
rect 356448 130170 356518 130226
rect 356574 130170 356642 130226
rect 356698 130170 356768 130226
rect 356448 130102 356768 130170
rect 356448 130046 356518 130102
rect 356574 130046 356642 130102
rect 356698 130046 356768 130102
rect 356448 129978 356768 130046
rect 356448 129922 356518 129978
rect 356574 129922 356642 129978
rect 356698 129922 356768 129978
rect 356448 129888 356768 129922
rect 374058 130350 374678 147922
rect 374058 130294 374154 130350
rect 374210 130294 374278 130350
rect 374334 130294 374402 130350
rect 374458 130294 374526 130350
rect 374582 130294 374678 130350
rect 374058 130226 374678 130294
rect 374058 130170 374154 130226
rect 374210 130170 374278 130226
rect 374334 130170 374402 130226
rect 374458 130170 374526 130226
rect 374582 130170 374678 130226
rect 374058 130102 374678 130170
rect 374058 130046 374154 130102
rect 374210 130046 374278 130102
rect 374334 130046 374402 130102
rect 374458 130046 374526 130102
rect 374582 130046 374678 130102
rect 374058 129978 374678 130046
rect 374058 129922 374154 129978
rect 374210 129922 374278 129978
rect 374334 129922 374402 129978
rect 374458 129922 374526 129978
rect 374582 129922 374678 129978
rect 352716 128458 352772 128468
rect 352604 128436 352716 128458
rect 352660 128402 352716 128436
rect 352716 128392 352772 128402
rect 352604 128370 352660 128380
rect 351932 120832 351988 120842
rect 352268 122836 352324 122846
rect 351820 114212 351988 114268
rect 350252 71474 350308 71484
rect 350364 109956 350420 109966
rect 350364 68068 350420 109900
rect 351148 104356 351204 104366
rect 350476 103796 350532 103806
rect 350476 79940 350532 103740
rect 351148 101668 351204 104300
rect 351148 101602 351204 101612
rect 351932 96852 351988 114212
rect 351932 96786 351988 96796
rect 350476 79874 350532 79884
rect 352268 78260 352324 122780
rect 374058 121870 374678 129922
rect 377778 208350 378398 225922
rect 396172 228116 396228 228126
rect 377778 208294 377874 208350
rect 377930 208294 377998 208350
rect 378054 208294 378122 208350
rect 378178 208294 378246 208350
rect 378302 208294 378398 208350
rect 377778 208226 378398 208294
rect 377778 208170 377874 208226
rect 377930 208170 377998 208226
rect 378054 208170 378122 208226
rect 378178 208170 378246 208226
rect 378302 208170 378398 208226
rect 377778 208102 378398 208170
rect 377778 208046 377874 208102
rect 377930 208046 377998 208102
rect 378054 208046 378122 208102
rect 378178 208046 378246 208102
rect 378302 208046 378398 208102
rect 377778 207978 378398 208046
rect 377778 207922 377874 207978
rect 377930 207922 377998 207978
rect 378054 207922 378122 207978
rect 378178 207922 378246 207978
rect 378302 207922 378398 207978
rect 377778 190350 378398 207922
rect 395836 213108 395892 213118
rect 387168 202350 387488 202384
rect 387168 202294 387238 202350
rect 387294 202294 387362 202350
rect 387418 202294 387488 202350
rect 387168 202226 387488 202294
rect 387168 202170 387238 202226
rect 387294 202170 387362 202226
rect 387418 202170 387488 202226
rect 387168 202102 387488 202170
rect 387168 202046 387238 202102
rect 387294 202046 387362 202102
rect 387418 202046 387488 202102
rect 387168 201978 387488 202046
rect 387168 201922 387238 201978
rect 387294 201922 387362 201978
rect 387418 201922 387488 201978
rect 387168 201888 387488 201922
rect 395836 196644 395892 213052
rect 396172 213108 396228 228060
rect 396172 213042 396228 213052
rect 396732 214340 396788 214350
rect 396620 212660 396676 212670
rect 396396 211316 396452 211326
rect 396396 199948 396452 211260
rect 396396 199892 396564 199948
rect 396508 199220 396564 199892
rect 396508 199154 396564 199164
rect 395836 196578 395892 196588
rect 396508 196644 396564 196654
rect 377778 190294 377874 190350
rect 377930 190294 377998 190350
rect 378054 190294 378122 190350
rect 378178 190294 378246 190350
rect 378302 190294 378398 190350
rect 377778 190226 378398 190294
rect 377778 190170 377874 190226
rect 377930 190170 377998 190226
rect 378054 190170 378122 190226
rect 378178 190170 378246 190226
rect 378302 190170 378398 190226
rect 377778 190102 378398 190170
rect 377778 190046 377874 190102
rect 377930 190046 377998 190102
rect 378054 190046 378122 190102
rect 378178 190046 378246 190102
rect 378302 190046 378398 190102
rect 377778 189978 378398 190046
rect 377778 189922 377874 189978
rect 377930 189922 377998 189978
rect 378054 189922 378122 189978
rect 378178 189922 378246 189978
rect 378302 189922 378398 189978
rect 377778 172350 378398 189922
rect 394828 196532 394884 196542
rect 394828 188938 394884 196476
rect 396508 193438 396564 196588
rect 396620 193618 396676 212604
rect 396732 195188 396788 214284
rect 400652 210980 400708 236460
rect 400652 210914 400708 210924
rect 404778 220350 405398 237922
rect 404778 220294 404874 220350
rect 404930 220294 404998 220350
rect 405054 220294 405122 220350
rect 405178 220294 405246 220350
rect 405302 220294 405398 220350
rect 404778 220226 405398 220294
rect 404778 220170 404874 220226
rect 404930 220170 404998 220226
rect 405054 220170 405122 220226
rect 405178 220170 405246 220226
rect 405302 220170 405398 220226
rect 404778 220102 405398 220170
rect 404778 220046 404874 220102
rect 404930 220046 404998 220102
rect 405054 220046 405122 220102
rect 405178 220046 405246 220102
rect 405302 220046 405398 220102
rect 404778 219978 405398 220046
rect 404778 219922 404874 219978
rect 404930 219922 404998 219978
rect 405054 219922 405122 219978
rect 405178 219922 405246 219978
rect 405302 219922 405398 219978
rect 396732 195122 396788 195132
rect 396844 210756 396900 210766
rect 396620 193562 396788 193618
rect 396508 193382 396676 193438
rect 394828 188872 394884 188882
rect 396508 193172 396564 193182
rect 396508 187318 396564 193116
rect 396620 189140 396676 193382
rect 396732 191828 396788 193562
rect 396732 191762 396788 191772
rect 396620 189074 396676 189084
rect 396844 188468 396900 210700
rect 404778 202350 405398 219922
rect 408498 244350 409118 261922
rect 410732 268436 410788 268446
rect 410732 245812 410788 268380
rect 428316 265438 428372 268802
rect 429212 267418 429268 267428
rect 429212 266338 429268 267362
rect 429212 266272 429268 266282
rect 428316 265372 428372 265382
rect 428428 263818 428484 263828
rect 428428 260398 428484 263762
rect 433808 262350 434128 262384
rect 433808 262294 433878 262350
rect 433934 262294 434002 262350
rect 434058 262294 434128 262350
rect 433808 262226 434128 262294
rect 433808 262170 433878 262226
rect 433934 262170 434002 262226
rect 434058 262170 434128 262226
rect 433808 262102 434128 262170
rect 433808 262046 433878 262102
rect 433934 262046 434002 262102
rect 434058 262046 434128 262102
rect 433808 261978 434128 262046
rect 433808 261922 433878 261978
rect 433934 261922 434002 261978
rect 434058 261922 434128 261978
rect 433808 261888 434128 261922
rect 428428 260332 428484 260342
rect 418448 256350 418768 256384
rect 418448 256294 418518 256350
rect 418574 256294 418642 256350
rect 418698 256294 418768 256350
rect 418448 256226 418768 256294
rect 418448 256170 418518 256226
rect 418574 256170 418642 256226
rect 418698 256170 418768 256226
rect 418448 256102 418768 256170
rect 418448 256046 418518 256102
rect 418574 256046 418642 256102
rect 418698 256046 418768 256102
rect 418448 255978 418768 256046
rect 418448 255922 418518 255978
rect 418574 255922 418642 255978
rect 418698 255922 418768 255978
rect 418448 255888 418768 255922
rect 435498 256350 436118 273922
rect 435498 256294 435594 256350
rect 435650 256294 435718 256350
rect 435774 256294 435842 256350
rect 435898 256294 435966 256350
rect 436022 256294 436118 256350
rect 435498 256226 436118 256294
rect 435498 256170 435594 256226
rect 435650 256170 435718 256226
rect 435774 256170 435842 256226
rect 435898 256170 435966 256226
rect 436022 256170 436118 256226
rect 435498 256102 436118 256170
rect 435498 256046 435594 256102
rect 435650 256046 435718 256102
rect 435774 256046 435842 256102
rect 435898 256046 435966 256102
rect 436022 256046 436118 256102
rect 435498 255978 436118 256046
rect 435498 255922 435594 255978
rect 435650 255922 435718 255978
rect 435774 255922 435842 255978
rect 435898 255922 435966 255978
rect 436022 255922 436118 255978
rect 410732 245746 410788 245756
rect 408498 244294 408594 244350
rect 408650 244294 408718 244350
rect 408774 244294 408842 244350
rect 408898 244294 408966 244350
rect 409022 244294 409118 244350
rect 408498 244226 409118 244294
rect 408498 244170 408594 244226
rect 408650 244170 408718 244226
rect 408774 244170 408842 244226
rect 408898 244170 408966 244226
rect 409022 244170 409118 244226
rect 408498 244102 409118 244170
rect 408498 244046 408594 244102
rect 408650 244046 408718 244102
rect 408774 244046 408842 244102
rect 408898 244046 408966 244102
rect 409022 244046 409118 244102
rect 408498 243978 409118 244046
rect 408498 243922 408594 243978
rect 408650 243922 408718 243978
rect 408774 243922 408842 243978
rect 408898 243922 408966 243978
rect 409022 243922 409118 243978
rect 408498 226350 409118 243922
rect 435498 238350 436118 255922
rect 435498 238294 435594 238350
rect 435650 238294 435718 238350
rect 435774 238294 435842 238350
rect 435898 238294 435966 238350
rect 436022 238294 436118 238350
rect 435498 238226 436118 238294
rect 435498 238170 435594 238226
rect 435650 238170 435718 238226
rect 435774 238170 435842 238226
rect 435898 238170 435966 238226
rect 436022 238170 436118 238226
rect 435498 238102 436118 238170
rect 435498 238046 435594 238102
rect 435650 238046 435718 238102
rect 435774 238046 435842 238102
rect 435898 238046 435966 238102
rect 436022 238046 436118 238102
rect 435498 237978 436118 238046
rect 435498 237922 435594 237978
rect 435650 237922 435718 237978
rect 435774 237922 435842 237978
rect 435898 237922 435966 237978
rect 436022 237922 436118 237978
rect 408498 226294 408594 226350
rect 408650 226294 408718 226350
rect 408774 226294 408842 226350
rect 408898 226294 408966 226350
rect 409022 226294 409118 226350
rect 408498 226226 409118 226294
rect 408498 226170 408594 226226
rect 408650 226170 408718 226226
rect 408774 226170 408842 226226
rect 408898 226170 408966 226226
rect 409022 226170 409118 226226
rect 408498 226102 409118 226170
rect 408498 226046 408594 226102
rect 408650 226046 408718 226102
rect 408774 226046 408842 226102
rect 408898 226046 408966 226102
rect 409022 226046 409118 226102
rect 408498 225978 409118 226046
rect 408498 225922 408594 225978
rect 408650 225922 408718 225978
rect 408774 225922 408842 225978
rect 408898 225922 408966 225978
rect 409022 225922 409118 225978
rect 404778 202294 404874 202350
rect 404930 202294 404998 202350
rect 405054 202294 405122 202350
rect 405178 202294 405246 202350
rect 405302 202294 405398 202350
rect 404778 202226 405398 202294
rect 404778 202170 404874 202226
rect 404930 202170 404998 202226
rect 405054 202170 405122 202226
rect 405178 202170 405246 202226
rect 405302 202170 405398 202226
rect 404778 202102 405398 202170
rect 404778 202046 404874 202102
rect 404930 202046 404998 202102
rect 405054 202046 405122 202102
rect 405178 202046 405246 202102
rect 405302 202046 405398 202102
rect 404778 201978 405398 202046
rect 404778 201922 404874 201978
rect 404930 201922 404998 201978
rect 405054 201922 405122 201978
rect 405178 201922 405246 201978
rect 405302 201922 405398 201978
rect 403116 198478 403172 198488
rect 401436 198298 401492 198308
rect 401436 195778 401492 198242
rect 401436 195712 401492 195722
rect 403116 194878 403172 198422
rect 403116 194812 403172 194822
rect 403228 195058 403284 195068
rect 403228 189658 403284 195002
rect 403228 189592 403284 189602
rect 396844 188402 396900 188412
rect 396508 187252 396564 187262
rect 393260 186452 393316 186462
rect 393260 186238 393316 186396
rect 393260 186172 393316 186182
rect 387168 184350 387488 184384
rect 387168 184294 387238 184350
rect 387294 184294 387362 184350
rect 387418 184294 387488 184350
rect 387168 184226 387488 184294
rect 387168 184170 387238 184226
rect 387294 184170 387362 184226
rect 387418 184170 387488 184226
rect 387168 184102 387488 184170
rect 387168 184046 387238 184102
rect 387294 184046 387362 184102
rect 387418 184046 387488 184102
rect 387168 183978 387488 184046
rect 387168 183922 387238 183978
rect 387294 183922 387362 183978
rect 387418 183922 387488 183978
rect 387168 183888 387488 183922
rect 404778 184350 405398 201922
rect 407372 219716 407428 219726
rect 407372 191156 407428 219660
rect 407372 191090 407428 191100
rect 408498 208350 409118 225922
rect 418348 229236 418404 229246
rect 418348 224420 418404 229180
rect 418348 224354 418404 224364
rect 419132 223636 419188 223646
rect 408498 208294 408594 208350
rect 408650 208294 408718 208350
rect 408774 208294 408842 208350
rect 408898 208294 408966 208350
rect 409022 208294 409118 208350
rect 408498 208226 409118 208294
rect 408498 208170 408594 208226
rect 408650 208170 408718 208226
rect 408774 208170 408842 208226
rect 408898 208170 408966 208226
rect 409022 208170 409118 208226
rect 408498 208102 409118 208170
rect 408498 208046 408594 208102
rect 408650 208046 408718 208102
rect 408774 208046 408842 208102
rect 408898 208046 408966 208102
rect 409022 208046 409118 208102
rect 408498 207978 409118 208046
rect 408498 207922 408594 207978
rect 408650 207922 408718 207978
rect 408774 207922 408842 207978
rect 408898 207922 408966 207978
rect 409022 207922 409118 207978
rect 404778 184294 404874 184350
rect 404930 184294 404998 184350
rect 405054 184294 405122 184350
rect 405178 184294 405246 184350
rect 405302 184294 405398 184350
rect 404778 184226 405398 184294
rect 404778 184170 404874 184226
rect 404930 184170 404998 184226
rect 405054 184170 405122 184226
rect 405178 184170 405246 184226
rect 405302 184170 405398 184226
rect 404778 184102 405398 184170
rect 404778 184046 404874 184102
rect 404930 184046 404998 184102
rect 405054 184046 405122 184102
rect 405178 184046 405246 184102
rect 405302 184046 405398 184102
rect 404778 183978 405398 184046
rect 404778 183922 404874 183978
rect 404930 183922 404998 183978
rect 405054 183922 405122 183978
rect 405178 183922 405246 183978
rect 405302 183922 405398 183978
rect 377778 172294 377874 172350
rect 377930 172294 377998 172350
rect 378054 172294 378122 172350
rect 378178 172294 378246 172350
rect 378302 172294 378398 172350
rect 377778 172226 378398 172294
rect 377778 172170 377874 172226
rect 377930 172170 377998 172226
rect 378054 172170 378122 172226
rect 378178 172170 378246 172226
rect 378302 172170 378398 172226
rect 377778 172102 378398 172170
rect 377778 172046 377874 172102
rect 377930 172046 377998 172102
rect 378054 172046 378122 172102
rect 378178 172046 378246 172102
rect 378302 172046 378398 172102
rect 377778 171978 378398 172046
rect 377778 171922 377874 171978
rect 377930 171922 377998 171978
rect 378054 171922 378122 171978
rect 378178 171922 378246 171978
rect 378302 171922 378398 171978
rect 377778 154350 378398 171922
rect 377778 154294 377874 154350
rect 377930 154294 377998 154350
rect 378054 154294 378122 154350
rect 378178 154294 378246 154350
rect 378302 154294 378398 154350
rect 377778 154226 378398 154294
rect 377778 154170 377874 154226
rect 377930 154170 377998 154226
rect 378054 154170 378122 154226
rect 378178 154170 378246 154226
rect 378302 154170 378398 154226
rect 377778 154102 378398 154170
rect 377778 154046 377874 154102
rect 377930 154046 377998 154102
rect 378054 154046 378122 154102
rect 378178 154046 378246 154102
rect 378302 154046 378398 154102
rect 377778 153978 378398 154046
rect 377778 153922 377874 153978
rect 377930 153922 377998 153978
rect 378054 153922 378122 153978
rect 378178 153922 378246 153978
rect 378302 153922 378398 153978
rect 377778 136350 378398 153922
rect 380492 170996 380548 171006
rect 380492 152180 380548 170940
rect 404778 166350 405398 183922
rect 404778 166294 404874 166350
rect 404930 166294 404998 166350
rect 405054 166294 405122 166350
rect 405178 166294 405246 166350
rect 405302 166294 405398 166350
rect 404778 166226 405398 166294
rect 404778 166170 404874 166226
rect 404930 166170 404998 166226
rect 405054 166170 405122 166226
rect 405178 166170 405246 166226
rect 405302 166170 405398 166226
rect 404778 166102 405398 166170
rect 404778 166046 404874 166102
rect 404930 166046 404998 166102
rect 405054 166046 405122 166102
rect 405178 166046 405246 166102
rect 405302 166046 405398 166102
rect 404778 165978 405398 166046
rect 404778 165922 404874 165978
rect 404930 165922 404998 165978
rect 405054 165922 405122 165978
rect 405178 165922 405246 165978
rect 405302 165922 405398 165978
rect 390572 160356 390628 160366
rect 380492 152114 380548 152124
rect 390460 157556 390516 157566
rect 390460 149548 390516 157500
rect 390572 157332 390628 160300
rect 390572 157266 390628 157276
rect 395612 158116 395668 158126
rect 392252 154756 392308 154766
rect 390460 149492 390628 149548
rect 390572 142660 390628 149492
rect 392252 142772 392308 154700
rect 392252 142706 392308 142716
rect 390572 142594 390628 142604
rect 377778 136294 377874 136350
rect 377930 136294 377998 136350
rect 378054 136294 378122 136350
rect 378178 136294 378246 136350
rect 378302 136294 378398 136350
rect 377778 136226 378398 136294
rect 377778 136170 377874 136226
rect 377930 136170 377998 136226
rect 378054 136170 378122 136226
rect 378178 136170 378246 136226
rect 378302 136170 378398 136226
rect 377778 136102 378398 136170
rect 377778 136046 377874 136102
rect 377930 136046 377998 136102
rect 378054 136046 378122 136102
rect 378178 136046 378246 136102
rect 378302 136046 378398 136102
rect 377778 135978 378398 136046
rect 377778 135922 377874 135978
rect 377930 135922 377998 135978
rect 378054 135922 378122 135978
rect 378178 135922 378246 135978
rect 378302 135922 378398 135978
rect 371808 118350 372128 118384
rect 371808 118294 371878 118350
rect 371934 118294 372002 118350
rect 372058 118294 372128 118350
rect 371808 118226 372128 118294
rect 371808 118170 371878 118226
rect 371934 118170 372002 118226
rect 372058 118170 372128 118226
rect 371808 118102 372128 118170
rect 371808 118046 371878 118102
rect 371934 118046 372002 118102
rect 372058 118046 372128 118102
rect 371808 117978 372128 118046
rect 371808 117922 371878 117978
rect 371934 117922 372002 117978
rect 372058 117922 372128 117978
rect 371808 117888 372128 117922
rect 377778 118350 378398 135922
rect 387168 130350 387488 130384
rect 387168 130294 387238 130350
rect 387294 130294 387362 130350
rect 387418 130294 387488 130350
rect 387168 130226 387488 130294
rect 387168 130170 387238 130226
rect 387294 130170 387362 130226
rect 387418 130170 387488 130226
rect 387168 130102 387488 130170
rect 387168 130046 387238 130102
rect 387294 130046 387362 130102
rect 387418 130046 387488 130102
rect 387168 129978 387488 130046
rect 387168 129922 387238 129978
rect 387294 129922 387362 129978
rect 387418 129922 387488 129978
rect 387168 129888 387488 129922
rect 393260 126658 393316 126682
rect 393260 126578 393316 126588
rect 393372 125524 393428 125534
rect 393372 125398 393428 125468
rect 393372 125332 393428 125342
rect 395612 119140 395668 158060
rect 395724 156996 395780 157006
rect 395724 119364 395780 156940
rect 395836 155316 395892 155326
rect 395836 132692 395892 155260
rect 396508 151396 396564 151406
rect 396508 135380 396564 151340
rect 404778 148350 405398 165922
rect 404778 148294 404874 148350
rect 404930 148294 404998 148350
rect 405054 148294 405122 148350
rect 405178 148294 405246 148350
rect 405302 148294 405398 148350
rect 404778 148226 405398 148294
rect 404778 148170 404874 148226
rect 404930 148170 404998 148226
rect 405054 148170 405122 148226
rect 405178 148170 405246 148226
rect 405302 148170 405398 148226
rect 404778 148102 405398 148170
rect 404778 148046 404874 148102
rect 404930 148046 404998 148102
rect 405054 148046 405122 148102
rect 405178 148046 405246 148102
rect 405302 148046 405398 148102
rect 404778 147978 405398 148046
rect 404778 147922 404874 147978
rect 404930 147922 404998 147978
rect 405054 147922 405122 147978
rect 405178 147922 405246 147978
rect 405302 147922 405398 147978
rect 396508 135314 396564 135324
rect 396620 143780 396676 143790
rect 395836 132626 395892 132636
rect 396620 120596 396676 143724
rect 396956 142772 397012 142782
rect 396732 142660 396788 142670
rect 396732 124068 396788 142604
rect 396732 124002 396788 124012
rect 396844 140868 396900 140878
rect 396844 122500 396900 140812
rect 396844 122434 396900 122444
rect 396620 120530 396676 120540
rect 395724 119298 395780 119308
rect 395612 119074 395668 119084
rect 396508 119252 396564 119262
rect 377778 118294 377874 118350
rect 377930 118294 377998 118350
rect 378054 118294 378122 118350
rect 378178 118294 378246 118350
rect 378302 118294 378398 118350
rect 377778 118226 378398 118294
rect 377778 118170 377874 118226
rect 377930 118170 377998 118226
rect 378054 118170 378122 118226
rect 378178 118170 378246 118226
rect 378302 118170 378398 118226
rect 377778 118102 378398 118170
rect 377778 118046 377874 118102
rect 377930 118046 377998 118102
rect 378054 118046 378122 118102
rect 378178 118046 378246 118102
rect 378302 118046 378398 118102
rect 377778 117978 378398 118046
rect 377778 117922 377874 117978
rect 377930 117922 377998 117978
rect 378054 117922 378122 117978
rect 378178 117922 378246 117978
rect 378302 117922 378398 117978
rect 356448 112350 356768 112384
rect 356448 112294 356518 112350
rect 356574 112294 356642 112350
rect 356698 112294 356768 112350
rect 356448 112226 356768 112294
rect 356448 112170 356518 112226
rect 356574 112170 356642 112226
rect 356698 112170 356768 112226
rect 356448 112102 356768 112170
rect 356448 112046 356518 112102
rect 356574 112046 356642 112102
rect 356698 112046 356768 112102
rect 356448 111978 356768 112046
rect 356448 111922 356518 111978
rect 356574 111922 356642 111978
rect 356698 111922 356768 111978
rect 356448 111888 356768 111922
rect 374058 112350 374678 115218
rect 374058 112294 374154 112350
rect 374210 112294 374278 112350
rect 374334 112294 374402 112350
rect 374458 112294 374526 112350
rect 374582 112294 374678 112350
rect 374058 112226 374678 112294
rect 374058 112170 374154 112226
rect 374210 112170 374278 112226
rect 374334 112170 374402 112226
rect 374458 112170 374526 112226
rect 374582 112170 374678 112226
rect 374058 112102 374678 112170
rect 374058 112046 374154 112102
rect 374210 112046 374278 112102
rect 374334 112046 374402 112102
rect 374458 112046 374526 112102
rect 374582 112046 374678 112102
rect 374058 111978 374678 112046
rect 374058 111922 374154 111978
rect 374210 111922 374278 111978
rect 374334 111922 374402 111978
rect 374458 111922 374526 111978
rect 374582 111922 374678 111978
rect 352268 78194 352324 78204
rect 353612 103236 353668 103246
rect 353612 71764 353668 103180
rect 368172 101892 368228 101902
rect 368172 100772 368228 101836
rect 368172 100706 368228 100716
rect 368844 101780 368900 101790
rect 368844 100772 368900 101724
rect 368844 100706 368900 100716
rect 353612 71698 353668 71708
rect 374058 94350 374678 111922
rect 374058 94294 374154 94350
rect 374210 94294 374278 94350
rect 374334 94294 374402 94350
rect 374458 94294 374526 94350
rect 374582 94294 374678 94350
rect 374058 94226 374678 94294
rect 374058 94170 374154 94226
rect 374210 94170 374278 94226
rect 374334 94170 374402 94226
rect 374458 94170 374526 94226
rect 374582 94170 374678 94226
rect 374058 94102 374678 94170
rect 374058 94046 374154 94102
rect 374210 94046 374278 94102
rect 374334 94046 374402 94102
rect 374458 94046 374526 94102
rect 374582 94046 374678 94102
rect 374058 93978 374678 94046
rect 374058 93922 374154 93978
rect 374210 93922 374278 93978
rect 374334 93922 374402 93978
rect 374458 93922 374526 93978
rect 374582 93922 374678 93978
rect 374058 76350 374678 93922
rect 374058 76294 374154 76350
rect 374210 76294 374278 76350
rect 374334 76294 374402 76350
rect 374458 76294 374526 76350
rect 374582 76294 374678 76350
rect 374058 76226 374678 76294
rect 374058 76170 374154 76226
rect 374210 76170 374278 76226
rect 374334 76170 374402 76226
rect 374458 76170 374526 76226
rect 374582 76170 374678 76226
rect 374058 76102 374678 76170
rect 374058 76046 374154 76102
rect 374210 76046 374278 76102
rect 374334 76046 374402 76102
rect 374458 76046 374526 76102
rect 374582 76046 374678 76102
rect 374058 75978 374678 76046
rect 374058 75922 374154 75978
rect 374210 75922 374278 75978
rect 374334 75922 374402 75978
rect 374458 75922 374526 75978
rect 374582 75922 374678 75978
rect 371196 70756 371252 70766
rect 371196 69188 371252 70700
rect 371196 69122 371252 69132
rect 350364 68002 350420 68012
rect 347058 64294 347154 64350
rect 347210 64294 347278 64350
rect 347334 64294 347402 64350
rect 347458 64294 347526 64350
rect 347582 64294 347678 64350
rect 347058 64226 347678 64294
rect 347058 64170 347154 64226
rect 347210 64170 347278 64226
rect 347334 64170 347402 64226
rect 347458 64170 347526 64226
rect 347582 64170 347678 64226
rect 347058 64102 347678 64170
rect 347058 64046 347154 64102
rect 347210 64046 347278 64102
rect 347334 64046 347402 64102
rect 347458 64046 347526 64102
rect 347582 64046 347678 64102
rect 347058 63978 347678 64046
rect 347058 63922 347154 63978
rect 347210 63922 347278 63978
rect 347334 63922 347402 63978
rect 347458 63922 347526 63978
rect 347582 63922 347678 63978
rect 345212 47394 345268 47404
rect 343338 40294 343434 40350
rect 343490 40294 343558 40350
rect 343614 40294 343682 40350
rect 343738 40294 343806 40350
rect 343862 40294 343958 40350
rect 343338 40226 343958 40294
rect 343338 40170 343434 40226
rect 343490 40170 343558 40226
rect 343614 40170 343682 40226
rect 343738 40170 343806 40226
rect 343862 40170 343958 40226
rect 343338 40102 343958 40170
rect 343338 40046 343434 40102
rect 343490 40046 343558 40102
rect 343614 40046 343682 40102
rect 343738 40046 343806 40102
rect 343862 40046 343958 40102
rect 343338 39978 343958 40046
rect 343338 39922 343434 39978
rect 343490 39922 343558 39978
rect 343614 39922 343682 39978
rect 343738 39922 343806 39978
rect 343862 39922 343958 39978
rect 343338 22350 343958 39922
rect 343338 22294 343434 22350
rect 343490 22294 343558 22350
rect 343614 22294 343682 22350
rect 343738 22294 343806 22350
rect 343862 22294 343958 22350
rect 343338 22226 343958 22294
rect 343338 22170 343434 22226
rect 343490 22170 343558 22226
rect 343614 22170 343682 22226
rect 343738 22170 343806 22226
rect 343862 22170 343958 22226
rect 343338 22102 343958 22170
rect 343338 22046 343434 22102
rect 343490 22046 343558 22102
rect 343614 22046 343682 22102
rect 343738 22046 343806 22102
rect 343862 22046 343958 22102
rect 343338 21978 343958 22046
rect 343338 21922 343434 21978
rect 343490 21922 343558 21978
rect 343614 21922 343682 21978
rect 343738 21922 343806 21978
rect 343862 21922 343958 21978
rect 343338 4350 343958 21922
rect 343338 4294 343434 4350
rect 343490 4294 343558 4350
rect 343614 4294 343682 4350
rect 343738 4294 343806 4350
rect 343862 4294 343958 4350
rect 343338 4226 343958 4294
rect 343338 4170 343434 4226
rect 343490 4170 343558 4226
rect 343614 4170 343682 4226
rect 343738 4170 343806 4226
rect 343862 4170 343958 4226
rect 343338 4102 343958 4170
rect 343338 4046 343434 4102
rect 343490 4046 343558 4102
rect 343614 4046 343682 4102
rect 343738 4046 343806 4102
rect 343862 4046 343958 4102
rect 343338 3978 343958 4046
rect 343338 3922 343434 3978
rect 343490 3922 343558 3978
rect 343614 3922 343682 3978
rect 343738 3922 343806 3978
rect 343862 3922 343958 3978
rect 343338 -160 343958 3922
rect 343338 -216 343434 -160
rect 343490 -216 343558 -160
rect 343614 -216 343682 -160
rect 343738 -216 343806 -160
rect 343862 -216 343958 -160
rect 343338 -284 343958 -216
rect 343338 -340 343434 -284
rect 343490 -340 343558 -284
rect 343614 -340 343682 -284
rect 343738 -340 343806 -284
rect 343862 -340 343958 -284
rect 343338 -408 343958 -340
rect 343338 -464 343434 -408
rect 343490 -464 343558 -408
rect 343614 -464 343682 -408
rect 343738 -464 343806 -408
rect 343862 -464 343958 -408
rect 343338 -532 343958 -464
rect 343338 -588 343434 -532
rect 343490 -588 343558 -532
rect 343614 -588 343682 -532
rect 343738 -588 343806 -532
rect 343862 -588 343958 -532
rect 343338 -1644 343958 -588
rect 347058 46350 347678 63922
rect 371808 64350 372128 64384
rect 371808 64294 371878 64350
rect 371934 64294 372002 64350
rect 372058 64294 372128 64350
rect 371808 64226 372128 64294
rect 371808 64170 371878 64226
rect 371934 64170 372002 64226
rect 372058 64170 372128 64226
rect 371808 64102 372128 64170
rect 371808 64046 371878 64102
rect 371934 64046 372002 64102
rect 372058 64046 372128 64102
rect 371808 63978 372128 64046
rect 371808 63922 371878 63978
rect 371934 63922 372002 63978
rect 372058 63922 372128 63978
rect 371808 63888 372128 63922
rect 356448 58350 356768 58384
rect 356448 58294 356518 58350
rect 356574 58294 356642 58350
rect 356698 58294 356768 58350
rect 356448 58226 356768 58294
rect 356448 58170 356518 58226
rect 356574 58170 356642 58226
rect 356698 58170 356768 58226
rect 356448 58102 356768 58170
rect 356448 58046 356518 58102
rect 356574 58046 356642 58102
rect 356698 58046 356768 58102
rect 356448 57978 356768 58046
rect 356448 57922 356518 57978
rect 356574 57922 356642 57978
rect 356698 57922 356768 57978
rect 356448 57888 356768 57922
rect 374058 58350 374678 75922
rect 374058 58294 374154 58350
rect 374210 58294 374278 58350
rect 374334 58294 374402 58350
rect 374458 58294 374526 58350
rect 374582 58294 374678 58350
rect 374058 58226 374678 58294
rect 374058 58170 374154 58226
rect 374210 58170 374278 58226
rect 374334 58170 374402 58226
rect 374458 58170 374526 58226
rect 374582 58170 374678 58226
rect 374058 58102 374678 58170
rect 374058 58046 374154 58102
rect 374210 58046 374278 58102
rect 374334 58046 374402 58102
rect 374458 58046 374526 58102
rect 374582 58046 374678 58102
rect 374058 57978 374678 58046
rect 374058 57922 374154 57978
rect 374210 57922 374278 57978
rect 374334 57922 374402 57978
rect 374458 57922 374526 57978
rect 374582 57922 374678 57978
rect 349356 57092 349412 57102
rect 349356 56278 349412 57036
rect 352604 56308 352660 56318
rect 352716 56278 352772 56288
rect 352660 56252 352716 56278
rect 352604 56222 352716 56252
rect 349356 56212 349412 56222
rect 352716 56212 352772 56222
rect 347058 46294 347154 46350
rect 347210 46294 347278 46350
rect 347334 46294 347402 46350
rect 347458 46294 347526 46350
rect 347582 46294 347678 46350
rect 347058 46226 347678 46294
rect 347058 46170 347154 46226
rect 347210 46170 347278 46226
rect 347334 46170 347402 46226
rect 347458 46170 347526 46226
rect 347582 46170 347678 46226
rect 347058 46102 347678 46170
rect 347058 46046 347154 46102
rect 347210 46046 347278 46102
rect 347334 46046 347402 46102
rect 347458 46046 347526 46102
rect 347582 46046 347678 46102
rect 347058 45978 347678 46046
rect 347058 45922 347154 45978
rect 347210 45922 347278 45978
rect 347334 45922 347402 45978
rect 347458 45922 347526 45978
rect 347582 45922 347678 45978
rect 347058 28350 347678 45922
rect 371808 46350 372128 46384
rect 371808 46294 371878 46350
rect 371934 46294 372002 46350
rect 372058 46294 372128 46350
rect 371808 46226 372128 46294
rect 371808 46170 371878 46226
rect 371934 46170 372002 46226
rect 372058 46170 372128 46226
rect 371808 46102 372128 46170
rect 371808 46046 371878 46102
rect 371934 46046 372002 46102
rect 372058 46046 372128 46102
rect 371808 45978 372128 46046
rect 371808 45922 371878 45978
rect 371934 45922 372002 45978
rect 372058 45922 372128 45978
rect 371808 45888 372128 45922
rect 356448 40350 356768 40384
rect 356448 40294 356518 40350
rect 356574 40294 356642 40350
rect 356698 40294 356768 40350
rect 356448 40226 356768 40294
rect 356448 40170 356518 40226
rect 356574 40170 356642 40226
rect 356698 40170 356768 40226
rect 356448 40102 356768 40170
rect 356448 40046 356518 40102
rect 356574 40046 356642 40102
rect 356698 40046 356768 40102
rect 356448 39978 356768 40046
rect 356448 39922 356518 39978
rect 356574 39922 356642 39978
rect 356698 39922 356768 39978
rect 356448 39888 356768 39922
rect 374058 40350 374678 57922
rect 374058 40294 374154 40350
rect 374210 40294 374278 40350
rect 374334 40294 374402 40350
rect 374458 40294 374526 40350
rect 374582 40294 374678 40350
rect 374058 40226 374678 40294
rect 374058 40170 374154 40226
rect 374210 40170 374278 40226
rect 374334 40170 374402 40226
rect 374458 40170 374526 40226
rect 374582 40170 374678 40226
rect 374058 40102 374678 40170
rect 374058 40046 374154 40102
rect 374210 40046 374278 40102
rect 374334 40046 374402 40102
rect 374458 40046 374526 40102
rect 374582 40046 374678 40102
rect 374058 39978 374678 40046
rect 374058 39922 374154 39978
rect 374210 39922 374278 39978
rect 374334 39922 374402 39978
rect 374458 39922 374526 39978
rect 374582 39922 374678 39978
rect 347058 28294 347154 28350
rect 347210 28294 347278 28350
rect 347334 28294 347402 28350
rect 347458 28294 347526 28350
rect 347582 28294 347678 28350
rect 347058 28226 347678 28294
rect 347058 28170 347154 28226
rect 347210 28170 347278 28226
rect 347334 28170 347402 28226
rect 347458 28170 347526 28226
rect 347582 28170 347678 28226
rect 347058 28102 347678 28170
rect 347058 28046 347154 28102
rect 347210 28046 347278 28102
rect 347334 28046 347402 28102
rect 347458 28046 347526 28102
rect 347582 28046 347678 28102
rect 347058 27978 347678 28046
rect 347058 27922 347154 27978
rect 347210 27922 347278 27978
rect 347334 27922 347402 27978
rect 347458 27922 347526 27978
rect 347582 27922 347678 27978
rect 347058 10350 347678 27922
rect 347058 10294 347154 10350
rect 347210 10294 347278 10350
rect 347334 10294 347402 10350
rect 347458 10294 347526 10350
rect 347582 10294 347678 10350
rect 347058 10226 347678 10294
rect 347058 10170 347154 10226
rect 347210 10170 347278 10226
rect 347334 10170 347402 10226
rect 347458 10170 347526 10226
rect 347582 10170 347678 10226
rect 347058 10102 347678 10170
rect 347058 10046 347154 10102
rect 347210 10046 347278 10102
rect 347334 10046 347402 10102
rect 347458 10046 347526 10102
rect 347582 10046 347678 10102
rect 347058 9978 347678 10046
rect 347058 9922 347154 9978
rect 347210 9922 347278 9978
rect 347334 9922 347402 9978
rect 347458 9922 347526 9978
rect 347582 9922 347678 9978
rect 347058 -1120 347678 9922
rect 347058 -1176 347154 -1120
rect 347210 -1176 347278 -1120
rect 347334 -1176 347402 -1120
rect 347458 -1176 347526 -1120
rect 347582 -1176 347678 -1120
rect 347058 -1244 347678 -1176
rect 347058 -1300 347154 -1244
rect 347210 -1300 347278 -1244
rect 347334 -1300 347402 -1244
rect 347458 -1300 347526 -1244
rect 347582 -1300 347678 -1244
rect 347058 -1368 347678 -1300
rect 347058 -1424 347154 -1368
rect 347210 -1424 347278 -1368
rect 347334 -1424 347402 -1368
rect 347458 -1424 347526 -1368
rect 347582 -1424 347678 -1368
rect 347058 -1492 347678 -1424
rect 347058 -1548 347154 -1492
rect 347210 -1548 347278 -1492
rect 347334 -1548 347402 -1492
rect 347458 -1548 347526 -1492
rect 347582 -1548 347678 -1492
rect 347058 -1644 347678 -1548
rect 374058 22350 374678 39922
rect 374058 22294 374154 22350
rect 374210 22294 374278 22350
rect 374334 22294 374402 22350
rect 374458 22294 374526 22350
rect 374582 22294 374678 22350
rect 374058 22226 374678 22294
rect 374058 22170 374154 22226
rect 374210 22170 374278 22226
rect 374334 22170 374402 22226
rect 374458 22170 374526 22226
rect 374582 22170 374678 22226
rect 374058 22102 374678 22170
rect 374058 22046 374154 22102
rect 374210 22046 374278 22102
rect 374334 22046 374402 22102
rect 374458 22046 374526 22102
rect 374582 22046 374678 22102
rect 374058 21978 374678 22046
rect 374058 21922 374154 21978
rect 374210 21922 374278 21978
rect 374334 21922 374402 21978
rect 374458 21922 374526 21978
rect 374582 21922 374678 21978
rect 374058 4350 374678 21922
rect 374058 4294 374154 4350
rect 374210 4294 374278 4350
rect 374334 4294 374402 4350
rect 374458 4294 374526 4350
rect 374582 4294 374678 4350
rect 374058 4226 374678 4294
rect 374058 4170 374154 4226
rect 374210 4170 374278 4226
rect 374334 4170 374402 4226
rect 374458 4170 374526 4226
rect 374582 4170 374678 4226
rect 374058 4102 374678 4170
rect 374058 4046 374154 4102
rect 374210 4046 374278 4102
rect 374334 4046 374402 4102
rect 374458 4046 374526 4102
rect 374582 4046 374678 4102
rect 374058 3978 374678 4046
rect 374058 3922 374154 3978
rect 374210 3922 374278 3978
rect 374334 3922 374402 3978
rect 374458 3922 374526 3978
rect 374582 3922 374678 3978
rect 374058 -160 374678 3922
rect 374058 -216 374154 -160
rect 374210 -216 374278 -160
rect 374334 -216 374402 -160
rect 374458 -216 374526 -160
rect 374582 -216 374678 -160
rect 374058 -284 374678 -216
rect 374058 -340 374154 -284
rect 374210 -340 374278 -284
rect 374334 -340 374402 -284
rect 374458 -340 374526 -284
rect 374582 -340 374678 -284
rect 374058 -408 374678 -340
rect 374058 -464 374154 -408
rect 374210 -464 374278 -408
rect 374334 -464 374402 -408
rect 374458 -464 374526 -408
rect 374582 -464 374678 -408
rect 374058 -532 374678 -464
rect 374058 -588 374154 -532
rect 374210 -588 374278 -532
rect 374334 -588 374402 -532
rect 374458 -588 374526 -532
rect 374582 -588 374678 -532
rect 374058 -1644 374678 -588
rect 377778 100350 378398 117922
rect 396508 117460 396564 119196
rect 396508 117394 396564 117404
rect 396956 115780 397012 142716
rect 397068 132692 397124 132702
rect 397068 117124 397124 132636
rect 400652 131338 400708 131348
rect 400652 125938 400708 131282
rect 400652 125872 400708 125882
rect 404012 131158 404068 131168
rect 404012 119252 404068 131102
rect 404012 119186 404068 119196
rect 404778 130350 405398 147922
rect 404778 130294 404874 130350
rect 404930 130294 404998 130350
rect 405054 130294 405122 130350
rect 405178 130294 405246 130350
rect 405302 130294 405398 130350
rect 404778 130226 405398 130294
rect 404778 130170 404874 130226
rect 404930 130170 404998 130226
rect 405054 130170 405122 130226
rect 405178 130170 405246 130226
rect 405302 130170 405398 130226
rect 404778 130102 405398 130170
rect 404778 130046 404874 130102
rect 404930 130046 404998 130102
rect 405054 130046 405122 130102
rect 405178 130046 405246 130102
rect 405302 130046 405398 130102
rect 404778 129978 405398 130046
rect 404778 129922 404874 129978
rect 404930 129922 404998 129978
rect 405054 129922 405122 129978
rect 405178 129922 405246 129978
rect 405302 129922 405398 129978
rect 397068 117058 397124 117068
rect 396956 115714 397012 115724
rect 387168 112350 387488 112384
rect 387168 112294 387238 112350
rect 387294 112294 387362 112350
rect 387418 112294 387488 112350
rect 387168 112226 387488 112294
rect 387168 112170 387238 112226
rect 387294 112170 387362 112226
rect 387418 112170 387488 112226
rect 387168 112102 387488 112170
rect 387168 112046 387238 112102
rect 387294 112046 387362 112102
rect 387418 112046 387488 112102
rect 387168 111978 387488 112046
rect 387168 111922 387238 111978
rect 387294 111922 387362 111978
rect 387418 111922 387488 111978
rect 387168 111888 387488 111922
rect 404778 112350 405398 129922
rect 404778 112294 404874 112350
rect 404930 112294 404998 112350
rect 405054 112294 405122 112350
rect 405178 112294 405246 112350
rect 405302 112294 405398 112350
rect 404778 112226 405398 112294
rect 404778 112170 404874 112226
rect 404930 112170 404998 112226
rect 405054 112170 405122 112226
rect 405178 112170 405246 112226
rect 405302 112170 405398 112226
rect 404778 112102 405398 112170
rect 404778 112046 404874 112102
rect 404930 112046 404998 112102
rect 405054 112046 405122 112102
rect 405178 112046 405246 112102
rect 405302 112046 405398 112102
rect 404778 111978 405398 112046
rect 404778 111922 404874 111978
rect 404930 111922 404998 111978
rect 405054 111922 405122 111978
rect 405178 111922 405246 111978
rect 405302 111922 405398 111978
rect 377778 100294 377874 100350
rect 377930 100294 377998 100350
rect 378054 100294 378122 100350
rect 378178 100294 378246 100350
rect 378302 100294 378398 100350
rect 377778 100226 378398 100294
rect 377778 100170 377874 100226
rect 377930 100170 377998 100226
rect 378054 100170 378122 100226
rect 378178 100170 378246 100226
rect 378302 100170 378398 100226
rect 377778 100102 378398 100170
rect 377778 100046 377874 100102
rect 377930 100046 377998 100102
rect 378054 100046 378122 100102
rect 378178 100046 378246 100102
rect 378302 100046 378398 100102
rect 377778 99978 378398 100046
rect 377778 99922 377874 99978
rect 377930 99922 377998 99978
rect 378054 99922 378122 99978
rect 378178 99922 378246 99978
rect 378302 99922 378398 99978
rect 377778 82350 378398 99922
rect 399196 100884 399252 100894
rect 394828 98308 394884 98318
rect 377778 82294 377874 82350
rect 377930 82294 377998 82350
rect 378054 82294 378122 82350
rect 378178 82294 378246 82350
rect 378302 82294 378398 82350
rect 377778 82226 378398 82294
rect 377778 82170 377874 82226
rect 377930 82170 377998 82226
rect 378054 82170 378122 82226
rect 378178 82170 378246 82226
rect 378302 82170 378398 82226
rect 377778 82102 378398 82170
rect 377778 82046 377874 82102
rect 377930 82046 377998 82102
rect 378054 82046 378122 82102
rect 378178 82046 378246 82102
rect 378302 82046 378398 82102
rect 377778 81978 378398 82046
rect 377778 81922 377874 81978
rect 377930 81922 377998 81978
rect 378054 81922 378122 81978
rect 378178 81922 378246 81978
rect 378302 81922 378398 81978
rect 377778 64350 378398 81922
rect 392252 95396 392308 95406
rect 392252 72212 392308 95340
rect 392252 72146 392308 72156
rect 393932 71316 393988 71326
rect 393148 70196 393204 70206
rect 393148 67956 393204 70140
rect 393148 67890 393204 67900
rect 377778 64294 377874 64350
rect 377930 64294 377998 64350
rect 378054 64294 378122 64350
rect 378178 64294 378246 64350
rect 378302 64294 378398 64350
rect 377778 64226 378398 64294
rect 377778 64170 377874 64226
rect 377930 64170 377998 64226
rect 378054 64170 378122 64226
rect 378178 64170 378246 64226
rect 378302 64170 378398 64226
rect 377778 64102 378398 64170
rect 377778 64046 377874 64102
rect 377930 64046 377998 64102
rect 378054 64046 378122 64102
rect 378178 64046 378246 64102
rect 378302 64046 378398 64102
rect 377778 63978 378398 64046
rect 377778 63922 377874 63978
rect 377930 63922 377998 63978
rect 378054 63922 378122 63978
rect 378178 63922 378246 63978
rect 378302 63922 378398 63978
rect 377778 46350 378398 63922
rect 387168 58350 387488 58384
rect 387168 58294 387238 58350
rect 387294 58294 387362 58350
rect 387418 58294 387488 58350
rect 387168 58226 387488 58294
rect 387168 58170 387238 58226
rect 387294 58170 387362 58226
rect 387418 58170 387488 58226
rect 387168 58102 387488 58170
rect 387168 58046 387238 58102
rect 387294 58046 387362 58102
rect 387418 58046 387488 58102
rect 387168 57978 387488 58046
rect 387168 57922 387238 57978
rect 387294 57922 387362 57978
rect 387418 57922 387488 57978
rect 387168 57888 387488 57922
rect 393932 53284 393988 71260
rect 393932 53218 393988 53228
rect 394828 48132 394884 98252
rect 394940 97188 394996 97198
rect 394940 50148 394996 97132
rect 395612 93716 395668 93726
rect 395052 68628 395108 68638
rect 395052 60452 395108 68572
rect 395052 60386 395108 60396
rect 395612 52052 395668 93660
rect 396956 91700 397012 91710
rect 396620 72212 396676 72222
rect 395612 51986 395668 51996
rect 396508 52052 396564 52062
rect 394940 50082 394996 50092
rect 394828 48066 394884 48076
rect 377778 46294 377874 46350
rect 377930 46294 377998 46350
rect 378054 46294 378122 46350
rect 378178 46294 378246 46350
rect 378302 46294 378398 46350
rect 377778 46226 378398 46294
rect 377778 46170 377874 46226
rect 377930 46170 377998 46226
rect 378054 46170 378122 46226
rect 378178 46170 378246 46226
rect 378302 46170 378398 46226
rect 377778 46102 378398 46170
rect 377778 46046 377874 46102
rect 377930 46046 377998 46102
rect 378054 46046 378122 46102
rect 378178 46046 378246 46102
rect 378302 46046 378398 46102
rect 377778 45978 378398 46046
rect 377778 45922 377874 45978
rect 377930 45922 377998 45978
rect 378054 45922 378122 45978
rect 378178 45922 378246 45978
rect 378302 45922 378398 45978
rect 377778 28350 378398 45922
rect 396508 44772 396564 51996
rect 396620 46116 396676 72156
rect 396732 67956 396788 67966
rect 396732 53508 396788 67900
rect 396732 53442 396788 53452
rect 396844 60452 396900 60462
rect 396620 46050 396676 46060
rect 396844 45444 396900 60396
rect 396956 54180 397012 91644
rect 398076 74676 398132 74686
rect 398076 68292 398132 74620
rect 398076 68226 398132 68236
rect 396956 54114 397012 54124
rect 399196 48132 399252 100828
rect 404778 94350 405398 111922
rect 404778 94294 404874 94350
rect 404930 94294 404998 94350
rect 405054 94294 405122 94350
rect 405178 94294 405246 94350
rect 405302 94294 405398 94350
rect 404778 94226 405398 94294
rect 404778 94170 404874 94226
rect 404930 94170 404998 94226
rect 405054 94170 405122 94226
rect 405178 94170 405246 94226
rect 405302 94170 405398 94226
rect 404778 94102 405398 94170
rect 404778 94046 404874 94102
rect 404930 94046 404998 94102
rect 405054 94046 405122 94102
rect 405178 94046 405246 94102
rect 405302 94046 405398 94102
rect 404778 93978 405398 94046
rect 404778 93922 404874 93978
rect 404930 93922 404998 93978
rect 405054 93922 405122 93978
rect 405178 93922 405246 93978
rect 405302 93922 405398 93978
rect 404778 76350 405398 93922
rect 404778 76294 404874 76350
rect 404930 76294 404998 76350
rect 405054 76294 405122 76350
rect 405178 76294 405246 76350
rect 405302 76294 405398 76350
rect 404778 76226 405398 76294
rect 404778 76170 404874 76226
rect 404930 76170 404998 76226
rect 405054 76170 405122 76226
rect 405178 76170 405246 76226
rect 405302 76170 405398 76226
rect 404778 76102 405398 76170
rect 404778 76046 404874 76102
rect 404930 76046 404998 76102
rect 405054 76046 405122 76102
rect 405178 76046 405246 76102
rect 405302 76046 405398 76102
rect 404778 75978 405398 76046
rect 404778 75922 404874 75978
rect 404930 75922 404998 75978
rect 405054 75922 405122 75978
rect 405178 75922 405246 75978
rect 405302 75922 405398 75978
rect 402332 74676 402388 74686
rect 400652 68180 400708 68190
rect 400652 54852 400708 68124
rect 400652 54786 400708 54796
rect 402332 52836 402388 74620
rect 402332 52770 402388 52780
rect 404778 58350 405398 75922
rect 404778 58294 404874 58350
rect 404930 58294 404998 58350
rect 405054 58294 405122 58350
rect 405178 58294 405246 58350
rect 405302 58294 405398 58350
rect 404778 58226 405398 58294
rect 404778 58170 404874 58226
rect 404930 58170 404998 58226
rect 405054 58170 405122 58226
rect 405178 58170 405246 58226
rect 405302 58170 405398 58226
rect 404778 58102 405398 58170
rect 404778 58046 404874 58102
rect 404930 58046 404998 58102
rect 405054 58046 405122 58102
rect 405178 58046 405246 58102
rect 405302 58046 405398 58102
rect 404778 57978 405398 58046
rect 404778 57922 404874 57978
rect 404930 57922 404998 57978
rect 405054 57922 405122 57978
rect 405178 57922 405246 57978
rect 405302 57922 405398 57978
rect 399196 48066 399252 48076
rect 396844 45378 396900 45388
rect 396508 44706 396564 44716
rect 387168 40350 387488 40384
rect 387168 40294 387238 40350
rect 387294 40294 387362 40350
rect 387418 40294 387488 40350
rect 387168 40226 387488 40294
rect 387168 40170 387238 40226
rect 387294 40170 387362 40226
rect 387418 40170 387488 40226
rect 387168 40102 387488 40170
rect 387168 40046 387238 40102
rect 387294 40046 387362 40102
rect 387418 40046 387488 40102
rect 387168 39978 387488 40046
rect 387168 39922 387238 39978
rect 387294 39922 387362 39978
rect 387418 39922 387488 39978
rect 387168 39888 387488 39922
rect 404778 40350 405398 57922
rect 404778 40294 404874 40350
rect 404930 40294 404998 40350
rect 405054 40294 405122 40350
rect 405178 40294 405246 40350
rect 405302 40294 405398 40350
rect 404778 40226 405398 40294
rect 404778 40170 404874 40226
rect 404930 40170 404998 40226
rect 405054 40170 405122 40226
rect 405178 40170 405246 40226
rect 405302 40170 405398 40226
rect 404778 40102 405398 40170
rect 404778 40046 404874 40102
rect 404930 40046 404998 40102
rect 405054 40046 405122 40102
rect 405178 40046 405246 40102
rect 405302 40046 405398 40102
rect 404778 39978 405398 40046
rect 404778 39922 404874 39978
rect 404930 39922 404998 39978
rect 405054 39922 405122 39978
rect 405178 39922 405246 39978
rect 405302 39922 405398 39978
rect 377778 28294 377874 28350
rect 377930 28294 377998 28350
rect 378054 28294 378122 28350
rect 378178 28294 378246 28350
rect 378302 28294 378398 28350
rect 377778 28226 378398 28294
rect 377778 28170 377874 28226
rect 377930 28170 377998 28226
rect 378054 28170 378122 28226
rect 378178 28170 378246 28226
rect 378302 28170 378398 28226
rect 377778 28102 378398 28170
rect 377778 28046 377874 28102
rect 377930 28046 377998 28102
rect 378054 28046 378122 28102
rect 378178 28046 378246 28102
rect 378302 28046 378398 28102
rect 377778 27978 378398 28046
rect 377778 27922 377874 27978
rect 377930 27922 377998 27978
rect 378054 27922 378122 27978
rect 378178 27922 378246 27978
rect 378302 27922 378398 27978
rect 377778 10350 378398 27922
rect 377778 10294 377874 10350
rect 377930 10294 377998 10350
rect 378054 10294 378122 10350
rect 378178 10294 378246 10350
rect 378302 10294 378398 10350
rect 377778 10226 378398 10294
rect 377778 10170 377874 10226
rect 377930 10170 377998 10226
rect 378054 10170 378122 10226
rect 378178 10170 378246 10226
rect 378302 10170 378398 10226
rect 377778 10102 378398 10170
rect 377778 10046 377874 10102
rect 377930 10046 377998 10102
rect 378054 10046 378122 10102
rect 378178 10046 378246 10102
rect 378302 10046 378398 10102
rect 377778 9978 378398 10046
rect 377778 9922 377874 9978
rect 377930 9922 377998 9978
rect 378054 9922 378122 9978
rect 378178 9922 378246 9978
rect 378302 9922 378398 9978
rect 377778 -1120 378398 9922
rect 377778 -1176 377874 -1120
rect 377930 -1176 377998 -1120
rect 378054 -1176 378122 -1120
rect 378178 -1176 378246 -1120
rect 378302 -1176 378398 -1120
rect 377778 -1244 378398 -1176
rect 377778 -1300 377874 -1244
rect 377930 -1300 377998 -1244
rect 378054 -1300 378122 -1244
rect 378178 -1300 378246 -1244
rect 378302 -1300 378398 -1244
rect 377778 -1368 378398 -1300
rect 377778 -1424 377874 -1368
rect 377930 -1424 377998 -1368
rect 378054 -1424 378122 -1368
rect 378178 -1424 378246 -1368
rect 378302 -1424 378398 -1368
rect 377778 -1492 378398 -1424
rect 377778 -1548 377874 -1492
rect 377930 -1548 377998 -1492
rect 378054 -1548 378122 -1492
rect 378178 -1548 378246 -1492
rect 378302 -1548 378398 -1492
rect 377778 -1644 378398 -1548
rect 404778 22350 405398 39922
rect 404778 22294 404874 22350
rect 404930 22294 404998 22350
rect 405054 22294 405122 22350
rect 405178 22294 405246 22350
rect 405302 22294 405398 22350
rect 404778 22226 405398 22294
rect 404778 22170 404874 22226
rect 404930 22170 404998 22226
rect 405054 22170 405122 22226
rect 405178 22170 405246 22226
rect 405302 22170 405398 22226
rect 404778 22102 405398 22170
rect 404778 22046 404874 22102
rect 404930 22046 404998 22102
rect 405054 22046 405122 22102
rect 405178 22046 405246 22102
rect 405302 22046 405398 22102
rect 404778 21978 405398 22046
rect 404778 21922 404874 21978
rect 404930 21922 404998 21978
rect 405054 21922 405122 21978
rect 405178 21922 405246 21978
rect 405302 21922 405398 21978
rect 404778 4350 405398 21922
rect 404778 4294 404874 4350
rect 404930 4294 404998 4350
rect 405054 4294 405122 4350
rect 405178 4294 405246 4350
rect 405302 4294 405398 4350
rect 404778 4226 405398 4294
rect 404778 4170 404874 4226
rect 404930 4170 404998 4226
rect 405054 4170 405122 4226
rect 405178 4170 405246 4226
rect 405302 4170 405398 4226
rect 404778 4102 405398 4170
rect 404778 4046 404874 4102
rect 404930 4046 404998 4102
rect 405054 4046 405122 4102
rect 405178 4046 405246 4102
rect 405302 4046 405398 4102
rect 404778 3978 405398 4046
rect 404778 3922 404874 3978
rect 404930 3922 404998 3978
rect 405054 3922 405122 3978
rect 405178 3922 405246 3978
rect 405302 3922 405398 3978
rect 404778 -160 405398 3922
rect 404778 -216 404874 -160
rect 404930 -216 404998 -160
rect 405054 -216 405122 -160
rect 405178 -216 405246 -160
rect 405302 -216 405398 -160
rect 404778 -284 405398 -216
rect 404778 -340 404874 -284
rect 404930 -340 404998 -284
rect 405054 -340 405122 -284
rect 405178 -340 405246 -284
rect 405302 -340 405398 -284
rect 404778 -408 405398 -340
rect 404778 -464 404874 -408
rect 404930 -464 404998 -408
rect 405054 -464 405122 -408
rect 405178 -464 405246 -408
rect 405302 -464 405398 -408
rect 404778 -532 405398 -464
rect 404778 -588 404874 -532
rect 404930 -588 404998 -532
rect 405054 -588 405122 -532
rect 405178 -588 405246 -532
rect 405302 -588 405398 -532
rect 404778 -1644 405398 -588
rect 408498 190350 409118 207922
rect 410732 214452 410788 214462
rect 410732 191828 410788 214396
rect 419132 214340 419188 223580
rect 419132 214274 419188 214284
rect 435498 220350 436118 237922
rect 435498 220294 435594 220350
rect 435650 220294 435718 220350
rect 435774 220294 435842 220350
rect 435898 220294 435966 220350
rect 436022 220294 436118 220350
rect 435498 220226 436118 220294
rect 435498 220170 435594 220226
rect 435650 220170 435718 220226
rect 435774 220170 435842 220226
rect 435898 220170 435966 220226
rect 436022 220170 436118 220226
rect 435498 220102 436118 220170
rect 435498 220046 435594 220102
rect 435650 220046 435718 220102
rect 435774 220046 435842 220102
rect 435898 220046 435966 220102
rect 436022 220046 436118 220102
rect 435498 219978 436118 220046
rect 435498 219922 435594 219978
rect 435650 219922 435718 219978
rect 435774 219922 435842 219978
rect 435898 219922 435966 219978
rect 436022 219922 436118 219978
rect 410844 211204 410900 211214
rect 410844 196532 410900 211148
rect 433808 208350 434128 208384
rect 433808 208294 433878 208350
rect 433934 208294 434002 208350
rect 434058 208294 434128 208350
rect 433808 208226 434128 208294
rect 433808 208170 433878 208226
rect 433934 208170 434002 208226
rect 434058 208170 434128 208226
rect 433808 208102 434128 208170
rect 433808 208046 433878 208102
rect 433934 208046 434002 208102
rect 434058 208046 434128 208102
rect 433808 207978 434128 208046
rect 433808 207922 433878 207978
rect 433934 207922 434002 207978
rect 434058 207922 434128 207978
rect 433808 207888 434128 207922
rect 418448 202350 418768 202384
rect 418448 202294 418518 202350
rect 418574 202294 418642 202350
rect 418698 202294 418768 202350
rect 418448 202226 418768 202294
rect 418448 202170 418518 202226
rect 418574 202170 418642 202226
rect 418698 202170 418768 202226
rect 418448 202102 418768 202170
rect 418448 202046 418518 202102
rect 418574 202046 418642 202102
rect 418698 202046 418768 202102
rect 418448 201978 418768 202046
rect 418448 201922 418518 201978
rect 418574 201922 418642 201978
rect 418698 201922 418768 201978
rect 418448 201888 418768 201922
rect 435498 202350 436118 219922
rect 435498 202294 435594 202350
rect 435650 202294 435718 202350
rect 435774 202294 435842 202350
rect 435898 202294 435966 202350
rect 436022 202294 436118 202350
rect 435498 202226 436118 202294
rect 435498 202170 435594 202226
rect 435650 202170 435718 202226
rect 435774 202170 435842 202226
rect 435898 202170 435966 202226
rect 436022 202170 436118 202226
rect 435498 202102 436118 202170
rect 435498 202046 435594 202102
rect 435650 202046 435718 202102
rect 435774 202046 435842 202102
rect 435898 202046 435966 202102
rect 436022 202046 436118 202102
rect 435498 201978 436118 202046
rect 435498 201922 435594 201978
rect 435650 201922 435718 201978
rect 435774 201922 435842 201978
rect 435898 201922 435966 201978
rect 436022 201922 436118 201978
rect 414652 199108 414708 199118
rect 414652 198298 414708 199052
rect 414652 198232 414708 198242
rect 410844 196466 410900 196476
rect 411180 195238 411236 195248
rect 411180 195122 411236 195132
rect 411292 194516 411348 194526
rect 411292 192538 411348 194460
rect 411180 192500 411236 192510
rect 411292 192472 411348 192482
rect 411180 192358 411236 192444
rect 411180 192292 411236 192302
rect 410732 191762 410788 191772
rect 408498 190294 408594 190350
rect 408650 190294 408718 190350
rect 408774 190294 408842 190350
rect 408898 190294 408966 190350
rect 409022 190294 409118 190350
rect 408498 190226 409118 190294
rect 408498 190170 408594 190226
rect 408650 190170 408718 190226
rect 408774 190170 408842 190226
rect 408898 190170 408966 190226
rect 409022 190170 409118 190226
rect 408498 190102 409118 190170
rect 408498 190046 408594 190102
rect 408650 190046 408718 190102
rect 408774 190046 408842 190102
rect 408898 190046 408966 190102
rect 409022 190046 409118 190102
rect 408498 189978 409118 190046
rect 408498 189922 408594 189978
rect 408650 189922 408718 189978
rect 408774 189922 408842 189978
rect 408898 189922 408966 189978
rect 409022 189922 409118 189978
rect 408498 172350 409118 189922
rect 433808 190350 434128 190384
rect 433808 190294 433878 190350
rect 433934 190294 434002 190350
rect 434058 190294 434128 190350
rect 433808 190226 434128 190294
rect 433808 190170 433878 190226
rect 433934 190170 434002 190226
rect 434058 190170 434128 190226
rect 433808 190102 434128 190170
rect 433808 190046 433878 190102
rect 433934 190046 434002 190102
rect 434058 190046 434128 190102
rect 433808 189978 434128 190046
rect 433808 189922 433878 189978
rect 433934 189922 434002 189978
rect 434058 189922 434128 189978
rect 433808 189888 434128 189922
rect 418448 184350 418768 184384
rect 418448 184294 418518 184350
rect 418574 184294 418642 184350
rect 418698 184294 418768 184350
rect 418448 184226 418768 184294
rect 418448 184170 418518 184226
rect 418574 184170 418642 184226
rect 418698 184170 418768 184226
rect 418448 184102 418768 184170
rect 418448 184046 418518 184102
rect 418574 184046 418642 184102
rect 418698 184046 418768 184102
rect 418448 183978 418768 184046
rect 418448 183922 418518 183978
rect 418574 183922 418642 183978
rect 418698 183922 418768 183978
rect 418448 183888 418768 183922
rect 435498 184350 436118 201922
rect 435498 184294 435594 184350
rect 435650 184294 435718 184350
rect 435774 184294 435842 184350
rect 435898 184294 435966 184350
rect 436022 184294 436118 184350
rect 435498 184226 436118 184294
rect 435498 184170 435594 184226
rect 435650 184170 435718 184226
rect 435774 184170 435842 184226
rect 435898 184170 435966 184226
rect 436022 184170 436118 184226
rect 435498 184102 436118 184170
rect 435498 184046 435594 184102
rect 435650 184046 435718 184102
rect 435774 184046 435842 184102
rect 435898 184046 435966 184102
rect 436022 184046 436118 184102
rect 435498 183978 436118 184046
rect 435498 183922 435594 183978
rect 435650 183922 435718 183978
rect 435774 183922 435842 183978
rect 435898 183922 435966 183978
rect 436022 183922 436118 183978
rect 408498 172294 408594 172350
rect 408650 172294 408718 172350
rect 408774 172294 408842 172350
rect 408898 172294 408966 172350
rect 409022 172294 409118 172350
rect 408498 172226 409118 172294
rect 408498 172170 408594 172226
rect 408650 172170 408718 172226
rect 408774 172170 408842 172226
rect 408898 172170 408966 172226
rect 409022 172170 409118 172226
rect 408498 172102 409118 172170
rect 408498 172046 408594 172102
rect 408650 172046 408718 172102
rect 408774 172046 408842 172102
rect 408898 172046 408966 172102
rect 409022 172046 409118 172102
rect 408498 171978 409118 172046
rect 408498 171922 408594 171978
rect 408650 171922 408718 171978
rect 408774 171922 408842 171978
rect 408898 171922 408966 171978
rect 409022 171922 409118 171978
rect 408498 154350 409118 171922
rect 435498 166350 436118 183922
rect 435498 166294 435594 166350
rect 435650 166294 435718 166350
rect 435774 166294 435842 166350
rect 435898 166294 435966 166350
rect 436022 166294 436118 166350
rect 435498 166226 436118 166294
rect 435498 166170 435594 166226
rect 435650 166170 435718 166226
rect 435774 166170 435842 166226
rect 435898 166170 435966 166226
rect 436022 166170 436118 166226
rect 435498 166102 436118 166170
rect 435498 166046 435594 166102
rect 435650 166046 435718 166102
rect 435774 166046 435842 166102
rect 435898 166046 435966 166102
rect 436022 166046 436118 166102
rect 435498 165978 436118 166046
rect 435498 165922 435594 165978
rect 435650 165922 435718 165978
rect 435774 165922 435842 165978
rect 435898 165922 435966 165978
rect 436022 165922 436118 165978
rect 408498 154294 408594 154350
rect 408650 154294 408718 154350
rect 408774 154294 408842 154350
rect 408898 154294 408966 154350
rect 409022 154294 409118 154350
rect 408498 154226 409118 154294
rect 408498 154170 408594 154226
rect 408650 154170 408718 154226
rect 408774 154170 408842 154226
rect 408898 154170 408966 154226
rect 409022 154170 409118 154226
rect 408498 154102 409118 154170
rect 408498 154046 408594 154102
rect 408650 154046 408718 154102
rect 408774 154046 408842 154102
rect 408898 154046 408966 154102
rect 409022 154046 409118 154102
rect 408498 153978 409118 154046
rect 408498 153922 408594 153978
rect 408650 153922 408718 153978
rect 408774 153922 408842 153978
rect 408898 153922 408966 153978
rect 409022 153922 409118 153978
rect 408498 136350 409118 153922
rect 408498 136294 408594 136350
rect 408650 136294 408718 136350
rect 408774 136294 408842 136350
rect 408898 136294 408966 136350
rect 409022 136294 409118 136350
rect 408498 136226 409118 136294
rect 408498 136170 408594 136226
rect 408650 136170 408718 136226
rect 408774 136170 408842 136226
rect 408898 136170 408966 136226
rect 409022 136170 409118 136226
rect 408498 136102 409118 136170
rect 408498 136046 408594 136102
rect 408650 136046 408718 136102
rect 408774 136046 408842 136102
rect 408898 136046 408966 136102
rect 409022 136046 409118 136102
rect 408498 135978 409118 136046
rect 408498 135922 408594 135978
rect 408650 135922 408718 135978
rect 408774 135922 408842 135978
rect 408898 135922 408966 135978
rect 409022 135922 409118 135978
rect 408498 118350 409118 135922
rect 408498 118294 408594 118350
rect 408650 118294 408718 118350
rect 408774 118294 408842 118350
rect 408898 118294 408966 118350
rect 409022 118294 409118 118350
rect 408498 118226 409118 118294
rect 408498 118170 408594 118226
rect 408650 118170 408718 118226
rect 408774 118170 408842 118226
rect 408898 118170 408966 118226
rect 409022 118170 409118 118226
rect 408498 118102 409118 118170
rect 408498 118046 408594 118102
rect 408650 118046 408718 118102
rect 408774 118046 408842 118102
rect 408898 118046 408966 118102
rect 409022 118046 409118 118102
rect 408498 117978 409118 118046
rect 408498 117922 408594 117978
rect 408650 117922 408718 117978
rect 408774 117922 408842 117978
rect 408898 117922 408966 117978
rect 409022 117922 409118 117978
rect 408498 100350 409118 117922
rect 410844 157220 410900 157230
rect 410844 116564 410900 157164
rect 435498 148350 436118 165922
rect 435498 148294 435594 148350
rect 435650 148294 435718 148350
rect 435774 148294 435842 148350
rect 435898 148294 435966 148350
rect 436022 148294 436118 148350
rect 435498 148226 436118 148294
rect 435498 148170 435594 148226
rect 435650 148170 435718 148226
rect 435774 148170 435842 148226
rect 435898 148170 435966 148226
rect 436022 148170 436118 148226
rect 435498 148102 436118 148170
rect 435498 148046 435594 148102
rect 435650 148046 435718 148102
rect 435774 148046 435842 148102
rect 435898 148046 435966 148102
rect 436022 148046 436118 148102
rect 435498 147978 436118 148046
rect 435498 147922 435594 147978
rect 435650 147922 435718 147978
rect 435774 147922 435842 147978
rect 435898 147922 435966 147978
rect 436022 147922 436118 147978
rect 433808 136350 434128 136384
rect 433808 136294 433878 136350
rect 433934 136294 434002 136350
rect 434058 136294 434128 136350
rect 433808 136226 434128 136294
rect 433808 136170 433878 136226
rect 433934 136170 434002 136226
rect 434058 136170 434128 136226
rect 433808 136102 434128 136170
rect 433808 136046 433878 136102
rect 433934 136046 434002 136102
rect 434058 136046 434128 136102
rect 433808 135978 434128 136046
rect 433808 135922 433878 135978
rect 433934 135922 434002 135978
rect 434058 135922 434128 135978
rect 433808 135888 434128 135922
rect 418448 130350 418768 130384
rect 418448 130294 418518 130350
rect 418574 130294 418642 130350
rect 418698 130294 418768 130350
rect 418448 130226 418768 130294
rect 418448 130170 418518 130226
rect 418574 130170 418642 130226
rect 418698 130170 418768 130226
rect 418448 130102 418768 130170
rect 418448 130046 418518 130102
rect 418574 130046 418642 130102
rect 418698 130046 418768 130102
rect 418448 129978 418768 130046
rect 418448 129922 418518 129978
rect 418574 129922 418642 129978
rect 418698 129922 418768 129978
rect 418448 129888 418768 129922
rect 435498 130350 436118 147922
rect 435498 130294 435594 130350
rect 435650 130294 435718 130350
rect 435774 130294 435842 130350
rect 435898 130294 435966 130350
rect 436022 130294 436118 130350
rect 435498 130226 436118 130294
rect 435498 130170 435594 130226
rect 435650 130170 435718 130226
rect 435774 130170 435842 130226
rect 435898 130170 435966 130226
rect 436022 130170 436118 130226
rect 435498 130102 436118 130170
rect 435498 130046 435594 130102
rect 435650 130046 435718 130102
rect 435774 130046 435842 130102
rect 435898 130046 435966 130102
rect 436022 130046 436118 130102
rect 435498 129978 436118 130046
rect 435498 129922 435594 129978
rect 435650 129922 435718 129978
rect 435774 129922 435842 129978
rect 435898 129922 435966 129978
rect 436022 129922 436118 129978
rect 411516 128458 411572 128468
rect 411516 126028 411572 128402
rect 411516 125972 411684 126028
rect 411628 125906 411684 125916
rect 411180 122518 411236 122528
rect 411180 121268 411236 122462
rect 411180 121202 411236 121212
rect 435498 119854 436118 129922
rect 439218 388350 439838 404498
rect 455308 403396 455364 403406
rect 449168 400350 449488 400384
rect 449168 400294 449238 400350
rect 449294 400294 449362 400350
rect 449418 400294 449488 400350
rect 449168 400226 449488 400294
rect 449168 400170 449238 400226
rect 449294 400170 449362 400226
rect 449418 400170 449488 400226
rect 449168 400102 449488 400170
rect 449168 400046 449238 400102
rect 449294 400046 449362 400102
rect 449418 400046 449488 400102
rect 449168 399978 449488 400046
rect 449168 399922 449238 399978
rect 449294 399922 449362 399978
rect 449418 399922 449488 399978
rect 449168 399888 449488 399922
rect 439218 388294 439314 388350
rect 439370 388294 439438 388350
rect 439494 388294 439562 388350
rect 439618 388294 439686 388350
rect 439742 388294 439838 388350
rect 439218 388226 439838 388294
rect 439218 388170 439314 388226
rect 439370 388170 439438 388226
rect 439494 388170 439562 388226
rect 439618 388170 439686 388226
rect 439742 388170 439838 388226
rect 439218 388102 439838 388170
rect 439218 388046 439314 388102
rect 439370 388046 439438 388102
rect 439494 388046 439562 388102
rect 439618 388046 439686 388102
rect 439742 388046 439838 388102
rect 439218 387978 439838 388046
rect 439218 387922 439314 387978
rect 439370 387922 439438 387978
rect 439494 387922 439562 387978
rect 439618 387922 439686 387978
rect 439742 387922 439838 387978
rect 439218 370350 439838 387922
rect 439218 370294 439314 370350
rect 439370 370294 439438 370350
rect 439494 370294 439562 370350
rect 439618 370294 439686 370350
rect 439742 370294 439838 370350
rect 439218 370226 439838 370294
rect 439218 370170 439314 370226
rect 439370 370170 439438 370226
rect 439494 370170 439562 370226
rect 439618 370170 439686 370226
rect 439742 370170 439838 370226
rect 439218 370102 439838 370170
rect 439218 370046 439314 370102
rect 439370 370046 439438 370102
rect 439494 370046 439562 370102
rect 439618 370046 439686 370102
rect 439742 370046 439838 370102
rect 439218 369978 439838 370046
rect 439218 369922 439314 369978
rect 439370 369922 439438 369978
rect 439494 369922 439562 369978
rect 439618 369922 439686 369978
rect 439742 369922 439838 369978
rect 439218 352350 439838 369922
rect 455308 368676 455364 403340
rect 455420 402724 455476 402734
rect 455420 380548 455476 402668
rect 455532 394678 455588 407372
rect 455532 394612 455588 394622
rect 455532 391618 455588 391628
rect 455532 390516 455588 391562
rect 455532 390450 455588 390460
rect 455420 380482 455476 380492
rect 455308 368610 455364 368620
rect 456092 365316 456148 409388
rect 457100 406756 457156 406766
rect 456988 405412 457044 405422
rect 456988 396478 457044 405356
rect 456988 396412 457044 396422
rect 457100 366436 457156 406700
rect 457212 404068 457268 404078
rect 457212 369236 457268 404012
rect 457212 369170 457268 369180
rect 457324 367556 457380 410732
rect 458892 408772 458948 408782
rect 458780 408100 458836 408110
rect 458668 406084 458724 406094
rect 458668 398998 458724 406028
rect 458668 398932 458724 398942
rect 458780 375508 458836 408044
rect 458892 397378 458948 408716
rect 458892 397312 458948 397322
rect 459004 404740 459060 404750
rect 458780 375442 458836 375452
rect 457324 367490 457380 367500
rect 457100 366370 457156 366380
rect 459004 365428 459060 404684
rect 461132 404068 461188 404078
rect 461132 403138 461188 404012
rect 461132 403072 461188 403082
rect 461132 402052 461188 402062
rect 461132 375396 461188 401996
rect 461132 375330 461188 375340
rect 464492 372036 464548 411404
rect 464492 371970 464548 371980
rect 466218 400350 466838 417922
rect 469938 424350 470558 441922
rect 469938 424294 470034 424350
rect 470090 424294 470158 424350
rect 470214 424294 470282 424350
rect 470338 424294 470406 424350
rect 470462 424294 470558 424350
rect 469938 424226 470558 424294
rect 469938 424170 470034 424226
rect 470090 424170 470158 424226
rect 470214 424170 470282 424226
rect 470338 424170 470406 424226
rect 470462 424170 470558 424226
rect 469938 424102 470558 424170
rect 469938 424046 470034 424102
rect 470090 424046 470158 424102
rect 470214 424046 470282 424102
rect 470338 424046 470406 424102
rect 470462 424046 470558 424102
rect 469938 423978 470558 424046
rect 469938 423922 470034 423978
rect 470090 423922 470158 423978
rect 470214 423922 470282 423978
rect 470338 423922 470406 423978
rect 470462 423922 470558 423978
rect 466218 400294 466314 400350
rect 466370 400294 466438 400350
rect 466494 400294 466562 400350
rect 466618 400294 466686 400350
rect 466742 400294 466838 400350
rect 466218 400226 466838 400294
rect 466218 400170 466314 400226
rect 466370 400170 466438 400226
rect 466494 400170 466562 400226
rect 466618 400170 466686 400226
rect 466742 400170 466838 400226
rect 466218 400102 466838 400170
rect 466218 400046 466314 400102
rect 466370 400046 466438 400102
rect 466494 400046 466562 400102
rect 466618 400046 466686 400102
rect 466742 400046 466838 400102
rect 466218 399978 466838 400046
rect 466218 399922 466314 399978
rect 466370 399922 466438 399978
rect 466494 399922 466562 399978
rect 466618 399922 466686 399978
rect 466742 399922 466838 399978
rect 466218 382350 466838 399922
rect 466218 382294 466314 382350
rect 466370 382294 466438 382350
rect 466494 382294 466562 382350
rect 466618 382294 466686 382350
rect 466742 382294 466838 382350
rect 466218 382226 466838 382294
rect 466218 382170 466314 382226
rect 466370 382170 466438 382226
rect 466494 382170 466562 382226
rect 466618 382170 466686 382226
rect 466742 382170 466838 382226
rect 466218 382102 466838 382170
rect 466218 382046 466314 382102
rect 466370 382046 466438 382102
rect 466494 382046 466562 382102
rect 466618 382046 466686 382102
rect 466742 382046 466838 382102
rect 466218 381978 466838 382046
rect 466218 381922 466314 381978
rect 466370 381922 466438 381978
rect 466494 381922 466562 381978
rect 466618 381922 466686 381978
rect 466742 381922 466838 381978
rect 459004 365362 459060 365372
rect 456092 365250 456148 365260
rect 439218 352294 439314 352350
rect 439370 352294 439438 352350
rect 439494 352294 439562 352350
rect 439618 352294 439686 352350
rect 439742 352294 439838 352350
rect 439218 352226 439838 352294
rect 439218 352170 439314 352226
rect 439370 352170 439438 352226
rect 439494 352170 439562 352226
rect 439618 352170 439686 352226
rect 439742 352170 439838 352226
rect 439218 352102 439838 352170
rect 439218 352046 439314 352102
rect 439370 352046 439438 352102
rect 439494 352046 439562 352102
rect 439618 352046 439686 352102
rect 439742 352046 439838 352102
rect 439218 351978 439838 352046
rect 439218 351922 439314 351978
rect 439370 351922 439438 351978
rect 439494 351922 439562 351978
rect 439618 351922 439686 351978
rect 439742 351922 439838 351978
rect 439218 334350 439838 351922
rect 466218 364350 466838 381922
rect 467852 408772 467908 408782
rect 467852 372596 467908 408716
rect 467852 372530 467908 372540
rect 469938 406350 470558 423922
rect 496938 436350 497558 453922
rect 496938 436294 497034 436350
rect 497090 436294 497158 436350
rect 497214 436294 497282 436350
rect 497338 436294 497406 436350
rect 497462 436294 497558 436350
rect 496938 436226 497558 436294
rect 496938 436170 497034 436226
rect 497090 436170 497158 436226
rect 497214 436170 497282 436226
rect 497338 436170 497406 436226
rect 497462 436170 497558 436226
rect 496938 436102 497558 436170
rect 496938 436046 497034 436102
rect 497090 436046 497158 436102
rect 497214 436046 497282 436102
rect 497338 436046 497406 436102
rect 497462 436046 497558 436102
rect 496938 435978 497558 436046
rect 496938 435922 497034 435978
rect 497090 435922 497158 435978
rect 497214 435922 497282 435978
rect 497338 435922 497406 435978
rect 497462 435922 497558 435978
rect 472108 421540 472164 421550
rect 472108 420058 472164 421484
rect 472108 419992 472164 420002
rect 480448 418350 480768 418384
rect 480448 418294 480518 418350
rect 480574 418294 480642 418350
rect 480698 418294 480768 418350
rect 480448 418226 480768 418294
rect 480448 418170 480518 418226
rect 480574 418170 480642 418226
rect 480698 418170 480768 418226
rect 480448 418102 480768 418170
rect 480448 418046 480518 418102
rect 480574 418046 480642 418102
rect 480698 418046 480768 418102
rect 480448 417978 480768 418046
rect 480448 417922 480518 417978
rect 480574 417922 480642 417978
rect 480698 417922 480768 417978
rect 480448 417888 480768 417922
rect 496938 418350 497558 435922
rect 496938 418294 497034 418350
rect 497090 418294 497158 418350
rect 497214 418294 497282 418350
rect 497338 418294 497406 418350
rect 497462 418294 497558 418350
rect 496938 418226 497558 418294
rect 496938 418170 497034 418226
rect 497090 418170 497158 418226
rect 497214 418170 497282 418226
rect 497338 418170 497406 418226
rect 497462 418170 497558 418226
rect 496938 418102 497558 418170
rect 496938 418046 497034 418102
rect 497090 418046 497158 418102
rect 497214 418046 497282 418102
rect 497338 418046 497406 418102
rect 497462 418046 497558 418102
rect 496938 417978 497558 418046
rect 496938 417922 497034 417978
rect 497090 417922 497158 417978
rect 497214 417922 497282 417978
rect 497338 417922 497406 417978
rect 497462 417922 497558 417978
rect 472108 413476 472164 413486
rect 472108 413398 472164 413420
rect 472108 413332 472164 413342
rect 472108 412138 472164 412170
rect 472108 412066 472164 412076
rect 469938 406294 470034 406350
rect 470090 406294 470158 406350
rect 470214 406294 470282 406350
rect 470338 406294 470406 406350
rect 470462 406294 470558 406350
rect 469938 406226 470558 406294
rect 469938 406170 470034 406226
rect 470090 406170 470158 406226
rect 470214 406170 470282 406226
rect 470338 406170 470406 406226
rect 470462 406170 470558 406226
rect 469938 406102 470558 406170
rect 469938 406046 470034 406102
rect 470090 406046 470158 406102
rect 470214 406046 470282 406102
rect 470338 406046 470406 406102
rect 470462 406046 470558 406102
rect 473116 410788 473172 410798
rect 469938 405978 470558 406046
rect 469938 405922 470034 405978
rect 470090 405922 470158 405978
rect 470214 405922 470282 405978
rect 470338 405922 470406 405978
rect 470462 405922 470558 405978
rect 469938 388350 470558 405922
rect 472892 406084 472948 406094
rect 472108 404758 472164 404768
rect 472108 403396 472164 404702
rect 472108 403330 472164 403340
rect 469938 388294 470034 388350
rect 470090 388294 470158 388350
rect 470214 388294 470282 388350
rect 470338 388294 470406 388350
rect 470462 388294 470558 388350
rect 469938 388226 470558 388294
rect 469938 388170 470034 388226
rect 470090 388170 470158 388226
rect 470214 388170 470282 388226
rect 470338 388170 470406 388226
rect 470462 388170 470558 388226
rect 469938 388102 470558 388170
rect 469938 388046 470034 388102
rect 470090 388046 470158 388102
rect 470214 388046 470282 388102
rect 470338 388046 470406 388102
rect 470462 388046 470558 388102
rect 469938 387978 470558 388046
rect 469938 387922 470034 387978
rect 470090 387922 470158 387978
rect 470214 387922 470282 387978
rect 470338 387922 470406 387978
rect 470462 387922 470558 387978
rect 466218 364294 466314 364350
rect 466370 364294 466438 364350
rect 466494 364294 466562 364350
rect 466618 364294 466686 364350
rect 466742 364294 466838 364350
rect 466218 364226 466838 364294
rect 466218 364170 466314 364226
rect 466370 364170 466438 364226
rect 466494 364170 466562 364226
rect 466618 364170 466686 364226
rect 466742 364170 466838 364226
rect 466218 364102 466838 364170
rect 466218 364046 466314 364102
rect 466370 364046 466438 364102
rect 466494 364046 466562 364102
rect 466618 364046 466686 364102
rect 466742 364046 466838 364102
rect 466218 363978 466838 364046
rect 466218 363922 466314 363978
rect 466370 363922 466438 363978
rect 466494 363922 466562 363978
rect 466618 363922 466686 363978
rect 466742 363922 466838 363978
rect 449168 346350 449488 346384
rect 449168 346294 449238 346350
rect 449294 346294 449362 346350
rect 449418 346294 449488 346350
rect 449168 346226 449488 346294
rect 449168 346170 449238 346226
rect 449294 346170 449362 346226
rect 449418 346170 449488 346226
rect 449168 346102 449488 346170
rect 449168 346046 449238 346102
rect 449294 346046 449362 346102
rect 449418 346046 449488 346102
rect 449168 345978 449488 346046
rect 449168 345922 449238 345978
rect 449294 345922 449362 345978
rect 449418 345922 449488 345978
rect 449168 345888 449488 345922
rect 466218 346350 466838 363922
rect 466218 346294 466314 346350
rect 466370 346294 466438 346350
rect 466494 346294 466562 346350
rect 466618 346294 466686 346350
rect 466742 346294 466838 346350
rect 466218 346226 466838 346294
rect 466218 346170 466314 346226
rect 466370 346170 466438 346226
rect 466494 346170 466562 346226
rect 466618 346170 466686 346226
rect 466742 346170 466838 346226
rect 466218 346102 466838 346170
rect 466218 346046 466314 346102
rect 466370 346046 466438 346102
rect 466494 346046 466562 346102
rect 466618 346046 466686 346102
rect 466742 346046 466838 346102
rect 466218 345978 466838 346046
rect 466218 345922 466314 345978
rect 466370 345922 466438 345978
rect 466494 345922 466562 345978
rect 466618 345922 466686 345978
rect 466742 345922 466838 345978
rect 460236 344458 460292 344468
rect 455420 340452 455476 340462
rect 455420 339778 455476 340396
rect 460236 340138 460292 344402
rect 460236 340072 460292 340082
rect 461132 341398 461188 341408
rect 455420 339712 455476 339722
rect 455532 339668 455588 339678
rect 455420 339418 455476 339428
rect 455308 337876 455364 337886
rect 455308 337798 455364 337820
rect 455308 337732 455364 337742
rect 455420 337708 455476 339362
rect 455532 338878 455588 339612
rect 455532 338812 455588 338822
rect 457772 339556 457828 339566
rect 455420 337652 455588 337708
rect 455308 337078 455364 337088
rect 455308 336868 455364 337022
rect 455308 336802 455364 336812
rect 455532 335636 455588 337652
rect 455532 335570 455588 335580
rect 455644 336538 455700 336548
rect 439218 334294 439314 334350
rect 439370 334294 439438 334350
rect 439494 334294 439562 334350
rect 439618 334294 439686 334350
rect 439742 334294 439838 334350
rect 439218 334226 439838 334294
rect 439218 334170 439314 334226
rect 439370 334170 439438 334226
rect 439494 334170 439562 334226
rect 439618 334170 439686 334226
rect 439742 334170 439838 334226
rect 439218 334102 439838 334170
rect 439218 334046 439314 334102
rect 439370 334046 439438 334102
rect 439494 334046 439562 334102
rect 439618 334046 439686 334102
rect 439742 334046 439838 334102
rect 439218 333978 439838 334046
rect 439218 333922 439314 333978
rect 439370 333922 439438 333978
rect 439494 333922 439562 333978
rect 439618 333922 439686 333978
rect 439742 333922 439838 333978
rect 439218 316350 439838 333922
rect 455308 334738 455364 334748
rect 455308 332276 455364 334682
rect 455644 333620 455700 336482
rect 455644 333554 455700 333564
rect 455308 332210 455364 332220
rect 456092 333508 456148 333518
rect 455532 331858 455588 331868
rect 455308 331268 455364 331278
rect 455308 330958 455364 331212
rect 455308 330892 455364 330902
rect 455420 329878 455476 329888
rect 455420 328692 455476 329822
rect 455532 328916 455588 331802
rect 455532 328850 455588 328860
rect 455420 328626 455476 328636
rect 449168 328350 449488 328384
rect 449168 328294 449238 328350
rect 449294 328294 449362 328350
rect 449418 328294 449488 328350
rect 449168 328226 449488 328294
rect 449168 328170 449238 328226
rect 449294 328170 449362 328226
rect 449418 328170 449488 328226
rect 449168 328102 449488 328170
rect 449168 328046 449238 328102
rect 449294 328046 449362 328102
rect 449418 328046 449488 328102
rect 449168 327978 449488 328046
rect 449168 327922 449238 327978
rect 449294 327922 449362 327978
rect 449418 327922 449488 327978
rect 449168 327888 449488 327922
rect 439218 316294 439314 316350
rect 439370 316294 439438 316350
rect 439494 316294 439562 316350
rect 439618 316294 439686 316350
rect 439742 316294 439838 316350
rect 439218 316226 439838 316294
rect 439218 316170 439314 316226
rect 439370 316170 439438 316226
rect 439494 316170 439562 316226
rect 439618 316170 439686 316226
rect 439742 316170 439838 316226
rect 439218 316102 439838 316170
rect 439218 316046 439314 316102
rect 439370 316046 439438 316102
rect 439494 316046 439562 316102
rect 439618 316046 439686 316102
rect 439742 316046 439838 316102
rect 439218 315978 439838 316046
rect 439218 315922 439314 315978
rect 439370 315922 439438 315978
rect 439494 315922 439562 315978
rect 439618 315922 439686 315978
rect 439742 315922 439838 315978
rect 439218 298350 439838 315922
rect 456092 314916 456148 333452
rect 456876 318500 456932 318510
rect 456092 314850 456148 314860
rect 456204 318388 456260 318398
rect 456204 313236 456260 318332
rect 456876 315476 456932 318444
rect 456876 315410 456932 315420
rect 456204 313170 456260 313180
rect 457772 305956 457828 339500
rect 461132 339238 461188 341342
rect 461132 339172 461188 339182
rect 461132 334964 461188 334974
rect 460236 325018 460292 325028
rect 460236 322498 460292 324962
rect 460236 322432 460292 322442
rect 461132 319078 461188 334908
rect 464492 331138 464548 331148
rect 462812 330058 462868 330068
rect 462812 325918 462868 330002
rect 462812 325852 462868 325862
rect 464492 323938 464548 331082
rect 464492 323872 464548 323882
rect 466218 328350 466838 345922
rect 466218 328294 466314 328350
rect 466370 328294 466438 328350
rect 466494 328294 466562 328350
rect 466618 328294 466686 328350
rect 466742 328294 466838 328350
rect 466218 328226 466838 328294
rect 466218 328170 466314 328226
rect 466370 328170 466438 328226
rect 466494 328170 466562 328226
rect 466618 328170 466686 328226
rect 466742 328170 466838 328226
rect 466218 328102 466838 328170
rect 466218 328046 466314 328102
rect 466370 328046 466438 328102
rect 466494 328046 466562 328102
rect 466618 328046 466686 328102
rect 466742 328046 466838 328102
rect 466218 327978 466838 328046
rect 466218 327922 466314 327978
rect 466370 327922 466438 327978
rect 466494 327922 466562 327978
rect 466618 327922 466686 327978
rect 466742 327922 466838 327978
rect 461132 319012 461188 319022
rect 457772 305890 457828 305900
rect 466218 310350 466838 327922
rect 466218 310294 466314 310350
rect 466370 310294 466438 310350
rect 466494 310294 466562 310350
rect 466618 310294 466686 310350
rect 466742 310294 466838 310350
rect 466218 310226 466838 310294
rect 466218 310170 466314 310226
rect 466370 310170 466438 310226
rect 466494 310170 466562 310226
rect 466618 310170 466686 310226
rect 466742 310170 466838 310226
rect 466218 310102 466838 310170
rect 466218 310046 466314 310102
rect 466370 310046 466438 310102
rect 466494 310046 466562 310102
rect 466618 310046 466686 310102
rect 466742 310046 466838 310102
rect 466218 309978 466838 310046
rect 466218 309922 466314 309978
rect 466370 309922 466438 309978
rect 466494 309922 466562 309978
rect 466618 309922 466686 309978
rect 466742 309922 466838 309978
rect 439218 298294 439314 298350
rect 439370 298294 439438 298350
rect 439494 298294 439562 298350
rect 439618 298294 439686 298350
rect 439742 298294 439838 298350
rect 439218 298226 439838 298294
rect 439218 298170 439314 298226
rect 439370 298170 439438 298226
rect 439494 298170 439562 298226
rect 439618 298170 439686 298226
rect 439742 298170 439838 298226
rect 439218 298102 439838 298170
rect 439218 298046 439314 298102
rect 439370 298046 439438 298102
rect 439494 298046 439562 298102
rect 439618 298046 439686 298102
rect 439742 298046 439838 298102
rect 439218 297978 439838 298046
rect 439218 297922 439314 297978
rect 439370 297922 439438 297978
rect 439494 297922 439562 297978
rect 439618 297922 439686 297978
rect 439742 297922 439838 297978
rect 439218 280350 439838 297922
rect 466218 292350 466838 309922
rect 466218 292294 466314 292350
rect 466370 292294 466438 292350
rect 466494 292294 466562 292350
rect 466618 292294 466686 292350
rect 466742 292294 466838 292350
rect 466218 292226 466838 292294
rect 466218 292170 466314 292226
rect 466370 292170 466438 292226
rect 466494 292170 466562 292226
rect 466618 292170 466686 292226
rect 466742 292170 466838 292226
rect 466218 292102 466838 292170
rect 466218 292046 466314 292102
rect 466370 292046 466438 292102
rect 466494 292046 466562 292102
rect 466618 292046 466686 292102
rect 466742 292046 466838 292102
rect 466218 291978 466838 292046
rect 466218 291922 466314 291978
rect 466370 291922 466438 291978
rect 466494 291922 466562 291978
rect 466618 291922 466686 291978
rect 466742 291922 466838 291978
rect 449372 290276 449428 290286
rect 449372 284900 449428 290220
rect 449372 284834 449428 284844
rect 464492 285796 464548 285806
rect 456988 282996 457044 283006
rect 439218 280294 439314 280350
rect 439370 280294 439438 280350
rect 439494 280294 439562 280350
rect 439618 280294 439686 280350
rect 439742 280294 439838 280350
rect 439218 280226 439838 280294
rect 439218 280170 439314 280226
rect 439370 280170 439438 280226
rect 439494 280170 439562 280226
rect 439618 280170 439686 280226
rect 439742 280170 439838 280226
rect 439218 280102 439838 280170
rect 439218 280046 439314 280102
rect 439370 280046 439438 280102
rect 439494 280046 439562 280102
rect 439618 280046 439686 280102
rect 439742 280046 439838 280102
rect 439218 279978 439838 280046
rect 439218 279922 439314 279978
rect 439370 279922 439438 279978
rect 439494 279922 439562 279978
rect 439618 279922 439686 279978
rect 439742 279922 439838 279978
rect 439218 262350 439838 279922
rect 455308 282436 455364 282446
rect 455308 277318 455364 282380
rect 456092 281876 456148 281886
rect 455420 279412 455476 279422
rect 455420 278038 455476 279356
rect 455420 277972 455476 277982
rect 455308 277262 455476 277318
rect 455308 277172 455364 277182
rect 455308 277072 455364 277082
rect 449168 274350 449488 274384
rect 449168 274294 449238 274350
rect 449294 274294 449362 274350
rect 449418 274294 449488 274350
rect 449168 274226 449488 274294
rect 449168 274170 449238 274226
rect 449294 274170 449362 274226
rect 449418 274170 449488 274226
rect 449168 274102 449488 274170
rect 449168 274046 449238 274102
rect 449294 274046 449362 274102
rect 449418 274046 449488 274102
rect 449168 273978 449488 274046
rect 449168 273922 449238 273978
rect 449294 273922 449362 273978
rect 449418 273922 449488 273978
rect 449168 273888 449488 273922
rect 455420 267148 455476 277262
rect 455532 271018 455588 271028
rect 455532 268436 455588 270962
rect 455532 268370 455588 268380
rect 439218 262294 439314 262350
rect 439370 262294 439438 262350
rect 439494 262294 439562 262350
rect 439618 262294 439686 262350
rect 439742 262294 439838 262350
rect 439218 262226 439838 262294
rect 439218 262170 439314 262226
rect 439370 262170 439438 262226
rect 439494 262170 439562 262226
rect 439618 262170 439686 262226
rect 439742 262170 439838 262226
rect 439218 262102 439838 262170
rect 439218 262046 439314 262102
rect 439370 262046 439438 262102
rect 439494 262046 439562 262102
rect 439618 262046 439686 262102
rect 439742 262046 439838 262102
rect 439218 261978 439838 262046
rect 439218 261922 439314 261978
rect 439370 261922 439438 261978
rect 439494 261922 439562 261978
rect 439618 261922 439686 261978
rect 439742 261922 439838 261978
rect 439218 244350 439838 261922
rect 455308 267092 455476 267148
rect 455308 257684 455364 267092
rect 456092 258692 456148 281820
rect 456988 265748 457044 282940
rect 458780 281652 458836 281662
rect 457772 281540 457828 281550
rect 456988 265682 457044 265692
rect 457212 269780 457268 269790
rect 457100 261716 457156 261726
rect 456092 258626 456148 258636
rect 456876 259588 456932 259598
rect 456876 258238 456932 259532
rect 456876 258172 456932 258182
rect 455308 257618 455364 257628
rect 449168 256350 449488 256384
rect 449168 256294 449238 256350
rect 449294 256294 449362 256350
rect 449418 256294 449488 256350
rect 449168 256226 449488 256294
rect 449168 256170 449238 256226
rect 449294 256170 449362 256226
rect 449418 256170 449488 256226
rect 449168 256102 449488 256170
rect 449168 256046 449238 256102
rect 449294 256046 449362 256102
rect 449418 256046 449488 256102
rect 449168 255978 449488 256046
rect 449168 255922 449238 255978
rect 449294 255922 449362 255978
rect 449418 255922 449488 255978
rect 449168 255888 449488 255922
rect 457100 253558 457156 261660
rect 457100 253492 457156 253502
rect 457212 251938 457268 269724
rect 457772 268772 457828 281484
rect 457772 268706 457828 268716
rect 458668 268772 458724 268782
rect 458668 265076 458724 268716
rect 458668 265010 458724 265020
rect 458780 261044 458836 281596
rect 464492 271348 464548 285740
rect 464492 271282 464548 271292
rect 466218 274350 466838 291922
rect 466218 274294 466314 274350
rect 466370 274294 466438 274350
rect 466494 274294 466562 274350
rect 466618 274294 466686 274350
rect 466742 274294 466838 274350
rect 466218 274226 466838 274294
rect 466218 274170 466314 274226
rect 466370 274170 466438 274226
rect 466494 274170 466562 274226
rect 466618 274170 466686 274226
rect 466742 274170 466838 274226
rect 466218 274102 466838 274170
rect 466218 274046 466314 274102
rect 466370 274046 466438 274102
rect 466494 274046 466562 274102
rect 466618 274046 466686 274102
rect 466742 274046 466838 274102
rect 466218 273978 466838 274046
rect 466218 273922 466314 273978
rect 466370 273922 466438 273978
rect 466494 273922 466562 273978
rect 466618 273922 466686 273978
rect 466742 273922 466838 273978
rect 458780 260978 458836 260988
rect 458892 269108 458948 269118
rect 457212 251872 457268 251882
rect 458892 250318 458948 269052
rect 461132 265748 461188 265758
rect 461132 255178 461188 265692
rect 464492 264628 464548 264638
rect 464492 255358 464548 264572
rect 464492 255292 464548 255302
rect 466218 256350 466838 273922
rect 469938 370350 470558 387922
rect 472892 385588 472948 406028
rect 473116 404068 473172 410732
rect 495808 406350 496128 406384
rect 495808 406294 495878 406350
rect 495934 406294 496002 406350
rect 496058 406294 496128 406350
rect 495808 406226 496128 406294
rect 495808 406170 495878 406226
rect 495934 406170 496002 406226
rect 496058 406170 496128 406226
rect 495808 406102 496128 406170
rect 495808 406046 495878 406102
rect 495934 406046 496002 406102
rect 496058 406046 496128 406102
rect 495808 405978 496128 406046
rect 495808 405922 495878 405978
rect 495934 405922 496002 405978
rect 496058 405922 496128 405978
rect 495808 405888 496128 405922
rect 473116 404002 473172 404012
rect 480448 400350 480768 400384
rect 480448 400294 480518 400350
rect 480574 400294 480642 400350
rect 480698 400294 480768 400350
rect 480448 400226 480768 400294
rect 480448 400170 480518 400226
rect 480574 400170 480642 400226
rect 480698 400170 480768 400226
rect 480448 400102 480768 400170
rect 480448 400046 480518 400102
rect 480574 400046 480642 400102
rect 480698 400046 480768 400102
rect 480448 399978 480768 400046
rect 480448 399922 480518 399978
rect 480574 399922 480642 399978
rect 480698 399922 480768 399978
rect 480448 399888 480768 399922
rect 496938 400350 497558 417922
rect 500658 460350 501278 477922
rect 517468 480004 517524 480014
rect 511168 472350 511488 472384
rect 511168 472294 511238 472350
rect 511294 472294 511362 472350
rect 511418 472294 511488 472350
rect 511168 472226 511488 472294
rect 511168 472170 511238 472226
rect 511294 472170 511362 472226
rect 511418 472170 511488 472226
rect 511168 472102 511488 472170
rect 511168 472046 511238 472102
rect 511294 472046 511362 472102
rect 511418 472046 511488 472102
rect 511168 471978 511488 472046
rect 511168 471922 511238 471978
rect 511294 471922 511362 471978
rect 511418 471922 511488 471978
rect 511168 471888 511488 471922
rect 500658 460294 500754 460350
rect 500810 460294 500878 460350
rect 500934 460294 501002 460350
rect 501058 460294 501126 460350
rect 501182 460294 501278 460350
rect 500658 460226 501278 460294
rect 500658 460170 500754 460226
rect 500810 460170 500878 460226
rect 500934 460170 501002 460226
rect 501058 460170 501126 460226
rect 501182 460170 501278 460226
rect 500658 460102 501278 460170
rect 500658 460046 500754 460102
rect 500810 460046 500878 460102
rect 500934 460046 501002 460102
rect 501058 460046 501126 460102
rect 501182 460046 501278 460102
rect 500658 459978 501278 460046
rect 500658 459922 500754 459978
rect 500810 459922 500878 459978
rect 500934 459922 501002 459978
rect 501058 459922 501126 459978
rect 501182 459922 501278 459978
rect 500658 442350 501278 459922
rect 500658 442294 500754 442350
rect 500810 442294 500878 442350
rect 500934 442294 501002 442350
rect 501058 442294 501126 442350
rect 501182 442294 501278 442350
rect 500658 442226 501278 442294
rect 500658 442170 500754 442226
rect 500810 442170 500878 442226
rect 500934 442170 501002 442226
rect 501058 442170 501126 442226
rect 501182 442170 501278 442226
rect 500658 442102 501278 442170
rect 500658 442046 500754 442102
rect 500810 442046 500878 442102
rect 500934 442046 501002 442102
rect 501058 442046 501126 442102
rect 501182 442046 501278 442102
rect 500658 441978 501278 442046
rect 500658 441922 500754 441978
rect 500810 441922 500878 441978
rect 500934 441922 501002 441978
rect 501058 441922 501126 441978
rect 501182 441922 501278 441978
rect 500658 424350 501278 441922
rect 517468 432516 517524 479948
rect 518252 459396 518308 481852
rect 518252 459330 518308 459340
rect 518476 477204 518532 477214
rect 518476 458836 518532 477148
rect 518476 458770 518532 458780
rect 519148 433076 519204 483308
rect 523292 479668 523348 479678
rect 521164 479332 521220 479342
rect 519260 476644 519316 476654
rect 519260 433636 519316 476588
rect 520940 475972 520996 475982
rect 520940 449428 520996 475916
rect 521052 473956 521108 473966
rect 521052 466138 521108 473900
rect 521052 466072 521108 466082
rect 520940 449362 520996 449372
rect 521164 446180 521220 479276
rect 521164 446114 521220 446124
rect 523292 438116 523348 479612
rect 523292 438050 523348 438060
rect 527658 472350 528278 489922
rect 527658 472294 527754 472350
rect 527810 472294 527878 472350
rect 527934 472294 528002 472350
rect 528058 472294 528126 472350
rect 528182 472294 528278 472350
rect 527658 472226 528278 472294
rect 527658 472170 527754 472226
rect 527810 472170 527878 472226
rect 527934 472170 528002 472226
rect 528058 472170 528126 472226
rect 528182 472170 528278 472226
rect 527658 472102 528278 472170
rect 527658 472046 527754 472102
rect 527810 472046 527878 472102
rect 527934 472046 528002 472102
rect 528058 472046 528126 472102
rect 528182 472046 528278 472102
rect 527658 471978 528278 472046
rect 527658 471922 527754 471978
rect 527810 471922 527878 471978
rect 527934 471922 528002 471978
rect 528058 471922 528126 471978
rect 528182 471922 528278 471978
rect 527658 454350 528278 471922
rect 527658 454294 527754 454350
rect 527810 454294 527878 454350
rect 527934 454294 528002 454350
rect 528058 454294 528126 454350
rect 528182 454294 528278 454350
rect 527658 454226 528278 454294
rect 527658 454170 527754 454226
rect 527810 454170 527878 454226
rect 527934 454170 528002 454226
rect 528058 454170 528126 454226
rect 528182 454170 528278 454226
rect 527658 454102 528278 454170
rect 527658 454046 527754 454102
rect 527810 454046 527878 454102
rect 527934 454046 528002 454102
rect 528058 454046 528126 454102
rect 528182 454046 528278 454102
rect 527658 453978 528278 454046
rect 527658 453922 527754 453978
rect 527810 453922 527878 453978
rect 527934 453922 528002 453978
rect 528058 453922 528126 453978
rect 528182 453922 528278 453978
rect 519260 433570 519316 433580
rect 527658 436350 528278 453922
rect 527658 436294 527754 436350
rect 527810 436294 527878 436350
rect 527934 436294 528002 436350
rect 528058 436294 528126 436350
rect 528182 436294 528278 436350
rect 527658 436226 528278 436294
rect 527658 436170 527754 436226
rect 527810 436170 527878 436226
rect 527934 436170 528002 436226
rect 528058 436170 528126 436226
rect 528182 436170 528278 436226
rect 527658 436102 528278 436170
rect 527658 436046 527754 436102
rect 527810 436046 527878 436102
rect 527934 436046 528002 436102
rect 528058 436046 528126 436102
rect 528182 436046 528278 436102
rect 527658 435978 528278 436046
rect 527658 435922 527754 435978
rect 527810 435922 527878 435978
rect 527934 435922 528002 435978
rect 528058 435922 528126 435978
rect 528182 435922 528278 435978
rect 519148 433010 519204 433020
rect 517468 432450 517524 432460
rect 500658 424294 500754 424350
rect 500810 424294 500878 424350
rect 500934 424294 501002 424350
rect 501058 424294 501126 424350
rect 501182 424294 501278 424350
rect 500658 424226 501278 424294
rect 500658 424170 500754 424226
rect 500810 424170 500878 424226
rect 500934 424170 501002 424226
rect 501058 424170 501126 424226
rect 501182 424170 501278 424226
rect 500658 424102 501278 424170
rect 500658 424046 500754 424102
rect 500810 424046 500878 424102
rect 500934 424046 501002 424102
rect 501058 424046 501126 424102
rect 501182 424046 501278 424102
rect 500658 423978 501278 424046
rect 500658 423922 500754 423978
rect 500810 423922 500878 423978
rect 500934 423922 501002 423978
rect 501058 423922 501126 423978
rect 501182 423922 501278 423978
rect 500658 409246 501278 423922
rect 511168 418350 511488 418384
rect 511168 418294 511238 418350
rect 511294 418294 511362 418350
rect 511418 418294 511488 418350
rect 511168 418226 511488 418294
rect 511168 418170 511238 418226
rect 511294 418170 511362 418226
rect 511418 418170 511488 418226
rect 511168 418102 511488 418170
rect 511168 418046 511238 418102
rect 511294 418046 511362 418102
rect 511418 418046 511488 418102
rect 511168 417978 511488 418046
rect 511168 417922 511238 417978
rect 511294 417922 511362 417978
rect 511418 417922 511488 417978
rect 511168 417888 511488 417922
rect 527658 418350 528278 435922
rect 527658 418294 527754 418350
rect 527810 418294 527878 418350
rect 527934 418294 528002 418350
rect 528058 418294 528126 418350
rect 528182 418294 528278 418350
rect 527658 418226 528278 418294
rect 527658 418170 527754 418226
rect 527810 418170 527878 418226
rect 527934 418170 528002 418226
rect 528058 418170 528126 418226
rect 528182 418170 528278 418226
rect 527658 418102 528278 418170
rect 527658 418046 527754 418102
rect 527810 418046 527878 418102
rect 527934 418046 528002 418102
rect 528058 418046 528126 418102
rect 528182 418046 528278 418102
rect 527658 417978 528278 418046
rect 527658 417922 527754 417978
rect 527810 417922 527878 417978
rect 527934 417922 528002 417978
rect 528058 417922 528126 417978
rect 528182 417922 528278 417978
rect 523292 415018 523348 415028
rect 518252 413578 518308 413588
rect 518252 404038 518308 413522
rect 521052 410116 521108 410126
rect 518252 403972 518308 403982
rect 519148 408100 519204 408110
rect 496938 400294 497034 400350
rect 497090 400294 497158 400350
rect 497214 400294 497282 400350
rect 497338 400294 497406 400350
rect 497462 400294 497558 400350
rect 496938 400226 497558 400294
rect 496938 400170 497034 400226
rect 497090 400170 497158 400226
rect 497214 400170 497282 400226
rect 497338 400170 497406 400226
rect 497462 400170 497558 400226
rect 496938 400102 497558 400170
rect 496938 400046 497034 400102
rect 497090 400046 497158 400102
rect 497214 400046 497282 400102
rect 497338 400046 497406 400102
rect 497462 400046 497558 400102
rect 496938 399978 497558 400046
rect 496938 399922 497034 399978
rect 497090 399922 497158 399978
rect 497214 399922 497282 399978
rect 497338 399922 497406 399978
rect 497462 399922 497558 399978
rect 495808 388389 496128 388446
rect 495808 388333 495836 388389
rect 495892 388333 495940 388389
rect 495996 388333 496044 388389
rect 496100 388333 496128 388389
rect 495808 388276 496128 388333
rect 472892 385522 472948 385532
rect 476252 385588 476308 385598
rect 476252 377076 476308 385532
rect 476252 377010 476308 377020
rect 496938 382350 497558 399922
rect 496938 382294 497034 382350
rect 497090 382294 497158 382350
rect 497214 382294 497282 382350
rect 497338 382294 497406 382350
rect 497462 382294 497558 382350
rect 496938 382226 497558 382294
rect 496938 382170 497034 382226
rect 497090 382170 497158 382226
rect 497214 382170 497282 382226
rect 497338 382170 497406 382226
rect 497462 382170 497558 382226
rect 496938 382102 497558 382170
rect 496938 382046 497034 382102
rect 497090 382046 497158 382102
rect 497214 382046 497282 382102
rect 497338 382046 497406 382102
rect 497462 382046 497558 382102
rect 496938 381978 497558 382046
rect 496938 381922 497034 381978
rect 497090 381922 497158 381978
rect 497214 381922 497282 381978
rect 497338 381922 497406 381978
rect 497462 381922 497558 381978
rect 469938 370294 470034 370350
rect 470090 370294 470158 370350
rect 470214 370294 470282 370350
rect 470338 370294 470406 370350
rect 470462 370294 470558 370350
rect 469938 370226 470558 370294
rect 469938 370170 470034 370226
rect 470090 370170 470158 370226
rect 470214 370170 470282 370226
rect 470338 370170 470406 370226
rect 470462 370170 470558 370226
rect 469938 370102 470558 370170
rect 469938 370046 470034 370102
rect 470090 370046 470158 370102
rect 470214 370046 470282 370102
rect 470338 370046 470406 370102
rect 470462 370046 470558 370102
rect 469938 369978 470558 370046
rect 469938 369922 470034 369978
rect 470090 369922 470158 369978
rect 470214 369922 470282 369978
rect 470338 369922 470406 369978
rect 470462 369922 470558 369978
rect 469938 352350 470558 369922
rect 496938 364350 497558 381922
rect 496938 364294 497034 364350
rect 497090 364294 497158 364350
rect 497214 364294 497282 364350
rect 497338 364294 497406 364350
rect 497462 364294 497558 364350
rect 496938 364226 497558 364294
rect 496938 364170 497034 364226
rect 497090 364170 497158 364226
rect 497214 364170 497282 364226
rect 497338 364170 497406 364226
rect 497462 364170 497558 364226
rect 496938 364102 497558 364170
rect 496938 364046 497034 364102
rect 497090 364046 497158 364102
rect 497214 364046 497282 364102
rect 497338 364046 497406 364102
rect 497462 364046 497558 364102
rect 496938 363978 497558 364046
rect 496938 363922 497034 363978
rect 497090 363922 497158 363978
rect 497214 363922 497282 363978
rect 497338 363922 497406 363978
rect 497462 363922 497558 363978
rect 469938 352294 470034 352350
rect 470090 352294 470158 352350
rect 470214 352294 470282 352350
rect 470338 352294 470406 352350
rect 470462 352294 470558 352350
rect 469938 352226 470558 352294
rect 469938 352170 470034 352226
rect 470090 352170 470158 352226
rect 470214 352170 470282 352226
rect 470338 352170 470406 352226
rect 470462 352170 470558 352226
rect 469938 352102 470558 352170
rect 469938 352046 470034 352102
rect 470090 352046 470158 352102
rect 470214 352046 470282 352102
rect 470338 352046 470406 352102
rect 470462 352046 470558 352102
rect 469938 351978 470558 352046
rect 469938 351922 470034 351978
rect 470090 351922 470158 351978
rect 470214 351922 470282 351978
rect 470338 351922 470406 351978
rect 470462 351922 470558 351978
rect 469938 334350 470558 351922
rect 495808 352350 496128 352384
rect 495808 352294 495878 352350
rect 495934 352294 496002 352350
rect 496058 352294 496128 352350
rect 495808 352226 496128 352294
rect 495808 352170 495878 352226
rect 495934 352170 496002 352226
rect 496058 352170 496128 352226
rect 495808 352102 496128 352170
rect 495808 352046 495878 352102
rect 495934 352046 496002 352102
rect 496058 352046 496128 352102
rect 495808 351978 496128 352046
rect 495808 351922 495878 351978
rect 495934 351922 496002 351978
rect 496058 351922 496128 351978
rect 495808 351888 496128 351922
rect 473228 349748 473284 349758
rect 473228 348598 473284 349692
rect 473228 348532 473284 348542
rect 480448 346350 480768 346384
rect 480448 346294 480518 346350
rect 480574 346294 480642 346350
rect 480698 346294 480768 346350
rect 480448 346226 480768 346294
rect 480448 346170 480518 346226
rect 480574 346170 480642 346226
rect 480698 346170 480768 346226
rect 480448 346102 480768 346170
rect 480448 346046 480518 346102
rect 480574 346046 480642 346102
rect 480698 346046 480768 346102
rect 480448 345978 480768 346046
rect 480448 345922 480518 345978
rect 480574 345922 480642 345978
rect 480698 345922 480768 345978
rect 480448 345888 480768 345922
rect 496938 346350 497558 363922
rect 496938 346294 497034 346350
rect 497090 346294 497158 346350
rect 497214 346294 497282 346350
rect 497338 346294 497406 346350
rect 497462 346294 497558 346350
rect 496938 346226 497558 346294
rect 496938 346170 497034 346226
rect 497090 346170 497158 346226
rect 497214 346170 497282 346226
rect 497338 346170 497406 346226
rect 497462 346170 497558 346226
rect 496938 346102 497558 346170
rect 496938 346046 497034 346102
rect 497090 346046 497158 346102
rect 497214 346046 497282 346102
rect 497338 346046 497406 346102
rect 497462 346046 497558 346102
rect 496938 345978 497558 346046
rect 496938 345922 497034 345978
rect 497090 345922 497158 345978
rect 497214 345922 497282 345978
rect 497338 345922 497406 345978
rect 497462 345922 497558 345978
rect 476028 341758 476084 341768
rect 473676 341684 473732 341694
rect 473676 341218 473732 341628
rect 476028 341684 476084 341702
rect 476028 341618 476084 341628
rect 473676 341152 473732 341162
rect 473228 339668 473284 339678
rect 469938 334294 470034 334350
rect 470090 334294 470158 334350
rect 470214 334294 470282 334350
rect 470338 334294 470406 334350
rect 470462 334294 470558 334350
rect 469938 334226 470558 334294
rect 469938 334170 470034 334226
rect 470090 334170 470158 334226
rect 470214 334170 470282 334226
rect 470338 334170 470406 334226
rect 470462 334170 470558 334226
rect 469938 334102 470558 334170
rect 469938 334046 470034 334102
rect 470090 334046 470158 334102
rect 470214 334046 470282 334102
rect 470338 334046 470406 334102
rect 470462 334046 470558 334102
rect 469938 333978 470558 334046
rect 469938 333922 470034 333978
rect 470090 333922 470158 333978
rect 470214 333922 470282 333978
rect 470338 333922 470406 333978
rect 470462 333922 470558 333978
rect 469938 316350 470558 333922
rect 472892 338996 472948 339006
rect 472892 318388 472948 338940
rect 473116 333620 473172 333630
rect 473116 318500 473172 333564
rect 473228 333508 473284 339612
rect 496938 338718 497558 345922
rect 500658 388350 501278 403714
rect 517244 403318 517300 403328
rect 517244 401380 517300 403262
rect 517244 401314 517300 401324
rect 517468 402052 517524 402062
rect 511168 400350 511488 400384
rect 511168 400294 511238 400350
rect 511294 400294 511362 400350
rect 511418 400294 511488 400350
rect 511168 400226 511488 400294
rect 511168 400170 511238 400226
rect 511294 400170 511362 400226
rect 511418 400170 511488 400226
rect 511168 400102 511488 400170
rect 511168 400046 511238 400102
rect 511294 400046 511362 400102
rect 511418 400046 511488 400102
rect 511168 399978 511488 400046
rect 511168 399922 511238 399978
rect 511294 399922 511362 399978
rect 511418 399922 511488 399978
rect 511168 399888 511488 399922
rect 500658 388294 500754 388350
rect 500810 388294 500878 388350
rect 500934 388294 501002 388350
rect 501058 388294 501126 388350
rect 501182 388294 501278 388350
rect 500658 388226 501278 388294
rect 500658 388170 500754 388226
rect 500810 388170 500878 388226
rect 500934 388170 501002 388226
rect 501058 388170 501126 388226
rect 501182 388170 501278 388226
rect 500658 388102 501278 388170
rect 500658 388046 500754 388102
rect 500810 388046 500878 388102
rect 500934 388046 501002 388102
rect 501058 388046 501126 388102
rect 501182 388046 501278 388102
rect 500658 387978 501278 388046
rect 500658 387922 500754 387978
rect 500810 387922 500878 387978
rect 500934 387922 501002 387978
rect 501058 387922 501126 387978
rect 501182 387922 501278 387978
rect 500658 370350 501278 387922
rect 503132 385812 503188 385822
rect 503132 371476 503188 385756
rect 517468 373716 517524 401996
rect 519148 376516 519204 408044
rect 519148 376450 519204 376460
rect 519932 405300 519988 405310
rect 519932 375956 519988 405244
rect 520940 402724 520996 402734
rect 520940 385812 520996 402668
rect 520940 385746 520996 385756
rect 521052 385588 521108 410060
rect 523292 403138 523348 414962
rect 523292 403072 523348 403082
rect 521052 385522 521108 385532
rect 527658 400350 528278 417922
rect 531378 598172 531998 598268
rect 531378 598116 531474 598172
rect 531530 598116 531598 598172
rect 531654 598116 531722 598172
rect 531778 598116 531846 598172
rect 531902 598116 531998 598172
rect 531378 598048 531998 598116
rect 531378 597992 531474 598048
rect 531530 597992 531598 598048
rect 531654 597992 531722 598048
rect 531778 597992 531846 598048
rect 531902 597992 531998 598048
rect 531378 597924 531998 597992
rect 531378 597868 531474 597924
rect 531530 597868 531598 597924
rect 531654 597868 531722 597924
rect 531778 597868 531846 597924
rect 531902 597868 531998 597924
rect 531378 597800 531998 597868
rect 531378 597744 531474 597800
rect 531530 597744 531598 597800
rect 531654 597744 531722 597800
rect 531778 597744 531846 597800
rect 531902 597744 531998 597800
rect 531378 586350 531998 597744
rect 531378 586294 531474 586350
rect 531530 586294 531598 586350
rect 531654 586294 531722 586350
rect 531778 586294 531846 586350
rect 531902 586294 531998 586350
rect 531378 586226 531998 586294
rect 531378 586170 531474 586226
rect 531530 586170 531598 586226
rect 531654 586170 531722 586226
rect 531778 586170 531846 586226
rect 531902 586170 531998 586226
rect 531378 586102 531998 586170
rect 531378 586046 531474 586102
rect 531530 586046 531598 586102
rect 531654 586046 531722 586102
rect 531778 586046 531846 586102
rect 531902 586046 531998 586102
rect 531378 585978 531998 586046
rect 531378 585922 531474 585978
rect 531530 585922 531598 585978
rect 531654 585922 531722 585978
rect 531778 585922 531846 585978
rect 531902 585922 531998 585978
rect 531378 568350 531998 585922
rect 531378 568294 531474 568350
rect 531530 568294 531598 568350
rect 531654 568294 531722 568350
rect 531778 568294 531846 568350
rect 531902 568294 531998 568350
rect 531378 568226 531998 568294
rect 531378 568170 531474 568226
rect 531530 568170 531598 568226
rect 531654 568170 531722 568226
rect 531778 568170 531846 568226
rect 531902 568170 531998 568226
rect 531378 568102 531998 568170
rect 531378 568046 531474 568102
rect 531530 568046 531598 568102
rect 531654 568046 531722 568102
rect 531778 568046 531846 568102
rect 531902 568046 531998 568102
rect 531378 567978 531998 568046
rect 531378 567922 531474 567978
rect 531530 567922 531598 567978
rect 531654 567922 531722 567978
rect 531778 567922 531846 567978
rect 531902 567922 531998 567978
rect 531378 550350 531998 567922
rect 558378 597212 558998 598268
rect 558378 597156 558474 597212
rect 558530 597156 558598 597212
rect 558654 597156 558722 597212
rect 558778 597156 558846 597212
rect 558902 597156 558998 597212
rect 558378 597088 558998 597156
rect 558378 597032 558474 597088
rect 558530 597032 558598 597088
rect 558654 597032 558722 597088
rect 558778 597032 558846 597088
rect 558902 597032 558998 597088
rect 558378 596964 558998 597032
rect 558378 596908 558474 596964
rect 558530 596908 558598 596964
rect 558654 596908 558722 596964
rect 558778 596908 558846 596964
rect 558902 596908 558998 596964
rect 558378 596840 558998 596908
rect 558378 596784 558474 596840
rect 558530 596784 558598 596840
rect 558654 596784 558722 596840
rect 558778 596784 558846 596840
rect 558902 596784 558998 596840
rect 558378 580350 558998 596784
rect 558378 580294 558474 580350
rect 558530 580294 558598 580350
rect 558654 580294 558722 580350
rect 558778 580294 558846 580350
rect 558902 580294 558998 580350
rect 558378 580226 558998 580294
rect 558378 580170 558474 580226
rect 558530 580170 558598 580226
rect 558654 580170 558722 580226
rect 558778 580170 558846 580226
rect 558902 580170 558998 580226
rect 558378 580102 558998 580170
rect 558378 580046 558474 580102
rect 558530 580046 558598 580102
rect 558654 580046 558722 580102
rect 558778 580046 558846 580102
rect 558902 580046 558998 580102
rect 558378 579978 558998 580046
rect 558378 579922 558474 579978
rect 558530 579922 558598 579978
rect 558654 579922 558722 579978
rect 558778 579922 558846 579978
rect 558902 579922 558998 579978
rect 542448 562350 542768 562384
rect 542448 562294 542518 562350
rect 542574 562294 542642 562350
rect 542698 562294 542768 562350
rect 542448 562226 542768 562294
rect 542448 562170 542518 562226
rect 542574 562170 542642 562226
rect 542698 562170 542768 562226
rect 542448 562102 542768 562170
rect 542448 562046 542518 562102
rect 542574 562046 542642 562102
rect 542698 562046 542768 562102
rect 542448 561978 542768 562046
rect 542448 561922 542518 561978
rect 542574 561922 542642 561978
rect 542698 561922 542768 561978
rect 542448 561888 542768 561922
rect 558378 562350 558998 579922
rect 558378 562294 558474 562350
rect 558530 562294 558598 562350
rect 558654 562294 558722 562350
rect 558778 562294 558846 562350
rect 558902 562294 558998 562350
rect 558378 562226 558998 562294
rect 558378 562170 558474 562226
rect 558530 562170 558598 562226
rect 558654 562170 558722 562226
rect 558778 562170 558846 562226
rect 558902 562170 558998 562226
rect 558378 562102 558998 562170
rect 558378 562046 558474 562102
rect 558530 562046 558598 562102
rect 558654 562046 558722 562102
rect 558778 562046 558846 562102
rect 558902 562046 558998 562102
rect 558378 561978 558998 562046
rect 558378 561922 558474 561978
rect 558530 561922 558598 561978
rect 558654 561922 558722 561978
rect 558778 561922 558846 561978
rect 558902 561922 558998 561978
rect 535500 552580 535556 552590
rect 531378 550294 531474 550350
rect 531530 550294 531598 550350
rect 531654 550294 531722 550350
rect 531778 550294 531846 550350
rect 531902 550294 531998 550350
rect 531378 550226 531998 550294
rect 531378 550170 531474 550226
rect 531530 550170 531598 550226
rect 531654 550170 531722 550226
rect 531778 550170 531846 550226
rect 531902 550170 531998 550226
rect 531378 550102 531998 550170
rect 531378 550046 531474 550102
rect 531530 550046 531598 550102
rect 531654 550046 531722 550102
rect 531778 550046 531846 550102
rect 531902 550046 531998 550102
rect 531378 549978 531998 550046
rect 531378 549922 531474 549978
rect 531530 549922 531598 549978
rect 531654 549922 531722 549978
rect 531778 549922 531846 549978
rect 531902 549922 531998 549978
rect 531378 532350 531998 549922
rect 535276 551236 535332 551246
rect 534268 549892 534324 549902
rect 534268 548548 534324 549836
rect 534268 548482 534324 548492
rect 535164 547876 535220 547886
rect 531378 532294 531474 532350
rect 531530 532294 531598 532350
rect 531654 532294 531722 532350
rect 531778 532294 531846 532350
rect 531902 532294 531998 532350
rect 531378 532226 531998 532294
rect 531378 532170 531474 532226
rect 531530 532170 531598 532226
rect 531654 532170 531722 532226
rect 531778 532170 531846 532226
rect 531902 532170 531998 532226
rect 531378 532102 531998 532170
rect 531378 532046 531474 532102
rect 531530 532046 531598 532102
rect 531654 532046 531722 532102
rect 531778 532046 531846 532102
rect 531902 532046 531998 532102
rect 531378 531978 531998 532046
rect 531378 531922 531474 531978
rect 531530 531922 531598 531978
rect 531654 531922 531722 531978
rect 531778 531922 531846 531978
rect 531902 531922 531998 531978
rect 531378 514350 531998 531922
rect 531378 514294 531474 514350
rect 531530 514294 531598 514350
rect 531654 514294 531722 514350
rect 531778 514294 531846 514350
rect 531902 514294 531998 514350
rect 531378 514226 531998 514294
rect 531378 514170 531474 514226
rect 531530 514170 531598 514226
rect 531654 514170 531722 514226
rect 531778 514170 531846 514226
rect 531902 514170 531998 514226
rect 531378 514102 531998 514170
rect 531378 514046 531474 514102
rect 531530 514046 531598 514102
rect 531654 514046 531722 514102
rect 531778 514046 531846 514102
rect 531902 514046 531998 514102
rect 531378 513978 531998 514046
rect 531378 513922 531474 513978
rect 531530 513922 531598 513978
rect 531654 513922 531722 513978
rect 531778 513922 531846 513978
rect 531902 513922 531998 513978
rect 531378 496350 531998 513922
rect 535052 547204 535108 547214
rect 535052 506660 535108 547148
rect 535164 509908 535220 547820
rect 535276 516740 535332 551180
rect 535388 543844 535444 543854
rect 535388 533428 535444 543788
rect 535388 533362 535444 533372
rect 535500 528052 535556 552524
rect 558378 550974 558998 561922
rect 562098 598172 562718 598268
rect 562098 598116 562194 598172
rect 562250 598116 562318 598172
rect 562374 598116 562442 598172
rect 562498 598116 562566 598172
rect 562622 598116 562718 598172
rect 562098 598048 562718 598116
rect 562098 597992 562194 598048
rect 562250 597992 562318 598048
rect 562374 597992 562442 598048
rect 562498 597992 562566 598048
rect 562622 597992 562718 598048
rect 562098 597924 562718 597992
rect 562098 597868 562194 597924
rect 562250 597868 562318 597924
rect 562374 597868 562442 597924
rect 562498 597868 562566 597924
rect 562622 597868 562718 597924
rect 562098 597800 562718 597868
rect 562098 597744 562194 597800
rect 562250 597744 562318 597800
rect 562374 597744 562442 597800
rect 562498 597744 562566 597800
rect 562622 597744 562718 597800
rect 562098 586350 562718 597744
rect 562098 586294 562194 586350
rect 562250 586294 562318 586350
rect 562374 586294 562442 586350
rect 562498 586294 562566 586350
rect 562622 586294 562718 586350
rect 562098 586226 562718 586294
rect 562098 586170 562194 586226
rect 562250 586170 562318 586226
rect 562374 586170 562442 586226
rect 562498 586170 562566 586226
rect 562622 586170 562718 586226
rect 562098 586102 562718 586170
rect 562098 586046 562194 586102
rect 562250 586046 562318 586102
rect 562374 586046 562442 586102
rect 562498 586046 562566 586102
rect 562622 586046 562718 586102
rect 562098 585978 562718 586046
rect 562098 585922 562194 585978
rect 562250 585922 562318 585978
rect 562374 585922 562442 585978
rect 562498 585922 562566 585978
rect 562622 585922 562718 585978
rect 562098 568350 562718 585922
rect 562098 568294 562194 568350
rect 562250 568294 562318 568350
rect 562374 568294 562442 568350
rect 562498 568294 562566 568350
rect 562622 568294 562718 568350
rect 562098 568226 562718 568294
rect 562098 568170 562194 568226
rect 562250 568170 562318 568226
rect 562374 568170 562442 568226
rect 562498 568170 562566 568226
rect 562622 568170 562718 568226
rect 562098 568102 562718 568170
rect 562098 568046 562194 568102
rect 562250 568046 562318 568102
rect 562374 568046 562442 568102
rect 562498 568046 562566 568102
rect 562622 568046 562718 568102
rect 562098 567978 562718 568046
rect 562098 567922 562194 567978
rect 562250 567922 562318 567978
rect 562374 567922 562442 567978
rect 562498 567922 562566 567978
rect 562622 567922 562718 567978
rect 557808 550350 558128 550384
rect 557808 550294 557878 550350
rect 557934 550294 558002 550350
rect 558058 550294 558128 550350
rect 557808 550226 558128 550294
rect 557808 550170 557878 550226
rect 557934 550170 558002 550226
rect 558058 550170 558128 550226
rect 557808 550102 558128 550170
rect 557808 550046 557878 550102
rect 557934 550046 558002 550102
rect 558058 550046 558128 550102
rect 557808 549978 558128 550046
rect 557808 549922 557878 549978
rect 557934 549922 558002 549978
rect 558058 549922 558128 549978
rect 557808 549888 558128 549922
rect 562098 550350 562718 567922
rect 589098 597212 589718 598268
rect 589098 597156 589194 597212
rect 589250 597156 589318 597212
rect 589374 597156 589442 597212
rect 589498 597156 589566 597212
rect 589622 597156 589718 597212
rect 589098 597088 589718 597156
rect 589098 597032 589194 597088
rect 589250 597032 589318 597088
rect 589374 597032 589442 597088
rect 589498 597032 589566 597088
rect 589622 597032 589718 597088
rect 589098 596964 589718 597032
rect 589098 596908 589194 596964
rect 589250 596908 589318 596964
rect 589374 596908 589442 596964
rect 589498 596908 589566 596964
rect 589622 596908 589718 596964
rect 589098 596840 589718 596908
rect 589098 596784 589194 596840
rect 589250 596784 589318 596840
rect 589374 596784 589442 596840
rect 589498 596784 589566 596840
rect 589622 596784 589718 596840
rect 589098 580350 589718 596784
rect 589098 580294 589194 580350
rect 589250 580294 589318 580350
rect 589374 580294 589442 580350
rect 589498 580294 589566 580350
rect 589622 580294 589718 580350
rect 589098 580226 589718 580294
rect 589098 580170 589194 580226
rect 589250 580170 589318 580226
rect 589374 580170 589442 580226
rect 589498 580170 589566 580226
rect 589622 580170 589718 580226
rect 589098 580102 589718 580170
rect 589098 580046 589194 580102
rect 589250 580046 589318 580102
rect 589374 580046 589442 580102
rect 589498 580046 589566 580102
rect 589622 580046 589718 580102
rect 589098 579978 589718 580046
rect 589098 579922 589194 579978
rect 589250 579922 589318 579978
rect 589374 579922 589442 579978
rect 589498 579922 589566 579978
rect 589622 579922 589718 579978
rect 585452 566938 585508 566948
rect 583212 564004 583268 564014
rect 573168 562350 573488 562384
rect 573168 562294 573238 562350
rect 573294 562294 573362 562350
rect 573418 562294 573488 562350
rect 573168 562226 573488 562294
rect 573168 562170 573238 562226
rect 573294 562170 573362 562226
rect 573418 562170 573488 562226
rect 573168 562102 573488 562170
rect 573168 562046 573238 562102
rect 573294 562046 573362 562102
rect 573418 562046 573488 562102
rect 573168 561978 573488 562046
rect 573168 561922 573238 561978
rect 573294 561922 573362 561978
rect 573418 561922 573488 561978
rect 573168 561888 573488 561922
rect 562098 550294 562194 550350
rect 562250 550294 562318 550350
rect 562374 550294 562442 550350
rect 562498 550294 562566 550350
rect 562622 550294 562718 550350
rect 562098 550226 562718 550294
rect 562098 550170 562194 550226
rect 562250 550170 562318 550226
rect 562374 550170 562442 550226
rect 562498 550170 562566 550226
rect 562622 550170 562718 550226
rect 562098 550102 562718 550170
rect 562098 550046 562194 550102
rect 562250 550046 562318 550102
rect 562374 550046 562442 550102
rect 562498 550046 562566 550102
rect 562622 550046 562718 550102
rect 562098 549978 562718 550046
rect 562098 549922 562194 549978
rect 562250 549922 562318 549978
rect 562374 549922 562442 549978
rect 562498 549922 562566 549978
rect 562622 549922 562718 549978
rect 542448 544350 542768 544384
rect 542448 544294 542518 544350
rect 542574 544294 542642 544350
rect 542698 544294 542768 544350
rect 542448 544226 542768 544294
rect 542448 544170 542518 544226
rect 542574 544170 542642 544226
rect 542698 544170 542768 544226
rect 542448 544102 542768 544170
rect 542448 544046 542518 544102
rect 542574 544046 542642 544102
rect 542698 544046 542768 544102
rect 542448 543978 542768 544046
rect 542448 543922 542518 543978
rect 542574 543922 542642 543978
rect 542698 543922 542768 543978
rect 542448 543888 542768 543922
rect 558378 544350 558998 545554
rect 558378 544294 558474 544350
rect 558530 544294 558598 544350
rect 558654 544294 558722 544350
rect 558778 544294 558846 544350
rect 558902 544294 558998 544350
rect 558378 544226 558998 544294
rect 558378 544170 558474 544226
rect 558530 544170 558598 544226
rect 558654 544170 558722 544226
rect 558778 544170 558846 544226
rect 558902 544170 558998 544226
rect 558378 544102 558998 544170
rect 558378 544046 558474 544102
rect 558530 544046 558598 544102
rect 558654 544046 558722 544102
rect 558778 544046 558846 544102
rect 558902 544046 558998 544102
rect 558378 543978 558998 544046
rect 558378 543922 558474 543978
rect 558530 543922 558598 543978
rect 558654 543922 558722 543978
rect 558778 543922 558846 543978
rect 558902 543922 558998 543978
rect 557808 532350 558128 532384
rect 557808 532294 557878 532350
rect 557934 532294 558002 532350
rect 558058 532294 558128 532350
rect 557808 532226 558128 532294
rect 557808 532170 557878 532226
rect 557934 532170 558002 532226
rect 558058 532170 558128 532226
rect 557808 532102 558128 532170
rect 557808 532046 557878 532102
rect 557934 532046 558002 532102
rect 558058 532046 558128 532102
rect 557808 531978 558128 532046
rect 557808 531922 557878 531978
rect 557934 531922 558002 531978
rect 558058 531922 558128 531978
rect 557808 531888 558128 531922
rect 535500 527986 535556 527996
rect 535276 516674 535332 516684
rect 558378 526350 558998 543922
rect 558378 526294 558474 526350
rect 558530 526294 558598 526350
rect 558654 526294 558722 526350
rect 558778 526294 558846 526350
rect 558902 526294 558998 526350
rect 558378 526226 558998 526294
rect 558378 526170 558474 526226
rect 558530 526170 558598 526226
rect 558654 526170 558722 526226
rect 558778 526170 558846 526226
rect 558902 526170 558998 526226
rect 558378 526102 558998 526170
rect 558378 526046 558474 526102
rect 558530 526046 558598 526102
rect 558654 526046 558722 526102
rect 558778 526046 558846 526102
rect 558902 526046 558998 526102
rect 558378 525978 558998 526046
rect 558378 525922 558474 525978
rect 558530 525922 558598 525978
rect 558654 525922 558722 525978
rect 558778 525922 558846 525978
rect 558902 525922 558998 525978
rect 535164 509842 535220 509852
rect 535052 506594 535108 506604
rect 558378 508350 558998 525922
rect 558378 508294 558474 508350
rect 558530 508294 558598 508350
rect 558654 508294 558722 508350
rect 558778 508294 558846 508350
rect 558902 508294 558998 508350
rect 558378 508226 558998 508294
rect 558378 508170 558474 508226
rect 558530 508170 558598 508226
rect 558654 508170 558722 508226
rect 558778 508170 558846 508226
rect 558902 508170 558998 508226
rect 558378 508102 558998 508170
rect 558378 508046 558474 508102
rect 558530 508046 558598 508102
rect 558654 508046 558722 508102
rect 558778 508046 558846 508102
rect 558902 508046 558998 508102
rect 558378 507978 558998 508046
rect 558378 507922 558474 507978
rect 558530 507922 558598 507978
rect 558654 507922 558722 507978
rect 558778 507922 558846 507978
rect 558902 507922 558998 507978
rect 531378 496294 531474 496350
rect 531530 496294 531598 496350
rect 531654 496294 531722 496350
rect 531778 496294 531846 496350
rect 531902 496294 531998 496350
rect 531378 496226 531998 496294
rect 531378 496170 531474 496226
rect 531530 496170 531598 496226
rect 531654 496170 531722 496226
rect 531778 496170 531846 496226
rect 531902 496170 531998 496226
rect 531378 496102 531998 496170
rect 531378 496046 531474 496102
rect 531530 496046 531598 496102
rect 531654 496046 531722 496102
rect 531778 496046 531846 496102
rect 531902 496046 531998 496102
rect 531378 495978 531998 496046
rect 531378 495922 531474 495978
rect 531530 495922 531598 495978
rect 531654 495922 531722 495978
rect 531778 495922 531846 495978
rect 531902 495922 531998 495978
rect 531378 478350 531998 495922
rect 542448 490350 542768 490384
rect 542448 490294 542518 490350
rect 542574 490294 542642 490350
rect 542698 490294 542768 490350
rect 542448 490226 542768 490294
rect 542448 490170 542518 490226
rect 542574 490170 542642 490226
rect 542698 490170 542768 490226
rect 542448 490102 542768 490170
rect 542448 490046 542518 490102
rect 542574 490046 542642 490102
rect 542698 490046 542768 490102
rect 542448 489978 542768 490046
rect 542448 489922 542518 489978
rect 542574 489922 542642 489978
rect 542698 489922 542768 489978
rect 542448 489888 542768 489922
rect 558378 490350 558998 507922
rect 558378 490294 558474 490350
rect 558530 490294 558598 490350
rect 558654 490294 558722 490350
rect 558778 490294 558846 490350
rect 558902 490294 558998 490350
rect 558378 490226 558998 490294
rect 558378 490170 558474 490226
rect 558530 490170 558598 490226
rect 558654 490170 558722 490226
rect 558778 490170 558846 490226
rect 558902 490170 558998 490226
rect 558378 490102 558998 490170
rect 558378 490046 558474 490102
rect 558530 490046 558598 490102
rect 558654 490046 558722 490102
rect 558778 490046 558846 490102
rect 558902 490046 558998 490102
rect 558378 489978 558998 490046
rect 558378 489922 558474 489978
rect 558530 489922 558598 489978
rect 558654 489922 558722 489978
rect 558778 489922 558846 489978
rect 558902 489922 558998 489978
rect 534268 484708 534324 484718
rect 534268 484612 534324 484622
rect 534268 482020 534324 482030
rect 558378 482014 558998 489922
rect 562098 532350 562718 549922
rect 579628 551236 579684 551246
rect 573168 544350 573488 544384
rect 573168 544294 573238 544350
rect 573294 544294 573362 544350
rect 573418 544294 573488 544350
rect 573168 544226 573488 544294
rect 573168 544170 573238 544226
rect 573294 544170 573362 544226
rect 573418 544170 573488 544226
rect 573168 544102 573488 544170
rect 573168 544046 573238 544102
rect 573294 544046 573362 544102
rect 573418 544046 573488 544102
rect 573168 543978 573488 544046
rect 573168 543922 573238 543978
rect 573294 543922 573362 543978
rect 573418 543922 573488 543978
rect 573168 543888 573488 543922
rect 562098 532294 562194 532350
rect 562250 532294 562318 532350
rect 562374 532294 562442 532350
rect 562498 532294 562566 532350
rect 562622 532294 562718 532350
rect 562098 532226 562718 532294
rect 562098 532170 562194 532226
rect 562250 532170 562318 532226
rect 562374 532170 562442 532226
rect 562498 532170 562566 532226
rect 562622 532170 562718 532226
rect 562098 532102 562718 532170
rect 562098 532046 562194 532102
rect 562250 532046 562318 532102
rect 562374 532046 562442 532102
rect 562498 532046 562566 532102
rect 562622 532046 562718 532102
rect 562098 531978 562718 532046
rect 562098 531922 562194 531978
rect 562250 531922 562318 531978
rect 562374 531922 562442 531978
rect 562498 531922 562566 531978
rect 562622 531922 562718 531978
rect 562098 514350 562718 531922
rect 562098 514294 562194 514350
rect 562250 514294 562318 514350
rect 562374 514294 562442 514350
rect 562498 514294 562566 514350
rect 562622 514294 562718 514350
rect 562098 514226 562718 514294
rect 562098 514170 562194 514226
rect 562250 514170 562318 514226
rect 562374 514170 562442 514226
rect 562498 514170 562566 514226
rect 562622 514170 562718 514226
rect 562098 514102 562718 514170
rect 562098 514046 562194 514102
rect 562250 514046 562318 514102
rect 562374 514046 562442 514102
rect 562498 514046 562566 514102
rect 562622 514046 562718 514102
rect 562098 513978 562718 514046
rect 562098 513922 562194 513978
rect 562250 513922 562318 513978
rect 562374 513922 562442 513978
rect 562498 513922 562566 513978
rect 562622 513922 562718 513978
rect 562098 496350 562718 513922
rect 579628 498036 579684 551180
rect 582428 551124 582484 551134
rect 581308 546532 581364 546542
rect 581308 498596 581364 546476
rect 581420 545860 581476 545870
rect 581420 500276 581476 545804
rect 582428 529956 582484 551068
rect 582428 529890 582484 529900
rect 583100 548548 583156 548558
rect 583100 513268 583156 548492
rect 583212 530180 583268 563948
rect 583436 553252 583492 553262
rect 583212 530114 583268 530124
rect 583324 552580 583380 552590
rect 583324 518308 583380 552524
rect 583324 518242 583380 518252
rect 583100 513202 583156 513212
rect 583436 503188 583492 553196
rect 583436 503122 583492 503132
rect 581420 500210 581476 500220
rect 581308 498530 581364 498540
rect 579628 497970 579684 497980
rect 562098 496294 562194 496350
rect 562250 496294 562318 496350
rect 562374 496294 562442 496350
rect 562498 496294 562566 496350
rect 562622 496294 562718 496350
rect 562098 496226 562718 496294
rect 562098 496170 562194 496226
rect 562250 496170 562318 496226
rect 562374 496170 562442 496226
rect 562498 496170 562566 496226
rect 562622 496170 562718 496226
rect 562098 496102 562718 496170
rect 562098 496046 562194 496102
rect 562250 496046 562318 496102
rect 562374 496046 562442 496102
rect 562498 496046 562566 496102
rect 562622 496046 562718 496102
rect 562098 495978 562718 496046
rect 562098 495922 562194 495978
rect 562250 495922 562318 495978
rect 562374 495922 562442 495978
rect 562498 495922 562566 495978
rect 562622 495922 562718 495978
rect 534268 479668 534324 481964
rect 534268 479602 534324 479612
rect 535052 481348 535108 481358
rect 531378 478294 531474 478350
rect 531530 478294 531598 478350
rect 531654 478294 531722 478350
rect 531778 478294 531846 478350
rect 531902 478294 531998 478350
rect 531378 478226 531998 478294
rect 531378 478170 531474 478226
rect 531530 478170 531598 478226
rect 531654 478170 531722 478226
rect 531778 478170 531846 478226
rect 531902 478170 531998 478226
rect 531378 478102 531998 478170
rect 531378 478046 531474 478102
rect 531530 478046 531598 478102
rect 531654 478046 531722 478102
rect 531778 478046 531846 478102
rect 531902 478046 531998 478102
rect 531378 477978 531998 478046
rect 531378 477922 531474 477978
rect 531530 477922 531598 477978
rect 531654 477922 531722 477978
rect 531778 477922 531846 477978
rect 531902 477922 531998 477978
rect 531378 460350 531998 477922
rect 531378 460294 531474 460350
rect 531530 460294 531598 460350
rect 531654 460294 531722 460350
rect 531778 460294 531846 460350
rect 531902 460294 531998 460350
rect 531378 460226 531998 460294
rect 531378 460170 531474 460226
rect 531530 460170 531598 460226
rect 531654 460170 531722 460226
rect 531778 460170 531846 460226
rect 531902 460170 531998 460226
rect 531378 460102 531998 460170
rect 531378 460046 531474 460102
rect 531530 460046 531598 460102
rect 531654 460046 531722 460102
rect 531778 460046 531846 460102
rect 531902 460046 531998 460102
rect 531378 459978 531998 460046
rect 531378 459922 531474 459978
rect 531530 459922 531598 459978
rect 531654 459922 531722 459978
rect 531778 459922 531846 459978
rect 531902 459922 531998 459978
rect 531378 442350 531998 459922
rect 535052 449540 535108 481292
rect 554316 480538 554372 480548
rect 535052 449474 535108 449484
rect 535164 474628 535220 474638
rect 535164 447748 535220 474572
rect 554316 473698 554372 480482
rect 557808 478350 558128 478384
rect 557808 478294 557878 478350
rect 557934 478294 558002 478350
rect 558058 478294 558128 478350
rect 557808 478226 558128 478294
rect 557808 478170 557878 478226
rect 557934 478170 558002 478226
rect 558058 478170 558128 478226
rect 557808 478102 558128 478170
rect 557808 478046 557878 478102
rect 557934 478046 558002 478102
rect 558058 478046 558128 478102
rect 557808 477978 558128 478046
rect 557808 477922 557878 477978
rect 557934 477922 558002 477978
rect 558058 477922 558128 477978
rect 557808 477888 558128 477922
rect 562098 478350 562718 495922
rect 573168 490350 573488 490384
rect 573168 490294 573238 490350
rect 573294 490294 573362 490350
rect 573418 490294 573488 490350
rect 573168 490226 573488 490294
rect 573168 490170 573238 490226
rect 573294 490170 573362 490226
rect 573418 490170 573488 490226
rect 573168 490102 573488 490170
rect 573168 490046 573238 490102
rect 573294 490046 573362 490102
rect 573418 490046 573488 490102
rect 573168 489978 573488 490046
rect 573168 489922 573238 489978
rect 573294 489922 573362 489978
rect 573418 489922 573488 489978
rect 573168 489888 573488 489922
rect 581308 482692 581364 482702
rect 579628 480538 579684 480548
rect 579628 478436 579684 480482
rect 579628 478370 579684 478380
rect 562098 478294 562194 478350
rect 562250 478294 562318 478350
rect 562374 478294 562442 478350
rect 562498 478294 562566 478350
rect 562622 478294 562718 478350
rect 562098 478226 562718 478294
rect 562098 478170 562194 478226
rect 562250 478170 562318 478226
rect 562374 478170 562442 478226
rect 562498 478170 562566 478226
rect 562622 478170 562718 478226
rect 562098 478102 562718 478170
rect 562098 478046 562194 478102
rect 562250 478046 562318 478102
rect 562374 478046 562442 478102
rect 562498 478046 562566 478102
rect 562622 478046 562718 478102
rect 562098 477978 562718 478046
rect 562098 477922 562194 477978
rect 562250 477922 562318 477978
rect 562374 477922 562442 477978
rect 562498 477922 562566 477978
rect 562622 477922 562718 477978
rect 554316 473632 554372 473642
rect 542448 472350 542768 472384
rect 542448 472294 542518 472350
rect 542574 472294 542642 472350
rect 542698 472294 542768 472350
rect 542448 472226 542768 472294
rect 542448 472170 542518 472226
rect 542574 472170 542642 472226
rect 542698 472170 542768 472226
rect 542448 472102 542768 472170
rect 542448 472046 542518 472102
rect 542574 472046 542642 472102
rect 542698 472046 542768 472102
rect 542448 471978 542768 472046
rect 542448 471922 542518 471978
rect 542574 471922 542642 471978
rect 542698 471922 542768 471978
rect 542448 471888 542768 471922
rect 554092 470458 554148 470468
rect 554092 468478 554148 470402
rect 554092 468412 554148 468422
rect 557808 460350 558128 460384
rect 557808 460294 557878 460350
rect 557934 460294 558002 460350
rect 558058 460294 558128 460350
rect 557808 460226 558128 460294
rect 557808 460170 557878 460226
rect 557934 460170 558002 460226
rect 558058 460170 558128 460226
rect 557808 460102 558128 460170
rect 557808 460046 557878 460102
rect 557934 460046 558002 460102
rect 558058 460046 558128 460102
rect 557808 459978 558128 460046
rect 557808 459922 557878 459978
rect 557934 459922 558002 459978
rect 558058 459922 558128 459978
rect 557808 459888 558128 459922
rect 535164 447682 535220 447692
rect 558378 454350 558998 468754
rect 558378 454294 558474 454350
rect 558530 454294 558598 454350
rect 558654 454294 558722 454350
rect 558778 454294 558846 454350
rect 558902 454294 558998 454350
rect 558378 454226 558998 454294
rect 558378 454170 558474 454226
rect 558530 454170 558598 454226
rect 558654 454170 558722 454226
rect 558778 454170 558846 454226
rect 558902 454170 558998 454226
rect 558378 454102 558998 454170
rect 558378 454046 558474 454102
rect 558530 454046 558598 454102
rect 558654 454046 558722 454102
rect 558778 454046 558846 454102
rect 558902 454046 558998 454102
rect 558378 453978 558998 454046
rect 558378 453922 558474 453978
rect 558530 453922 558598 453978
rect 558654 453922 558722 453978
rect 558778 453922 558846 453978
rect 558902 453922 558998 453978
rect 531378 442294 531474 442350
rect 531530 442294 531598 442350
rect 531654 442294 531722 442350
rect 531778 442294 531846 442350
rect 531902 442294 531998 442350
rect 531378 442226 531998 442294
rect 531378 442170 531474 442226
rect 531530 442170 531598 442226
rect 531654 442170 531722 442226
rect 531778 442170 531846 442226
rect 531902 442170 531998 442226
rect 531378 442102 531998 442170
rect 531378 442046 531474 442102
rect 531530 442046 531598 442102
rect 531654 442046 531722 442102
rect 531778 442046 531846 442102
rect 531902 442046 531998 442102
rect 531378 441978 531998 442046
rect 531378 441922 531474 441978
rect 531530 441922 531598 441978
rect 531654 441922 531722 441978
rect 531778 441922 531846 441978
rect 531902 441922 531998 441978
rect 531378 424350 531998 441922
rect 531378 424294 531474 424350
rect 531530 424294 531598 424350
rect 531654 424294 531722 424350
rect 531778 424294 531846 424350
rect 531902 424294 531998 424350
rect 531378 424226 531998 424294
rect 531378 424170 531474 424226
rect 531530 424170 531598 424226
rect 531654 424170 531722 424226
rect 531778 424170 531846 424226
rect 531902 424170 531998 424226
rect 531378 424102 531998 424170
rect 531378 424046 531474 424102
rect 531530 424046 531598 424102
rect 531654 424046 531722 424102
rect 531778 424046 531846 424102
rect 531902 424046 531998 424102
rect 531378 423978 531998 424046
rect 531378 423922 531474 423978
rect 531530 423922 531598 423978
rect 531654 423922 531722 423978
rect 531778 423922 531846 423978
rect 531902 423922 531998 423978
rect 527658 400294 527754 400350
rect 527810 400294 527878 400350
rect 527934 400294 528002 400350
rect 528058 400294 528126 400350
rect 528182 400294 528278 400350
rect 527658 400226 528278 400294
rect 527658 400170 527754 400226
rect 527810 400170 527878 400226
rect 527934 400170 528002 400226
rect 528058 400170 528126 400226
rect 528182 400170 528278 400226
rect 527658 400102 528278 400170
rect 527658 400046 527754 400102
rect 527810 400046 527878 400102
rect 527934 400046 528002 400102
rect 528058 400046 528126 400102
rect 528182 400046 528278 400102
rect 527658 399978 528278 400046
rect 527658 399922 527754 399978
rect 527810 399922 527878 399978
rect 527934 399922 528002 399978
rect 528058 399922 528126 399978
rect 528182 399922 528278 399978
rect 519932 375890 519988 375900
rect 527658 382350 528278 399922
rect 527658 382294 527754 382350
rect 527810 382294 527878 382350
rect 527934 382294 528002 382350
rect 528058 382294 528126 382350
rect 528182 382294 528278 382350
rect 527658 382226 528278 382294
rect 527658 382170 527754 382226
rect 527810 382170 527878 382226
rect 527934 382170 528002 382226
rect 528058 382170 528126 382226
rect 528182 382170 528278 382226
rect 527658 382102 528278 382170
rect 527658 382046 527754 382102
rect 527810 382046 527878 382102
rect 527934 382046 528002 382102
rect 528058 382046 528126 382102
rect 528182 382046 528278 382102
rect 527658 381978 528278 382046
rect 527658 381922 527754 381978
rect 527810 381922 527878 381978
rect 527934 381922 528002 381978
rect 528058 381922 528126 381978
rect 528182 381922 528278 381978
rect 517468 373650 517524 373660
rect 503132 371410 503188 371420
rect 500658 370294 500754 370350
rect 500810 370294 500878 370350
rect 500934 370294 501002 370350
rect 501058 370294 501126 370350
rect 501182 370294 501278 370350
rect 500658 370226 501278 370294
rect 500658 370170 500754 370226
rect 500810 370170 500878 370226
rect 500934 370170 501002 370226
rect 501058 370170 501126 370226
rect 501182 370170 501278 370226
rect 500658 370102 501278 370170
rect 500658 370046 500754 370102
rect 500810 370046 500878 370102
rect 500934 370046 501002 370102
rect 501058 370046 501126 370102
rect 501182 370046 501278 370102
rect 500658 369978 501278 370046
rect 500658 369922 500754 369978
rect 500810 369922 500878 369978
rect 500934 369922 501002 369978
rect 501058 369922 501126 369978
rect 501182 369922 501278 369978
rect 500658 352350 501278 369922
rect 527658 364350 528278 381922
rect 530012 410788 530068 410798
rect 530012 379316 530068 410732
rect 530012 379250 530068 379260
rect 531378 406350 531998 423922
rect 558378 436350 558998 453922
rect 558378 436294 558474 436350
rect 558530 436294 558598 436350
rect 558654 436294 558722 436350
rect 558778 436294 558846 436350
rect 558902 436294 558998 436350
rect 558378 436226 558998 436294
rect 558378 436170 558474 436226
rect 558530 436170 558598 436226
rect 558654 436170 558722 436226
rect 558778 436170 558846 436226
rect 558902 436170 558998 436226
rect 558378 436102 558998 436170
rect 558378 436046 558474 436102
rect 558530 436046 558598 436102
rect 558654 436046 558722 436102
rect 558778 436046 558846 436102
rect 558902 436046 558998 436102
rect 558378 435978 558998 436046
rect 558378 435922 558474 435978
rect 558530 435922 558598 435978
rect 558654 435922 558722 435978
rect 558778 435922 558846 435978
rect 558902 435922 558998 435978
rect 542448 418350 542768 418384
rect 542448 418294 542518 418350
rect 542574 418294 542642 418350
rect 542698 418294 542768 418350
rect 542448 418226 542768 418294
rect 542448 418170 542518 418226
rect 542574 418170 542642 418226
rect 542698 418170 542768 418226
rect 542448 418102 542768 418170
rect 542448 418046 542518 418102
rect 542574 418046 542642 418102
rect 542698 418046 542768 418102
rect 542448 417978 542768 418046
rect 542448 417922 542518 417978
rect 542574 417922 542642 417978
rect 542698 417922 542768 417978
rect 542448 417888 542768 417922
rect 558378 418350 558998 435922
rect 558378 418294 558474 418350
rect 558530 418294 558598 418350
rect 558654 418294 558722 418350
rect 558778 418294 558846 418350
rect 558902 418294 558998 418350
rect 558378 418226 558998 418294
rect 558378 418170 558474 418226
rect 558530 418170 558598 418226
rect 558654 418170 558722 418226
rect 558778 418170 558846 418226
rect 558902 418170 558998 418226
rect 558378 418102 558998 418170
rect 558378 418046 558474 418102
rect 558530 418046 558598 418102
rect 558654 418046 558722 418102
rect 558778 418046 558846 418102
rect 558902 418046 558998 418102
rect 558378 417978 558998 418046
rect 558378 417922 558474 417978
rect 558530 417922 558598 417978
rect 558654 417922 558722 417978
rect 558778 417922 558846 417978
rect 558902 417922 558998 417978
rect 534380 411460 534436 411470
rect 534268 410116 534324 410126
rect 534268 409618 534324 410060
rect 534380 409978 534436 411404
rect 534380 409912 534436 409922
rect 534268 409552 534324 409562
rect 531378 406294 531474 406350
rect 531530 406294 531598 406350
rect 531654 406294 531722 406350
rect 531778 406294 531846 406350
rect 531902 406294 531998 406350
rect 531378 406226 531998 406294
rect 531378 406170 531474 406226
rect 531530 406170 531598 406226
rect 531654 406170 531722 406226
rect 531778 406170 531846 406226
rect 531902 406170 531998 406226
rect 531378 406102 531998 406170
rect 531378 406046 531474 406102
rect 531530 406046 531598 406102
rect 531654 406046 531722 406102
rect 531778 406046 531846 406102
rect 531902 406046 531998 406102
rect 531378 405978 531998 406046
rect 531378 405922 531474 405978
rect 531530 405922 531598 405978
rect 531654 405922 531722 405978
rect 531778 405922 531846 405978
rect 531902 405922 531998 405978
rect 531378 388350 531998 405922
rect 531378 388294 531474 388350
rect 531530 388294 531598 388350
rect 531654 388294 531722 388350
rect 531778 388294 531846 388350
rect 531902 388294 531998 388350
rect 531378 388226 531998 388294
rect 531378 388170 531474 388226
rect 531530 388170 531598 388226
rect 531654 388170 531722 388226
rect 531778 388170 531846 388226
rect 531902 388170 531998 388226
rect 531378 388102 531998 388170
rect 531378 388046 531474 388102
rect 531530 388046 531598 388102
rect 531654 388046 531722 388102
rect 531778 388046 531846 388102
rect 531902 388046 531998 388102
rect 531378 387978 531998 388046
rect 531378 387922 531474 387978
rect 531530 387922 531598 387978
rect 531654 387922 531722 387978
rect 531778 387922 531846 387978
rect 531902 387922 531998 387978
rect 527658 364294 527754 364350
rect 527810 364294 527878 364350
rect 527934 364294 528002 364350
rect 528058 364294 528126 364350
rect 528182 364294 528278 364350
rect 527658 364226 528278 364294
rect 527658 364170 527754 364226
rect 527810 364170 527878 364226
rect 527934 364170 528002 364226
rect 528058 364170 528126 364226
rect 528182 364170 528278 364226
rect 527658 364102 528278 364170
rect 527658 364046 527754 364102
rect 527810 364046 527878 364102
rect 527934 364046 528002 364102
rect 528058 364046 528126 364102
rect 528182 364046 528278 364102
rect 527658 363978 528278 364046
rect 527658 363922 527754 363978
rect 527810 363922 527878 363978
rect 527934 363922 528002 363978
rect 528058 363922 528126 363978
rect 528182 363922 528278 363978
rect 500658 352294 500754 352350
rect 500810 352294 500878 352350
rect 500934 352294 501002 352350
rect 501058 352294 501126 352350
rect 501182 352294 501278 352350
rect 500658 352226 501278 352294
rect 500658 352170 500754 352226
rect 500810 352170 500878 352226
rect 500934 352170 501002 352226
rect 501058 352170 501126 352226
rect 501182 352170 501278 352226
rect 500658 352102 501278 352170
rect 500658 352046 500754 352102
rect 500810 352046 500878 352102
rect 500934 352046 501002 352102
rect 501058 352046 501126 352102
rect 501182 352046 501278 352102
rect 500658 351978 501278 352046
rect 500658 351922 500754 351978
rect 500810 351922 500878 351978
rect 500934 351922 501002 351978
rect 501058 351922 501126 351978
rect 501182 351922 501278 351978
rect 495808 334350 496128 334384
rect 495808 334294 495878 334350
rect 495934 334294 496002 334350
rect 496058 334294 496128 334350
rect 495808 334226 496128 334294
rect 495808 334170 495878 334226
rect 495934 334170 496002 334226
rect 496058 334170 496128 334226
rect 495808 334102 496128 334170
rect 495808 334046 495878 334102
rect 495934 334046 496002 334102
rect 496058 334046 496128 334102
rect 495808 333978 496128 334046
rect 495808 333922 495878 333978
rect 495934 333922 496002 333978
rect 496058 333922 496128 333978
rect 495808 333888 496128 333922
rect 500658 334350 501278 351922
rect 518252 355460 518308 355470
rect 511168 346350 511488 346384
rect 511168 346294 511238 346350
rect 511294 346294 511362 346350
rect 511418 346294 511488 346350
rect 511168 346226 511488 346294
rect 511168 346170 511238 346226
rect 511294 346170 511362 346226
rect 511418 346170 511488 346226
rect 511168 346102 511488 346170
rect 511168 346046 511238 346102
rect 511294 346046 511362 346102
rect 511418 346046 511488 346102
rect 511168 345978 511488 346046
rect 511168 345922 511238 345978
rect 511294 345922 511362 345978
rect 511418 345922 511488 345978
rect 511168 345888 511488 345922
rect 518252 340340 518308 355404
rect 523292 349498 523348 349508
rect 518252 340274 518308 340284
rect 521052 343558 521108 343568
rect 520940 340138 520996 340148
rect 517468 338878 517524 338888
rect 517468 338772 517524 338822
rect 517468 338706 517524 338716
rect 500658 334294 500754 334350
rect 500810 334294 500878 334350
rect 500934 334294 501002 334350
rect 501058 334294 501126 334350
rect 501182 334294 501278 334350
rect 500658 334226 501278 334294
rect 500658 334170 500754 334226
rect 500810 334170 500878 334226
rect 500934 334170 501002 334226
rect 501058 334170 501126 334226
rect 501182 334170 501278 334226
rect 500658 334102 501278 334170
rect 500658 334046 500754 334102
rect 500810 334046 500878 334102
rect 500934 334046 501002 334102
rect 501058 334046 501126 334102
rect 501182 334046 501278 334102
rect 500658 333978 501278 334046
rect 500658 333922 500754 333978
rect 500810 333922 500878 333978
rect 500934 333922 501002 333978
rect 501058 333922 501126 333978
rect 501182 333922 501278 333978
rect 473228 333442 473284 333452
rect 480448 328350 480768 328384
rect 480448 328294 480518 328350
rect 480574 328294 480642 328350
rect 480698 328294 480768 328350
rect 480448 328226 480768 328294
rect 480448 328170 480518 328226
rect 480574 328170 480642 328226
rect 480698 328170 480768 328226
rect 480448 328102 480768 328170
rect 480448 328046 480518 328102
rect 480574 328046 480642 328102
rect 480698 328046 480768 328102
rect 480448 327978 480768 328046
rect 480448 327922 480518 327978
rect 480574 327922 480642 327978
rect 480698 327922 480768 327978
rect 480448 327888 480768 327922
rect 496938 328350 497558 330274
rect 496938 328294 497034 328350
rect 497090 328294 497158 328350
rect 497214 328294 497282 328350
rect 497338 328294 497406 328350
rect 497462 328294 497558 328350
rect 496938 328226 497558 328294
rect 496938 328170 497034 328226
rect 497090 328170 497158 328226
rect 497214 328170 497282 328226
rect 497338 328170 497406 328226
rect 497462 328170 497558 328226
rect 496938 328102 497558 328170
rect 496938 328046 497034 328102
rect 497090 328046 497158 328102
rect 497214 328046 497282 328102
rect 497338 328046 497406 328102
rect 497462 328046 497558 328102
rect 496938 327978 497558 328046
rect 496938 327922 497034 327978
rect 497090 327922 497158 327978
rect 497214 327922 497282 327978
rect 497338 327922 497406 327978
rect 497462 327922 497558 327978
rect 473116 318434 473172 318444
rect 472892 318322 472948 318332
rect 469938 316294 470034 316350
rect 470090 316294 470158 316350
rect 470214 316294 470282 316350
rect 470338 316294 470406 316350
rect 470462 316294 470558 316350
rect 469938 316226 470558 316294
rect 469938 316170 470034 316226
rect 470090 316170 470158 316226
rect 470214 316170 470282 316226
rect 470338 316170 470406 316226
rect 470462 316170 470558 316226
rect 469938 316102 470558 316170
rect 469938 316046 470034 316102
rect 470090 316046 470158 316102
rect 470214 316046 470282 316102
rect 470338 316046 470406 316102
rect 470462 316046 470558 316102
rect 469938 315978 470558 316046
rect 469938 315922 470034 315978
rect 470090 315922 470158 315978
rect 470214 315922 470282 315978
rect 470338 315922 470406 315978
rect 470462 315922 470558 315978
rect 469938 298350 470558 315922
rect 469938 298294 470034 298350
rect 470090 298294 470158 298350
rect 470214 298294 470282 298350
rect 470338 298294 470406 298350
rect 470462 298294 470558 298350
rect 469938 298226 470558 298294
rect 469938 298170 470034 298226
rect 470090 298170 470158 298226
rect 470214 298170 470282 298226
rect 470338 298170 470406 298226
rect 470462 298170 470558 298226
rect 469938 298102 470558 298170
rect 469938 298046 470034 298102
rect 470090 298046 470158 298102
rect 470214 298046 470282 298102
rect 470338 298046 470406 298102
rect 470462 298046 470558 298102
rect 469938 297978 470558 298046
rect 469938 297922 470034 297978
rect 470090 297922 470158 297978
rect 470214 297922 470282 297978
rect 470338 297922 470406 297978
rect 470462 297922 470558 297978
rect 469938 280350 470558 297922
rect 496938 310350 497558 327922
rect 496938 310294 497034 310350
rect 497090 310294 497158 310350
rect 497214 310294 497282 310350
rect 497338 310294 497406 310350
rect 497462 310294 497558 310350
rect 496938 310226 497558 310294
rect 496938 310170 497034 310226
rect 497090 310170 497158 310226
rect 497214 310170 497282 310226
rect 497338 310170 497406 310226
rect 497462 310170 497558 310226
rect 496938 310102 497558 310170
rect 496938 310046 497034 310102
rect 497090 310046 497158 310102
rect 497214 310046 497282 310102
rect 497338 310046 497406 310102
rect 497462 310046 497558 310102
rect 496938 309978 497558 310046
rect 496938 309922 497034 309978
rect 497090 309922 497158 309978
rect 497214 309922 497282 309978
rect 497338 309922 497406 309978
rect 497462 309922 497558 309978
rect 496938 292350 497558 309922
rect 496938 292294 497034 292350
rect 497090 292294 497158 292350
rect 497214 292294 497282 292350
rect 497338 292294 497406 292350
rect 497462 292294 497558 292350
rect 496938 292226 497558 292294
rect 496938 292170 497034 292226
rect 497090 292170 497158 292226
rect 497214 292170 497282 292226
rect 497338 292170 497406 292226
rect 497462 292170 497558 292226
rect 496938 292102 497558 292170
rect 496938 292046 497034 292102
rect 497090 292046 497158 292102
rect 497214 292046 497282 292102
rect 497338 292046 497406 292102
rect 497462 292046 497558 292102
rect 496938 291978 497558 292046
rect 496938 291922 497034 291978
rect 497090 291922 497158 291978
rect 497214 291922 497282 291978
rect 497338 291922 497406 291978
rect 497462 291922 497558 291978
rect 473116 284564 473172 284574
rect 469938 280294 470034 280350
rect 470090 280294 470158 280350
rect 470214 280294 470282 280350
rect 470338 280294 470406 280350
rect 470462 280294 470558 280350
rect 469938 280226 470558 280294
rect 469938 280170 470034 280226
rect 470090 280170 470158 280226
rect 470214 280170 470282 280226
rect 470338 280170 470406 280226
rect 470462 280170 470558 280226
rect 469938 280102 470558 280170
rect 469938 280046 470034 280102
rect 470090 280046 470158 280102
rect 470214 280046 470282 280102
rect 470338 280046 470406 280102
rect 470462 280046 470558 280102
rect 469938 279978 470558 280046
rect 469938 279922 470034 279978
rect 470090 279922 470158 279978
rect 470214 279922 470282 279978
rect 470338 279922 470406 279978
rect 470462 279922 470558 279978
rect 469938 262350 470558 279922
rect 472892 283220 472948 283230
rect 472108 269108 472164 269118
rect 472108 269038 472164 269052
rect 472108 268972 472164 268982
rect 472108 268436 472164 268446
rect 472108 267418 472164 268380
rect 472108 267352 472164 267362
rect 472108 266420 472164 266430
rect 472108 264628 472164 266364
rect 472108 264562 472164 264572
rect 472892 263732 472948 283164
rect 473116 283220 473172 284508
rect 473116 283154 473172 283164
rect 495808 280350 496128 280384
rect 495808 280294 495878 280350
rect 495934 280294 496002 280350
rect 496058 280294 496128 280350
rect 495808 280226 496128 280294
rect 495808 280170 495878 280226
rect 495934 280170 496002 280226
rect 496058 280170 496128 280226
rect 495808 280102 496128 280170
rect 495808 280046 495878 280102
rect 495934 280046 496002 280102
rect 496058 280046 496128 280102
rect 495808 279978 496128 280046
rect 495808 279922 495878 279978
rect 495934 279922 496002 279978
rect 496058 279922 496128 279978
rect 495808 279888 496128 279922
rect 480448 274350 480768 274384
rect 480448 274294 480518 274350
rect 480574 274294 480642 274350
rect 480698 274294 480768 274350
rect 480448 274226 480768 274294
rect 480448 274170 480518 274226
rect 480574 274170 480642 274226
rect 480698 274170 480768 274226
rect 480448 274102 480768 274170
rect 480448 274046 480518 274102
rect 480574 274046 480642 274102
rect 480698 274046 480768 274102
rect 480448 273978 480768 274046
rect 480448 273922 480518 273978
rect 480574 273922 480642 273978
rect 480698 273922 480768 273978
rect 480448 273888 480768 273922
rect 496938 274350 497558 291922
rect 496938 274294 497034 274350
rect 497090 274294 497158 274350
rect 497214 274294 497282 274350
rect 497338 274294 497406 274350
rect 497462 274294 497558 274350
rect 496938 274226 497558 274294
rect 496938 274170 497034 274226
rect 497090 274170 497158 274226
rect 497214 274170 497282 274226
rect 497338 274170 497406 274226
rect 497462 274170 497558 274226
rect 496938 274102 497558 274170
rect 496938 274046 497034 274102
rect 497090 274046 497158 274102
rect 497214 274046 497282 274102
rect 497338 274046 497406 274102
rect 497462 274046 497558 274102
rect 496938 273978 497558 274046
rect 496938 273922 497034 273978
rect 497090 273922 497158 273978
rect 497214 273922 497282 273978
rect 497338 273922 497406 273978
rect 497462 273922 497558 273978
rect 473004 271348 473060 271358
rect 473004 264404 473060 271292
rect 473676 269780 473732 269790
rect 473676 269578 473732 269724
rect 473676 269512 473732 269522
rect 496938 268414 497558 273922
rect 500658 316350 501278 333922
rect 517468 337652 517524 337662
rect 511168 328350 511488 328384
rect 511168 328294 511238 328350
rect 511294 328294 511362 328350
rect 511418 328294 511488 328350
rect 511168 328226 511488 328294
rect 511168 328170 511238 328226
rect 511294 328170 511362 328226
rect 511418 328170 511488 328226
rect 511168 328102 511488 328170
rect 511168 328046 511238 328102
rect 511294 328046 511362 328102
rect 511418 328046 511488 328102
rect 511168 327978 511488 328046
rect 511168 327922 511238 327978
rect 511294 327922 511362 327978
rect 511418 327922 511488 327978
rect 511168 327888 511488 327922
rect 500658 316294 500754 316350
rect 500810 316294 500878 316350
rect 500934 316294 501002 316350
rect 501058 316294 501126 316350
rect 501182 316294 501278 316350
rect 500658 316226 501278 316294
rect 500658 316170 500754 316226
rect 500810 316170 500878 316226
rect 500934 316170 501002 316226
rect 501058 316170 501126 316226
rect 501182 316170 501278 316226
rect 500658 316102 501278 316170
rect 500658 316046 500754 316102
rect 500810 316046 500878 316102
rect 500934 316046 501002 316102
rect 501058 316046 501126 316102
rect 501182 316046 501278 316102
rect 500658 315978 501278 316046
rect 500658 315922 500754 315978
rect 500810 315922 500878 315978
rect 500934 315922 501002 315978
rect 501058 315922 501126 315978
rect 501182 315922 501278 315978
rect 500658 298350 501278 315922
rect 517468 314356 517524 337596
rect 520828 336980 520884 336990
rect 519148 335636 519204 335646
rect 519148 316596 519204 335580
rect 520828 317604 520884 336924
rect 520940 332276 520996 340082
rect 521052 332948 521108 343502
rect 521052 332882 521108 332892
rect 523292 332948 523348 349442
rect 523292 332882 523348 332892
rect 527658 346350 528278 363922
rect 527658 346294 527754 346350
rect 527810 346294 527878 346350
rect 527934 346294 528002 346350
rect 528058 346294 528126 346350
rect 528182 346294 528278 346350
rect 527658 346226 528278 346294
rect 527658 346170 527754 346226
rect 527810 346170 527878 346226
rect 527934 346170 528002 346226
rect 528058 346170 528126 346226
rect 528182 346170 528278 346226
rect 527658 346102 528278 346170
rect 527658 346046 527754 346102
rect 527810 346046 527878 346102
rect 527934 346046 528002 346102
rect 528058 346046 528126 346102
rect 528182 346046 528278 346102
rect 527658 345978 528278 346046
rect 527658 345922 527754 345978
rect 527810 345922 527878 345978
rect 527934 345922 528002 345978
rect 528058 345922 528126 345978
rect 528182 345922 528278 345978
rect 520940 332210 520996 332220
rect 523292 332276 523348 332286
rect 523292 324118 523348 332220
rect 523292 324052 523348 324062
rect 527658 328350 528278 345922
rect 527658 328294 527754 328350
rect 527810 328294 527878 328350
rect 527934 328294 528002 328350
rect 528058 328294 528126 328350
rect 528182 328294 528278 328350
rect 527658 328226 528278 328294
rect 527658 328170 527754 328226
rect 527810 328170 527878 328226
rect 527934 328170 528002 328226
rect 528058 328170 528126 328226
rect 528182 328170 528278 328226
rect 527658 328102 528278 328170
rect 527658 328046 527754 328102
rect 527810 328046 527878 328102
rect 527934 328046 528002 328102
rect 528058 328046 528126 328102
rect 528182 328046 528278 328102
rect 527658 327978 528278 328046
rect 527658 327922 527754 327978
rect 527810 327922 527878 327978
rect 527934 327922 528002 327978
rect 528058 327922 528126 327978
rect 528182 327922 528278 327978
rect 520828 317538 520884 317548
rect 519148 316530 519204 316540
rect 517468 314290 517524 314300
rect 500658 298294 500754 298350
rect 500810 298294 500878 298350
rect 500934 298294 501002 298350
rect 501058 298294 501126 298350
rect 501182 298294 501278 298350
rect 500658 298226 501278 298294
rect 500658 298170 500754 298226
rect 500810 298170 500878 298226
rect 500934 298170 501002 298226
rect 501058 298170 501126 298226
rect 501182 298170 501278 298226
rect 500658 298102 501278 298170
rect 500658 298046 500754 298102
rect 500810 298046 500878 298102
rect 500934 298046 501002 298102
rect 501058 298046 501126 298102
rect 501182 298046 501278 298102
rect 500658 297978 501278 298046
rect 500658 297922 500754 297978
rect 500810 297922 500878 297978
rect 500934 297922 501002 297978
rect 501058 297922 501126 297978
rect 501182 297922 501278 297978
rect 500658 280350 501278 297922
rect 527658 310350 528278 327922
rect 527658 310294 527754 310350
rect 527810 310294 527878 310350
rect 527934 310294 528002 310350
rect 528058 310294 528126 310350
rect 528182 310294 528278 310350
rect 527658 310226 528278 310294
rect 527658 310170 527754 310226
rect 527810 310170 527878 310226
rect 527934 310170 528002 310226
rect 528058 310170 528126 310226
rect 528182 310170 528278 310226
rect 527658 310102 528278 310170
rect 527658 310046 527754 310102
rect 527810 310046 527878 310102
rect 527934 310046 528002 310102
rect 528058 310046 528126 310102
rect 528182 310046 528278 310102
rect 527658 309978 528278 310046
rect 527658 309922 527754 309978
rect 527810 309922 527878 309978
rect 527934 309922 528002 309978
rect 528058 309922 528126 309978
rect 528182 309922 528278 309978
rect 523292 293076 523348 293086
rect 502348 291396 502404 291406
rect 502348 286468 502404 291340
rect 502348 286402 502404 286412
rect 517468 289828 517524 289838
rect 500658 280294 500754 280350
rect 500810 280294 500878 280350
rect 500934 280294 501002 280350
rect 501058 280294 501126 280350
rect 501182 280294 501278 280350
rect 500658 280226 501278 280294
rect 500658 280170 500754 280226
rect 500810 280170 500878 280226
rect 500934 280170 501002 280226
rect 501058 280170 501126 280226
rect 501182 280170 501278 280226
rect 500658 280102 501278 280170
rect 500658 280046 500754 280102
rect 500810 280046 500878 280102
rect 500934 280046 501002 280102
rect 501058 280046 501126 280102
rect 501182 280046 501278 280102
rect 500658 279978 501278 280046
rect 500658 279922 500754 279978
rect 500810 279922 500878 279978
rect 500934 279922 501002 279978
rect 501058 279922 501126 279978
rect 501182 279922 501278 279978
rect 500658 268414 501278 279922
rect 511168 274350 511488 274384
rect 511168 274294 511238 274350
rect 511294 274294 511362 274350
rect 511418 274294 511488 274350
rect 511168 274226 511488 274294
rect 511168 274170 511238 274226
rect 511294 274170 511362 274226
rect 511418 274170 511488 274226
rect 511168 274102 511488 274170
rect 511168 274046 511238 274102
rect 511294 274046 511362 274102
rect 511418 274046 511488 274102
rect 511168 273978 511488 274046
rect 511168 273922 511238 273978
rect 511294 273922 511362 273978
rect 511418 273922 511488 273978
rect 511168 273888 511488 273922
rect 517468 273718 517524 289772
rect 517580 289716 517636 289726
rect 517580 273868 517636 289660
rect 519148 289156 519204 289166
rect 517580 273812 517860 273868
rect 517468 273662 517748 273718
rect 517468 267316 517524 267326
rect 517468 267238 517524 267260
rect 517468 267172 517524 267182
rect 473004 264338 473060 264348
rect 472892 263666 472948 263676
rect 469938 262294 470034 262350
rect 470090 262294 470158 262350
rect 470214 262294 470282 262350
rect 470338 262294 470406 262350
rect 470462 262294 470558 262350
rect 469938 262226 470558 262294
rect 469938 262170 470034 262226
rect 470090 262170 470158 262226
rect 470214 262170 470282 262226
rect 470338 262170 470406 262226
rect 470462 262170 470558 262226
rect 469938 262102 470558 262170
rect 468636 262052 468692 262062
rect 468636 258598 468692 261996
rect 468636 258532 468692 258542
rect 469938 262046 470034 262102
rect 470090 262046 470158 262102
rect 470214 262046 470282 262102
rect 470338 262046 470406 262102
rect 470462 262046 470558 262102
rect 469938 261978 470558 262046
rect 469938 261922 470034 261978
rect 470090 261922 470158 261978
rect 470214 261922 470282 261978
rect 470338 261922 470406 261978
rect 470462 261922 470558 261978
rect 466218 256294 466314 256350
rect 466370 256294 466438 256350
rect 466494 256294 466562 256350
rect 466618 256294 466686 256350
rect 466742 256294 466838 256350
rect 466218 256226 466838 256294
rect 466218 256170 466314 256226
rect 466370 256170 466438 256226
rect 466494 256170 466562 256226
rect 466618 256170 466686 256226
rect 466742 256170 466838 256226
rect 466218 256102 466838 256170
rect 466218 256046 466314 256102
rect 466370 256046 466438 256102
rect 466494 256046 466562 256102
rect 466618 256046 466686 256102
rect 466742 256046 466838 256102
rect 466218 255978 466838 256046
rect 466218 255922 466314 255978
rect 466370 255922 466438 255978
rect 466494 255922 466562 255978
rect 466618 255922 466686 255978
rect 466742 255922 466838 255978
rect 461132 255112 461188 255122
rect 458892 250252 458948 250262
rect 439218 244294 439314 244350
rect 439370 244294 439438 244350
rect 439494 244294 439562 244350
rect 439618 244294 439686 244350
rect 439742 244294 439838 244350
rect 439218 244226 439838 244294
rect 439218 244170 439314 244226
rect 439370 244170 439438 244226
rect 439494 244170 439562 244226
rect 439618 244170 439686 244226
rect 439742 244170 439838 244226
rect 439218 244102 439838 244170
rect 439218 244046 439314 244102
rect 439370 244046 439438 244102
rect 439494 244046 439562 244102
rect 439618 244046 439686 244102
rect 439742 244046 439838 244102
rect 439218 243978 439838 244046
rect 439218 243922 439314 243978
rect 439370 243922 439438 243978
rect 439494 243922 439562 243978
rect 439618 243922 439686 243978
rect 439742 243922 439838 243978
rect 439218 226350 439838 243922
rect 466218 238350 466838 255922
rect 466218 238294 466314 238350
rect 466370 238294 466438 238350
rect 466494 238294 466562 238350
rect 466618 238294 466686 238350
rect 466742 238294 466838 238350
rect 466218 238226 466838 238294
rect 466218 238170 466314 238226
rect 466370 238170 466438 238226
rect 466494 238170 466562 238226
rect 466618 238170 466686 238226
rect 466742 238170 466838 238226
rect 466218 238102 466838 238170
rect 466218 238046 466314 238102
rect 466370 238046 466438 238102
rect 466494 238046 466562 238102
rect 466618 238046 466686 238102
rect 466742 238046 466838 238102
rect 466218 237978 466838 238046
rect 466218 237922 466314 237978
rect 466370 237922 466438 237978
rect 466494 237922 466562 237978
rect 466618 237922 466686 237978
rect 466742 237922 466838 237978
rect 439218 226294 439314 226350
rect 439370 226294 439438 226350
rect 439494 226294 439562 226350
rect 439618 226294 439686 226350
rect 439742 226294 439838 226350
rect 439218 226226 439838 226294
rect 439218 226170 439314 226226
rect 439370 226170 439438 226226
rect 439494 226170 439562 226226
rect 439618 226170 439686 226226
rect 439742 226170 439838 226226
rect 439218 226102 439838 226170
rect 439218 226046 439314 226102
rect 439370 226046 439438 226102
rect 439494 226046 439562 226102
rect 439618 226046 439686 226102
rect 439742 226046 439838 226102
rect 439218 225978 439838 226046
rect 439218 225922 439314 225978
rect 439370 225922 439438 225978
rect 439494 225922 439562 225978
rect 439618 225922 439686 225978
rect 439742 225922 439838 225978
rect 439218 208350 439838 225922
rect 459452 234276 459508 234286
rect 439218 208294 439314 208350
rect 439370 208294 439438 208350
rect 439494 208294 439562 208350
rect 439618 208294 439686 208350
rect 439742 208294 439838 208350
rect 439218 208226 439838 208294
rect 455308 222516 455364 222526
rect 455308 208348 455364 222460
rect 456988 217588 457044 217598
rect 455308 208292 455476 208348
rect 439218 208170 439314 208226
rect 439370 208170 439438 208226
rect 439494 208170 439562 208226
rect 439618 208170 439686 208226
rect 439742 208170 439838 208226
rect 439218 208102 439838 208170
rect 439218 208046 439314 208102
rect 439370 208046 439438 208102
rect 439494 208046 439562 208102
rect 439618 208046 439686 208102
rect 439742 208046 439838 208102
rect 439218 207978 439838 208046
rect 439218 207922 439314 207978
rect 439370 207922 439438 207978
rect 439494 207922 439562 207978
rect 439618 207922 439686 207978
rect 439742 207922 439838 207978
rect 439218 190350 439838 207922
rect 449168 202350 449488 202384
rect 449168 202294 449238 202350
rect 449294 202294 449362 202350
rect 449418 202294 449488 202350
rect 449168 202226 449488 202294
rect 449168 202170 449238 202226
rect 449294 202170 449362 202226
rect 449418 202170 449488 202226
rect 449168 202102 449488 202170
rect 449168 202046 449238 202102
rect 449294 202046 449362 202102
rect 449418 202046 449488 202102
rect 449168 201978 449488 202046
rect 449168 201922 449238 201978
rect 449294 201922 449362 201978
rect 449418 201922 449488 201978
rect 449168 201888 449488 201922
rect 455308 198548 455364 198558
rect 455308 198478 455364 198492
rect 455308 198412 455364 198422
rect 455420 196756 455476 208292
rect 455420 196690 455476 196700
rect 456092 196858 456148 196868
rect 455308 194068 455364 194078
rect 455308 193978 455364 194012
rect 455308 193912 455364 193922
rect 439218 190294 439314 190350
rect 439370 190294 439438 190350
rect 439494 190294 439562 190350
rect 439618 190294 439686 190350
rect 439742 190294 439838 190350
rect 439218 190226 439838 190294
rect 439218 190170 439314 190226
rect 439370 190170 439438 190226
rect 439494 190170 439562 190226
rect 439618 190170 439686 190226
rect 439742 190170 439838 190226
rect 439218 190102 439838 190170
rect 439218 190046 439314 190102
rect 439370 190046 439438 190102
rect 439494 190046 439562 190102
rect 439618 190046 439686 190102
rect 439742 190046 439838 190102
rect 439218 189978 439838 190046
rect 439218 189922 439314 189978
rect 439370 189922 439438 189978
rect 439494 189922 439562 189978
rect 439618 189922 439686 189978
rect 439742 189922 439838 189978
rect 439218 172350 439838 189922
rect 455420 192178 455476 192188
rect 455420 189028 455476 192122
rect 455420 188962 455476 188972
rect 455308 186452 455364 186462
rect 455308 186352 455364 186362
rect 456092 186340 456148 196802
rect 456988 193844 457044 217532
rect 458892 214340 458948 214350
rect 456988 193778 457044 193788
rect 458780 213220 458836 213230
rect 458780 191156 458836 213164
rect 458892 191828 458948 214284
rect 459452 214340 459508 234220
rect 459452 214274 459508 214284
rect 462812 232036 462868 232046
rect 462812 211204 462868 231980
rect 462812 211138 462868 211148
rect 466218 220350 466838 237922
rect 466218 220294 466314 220350
rect 466370 220294 466438 220350
rect 466494 220294 466562 220350
rect 466618 220294 466686 220350
rect 466742 220294 466838 220350
rect 466218 220226 466838 220294
rect 466218 220170 466314 220226
rect 466370 220170 466438 220226
rect 466494 220170 466562 220226
rect 466618 220170 466686 220226
rect 466742 220170 466838 220226
rect 466218 220102 466838 220170
rect 466218 220046 466314 220102
rect 466370 220046 466438 220102
rect 466494 220046 466562 220102
rect 466618 220046 466686 220102
rect 466742 220046 466838 220102
rect 466218 219978 466838 220046
rect 466218 219922 466314 219978
rect 466370 219922 466438 219978
rect 466494 219922 466562 219978
rect 466618 219922 466686 219978
rect 466742 219922 466838 219978
rect 466218 202350 466838 219922
rect 466218 202294 466314 202350
rect 466370 202294 466438 202350
rect 466494 202294 466562 202350
rect 466618 202294 466686 202350
rect 466742 202294 466838 202350
rect 466218 202226 466838 202294
rect 466218 202170 466314 202226
rect 466370 202170 466438 202226
rect 466494 202170 466562 202226
rect 466618 202170 466686 202226
rect 466742 202170 466838 202226
rect 466218 202102 466838 202170
rect 466218 202046 466314 202102
rect 466370 202046 466438 202102
rect 466494 202046 466562 202102
rect 466618 202046 466686 202102
rect 466742 202046 466838 202102
rect 466218 201978 466838 202046
rect 466218 201922 466314 201978
rect 466370 201922 466438 201978
rect 466494 201922 466562 201978
rect 466618 201922 466686 201978
rect 466742 201922 466838 201978
rect 463596 196678 463652 196688
rect 463596 192388 463652 196622
rect 463596 192322 463652 192332
rect 458892 191762 458948 191772
rect 458780 191090 458836 191100
rect 456092 186274 456148 186284
rect 449168 184350 449488 184384
rect 449168 184294 449238 184350
rect 449294 184294 449362 184350
rect 449418 184294 449488 184350
rect 449168 184226 449488 184294
rect 449168 184170 449238 184226
rect 449294 184170 449362 184226
rect 449418 184170 449488 184226
rect 449168 184102 449488 184170
rect 449168 184046 449238 184102
rect 449294 184046 449362 184102
rect 449418 184046 449488 184102
rect 449168 183978 449488 184046
rect 449168 183922 449238 183978
rect 449294 183922 449362 183978
rect 449418 183922 449488 183978
rect 449168 183888 449488 183922
rect 466218 184350 466838 201922
rect 469938 244350 470558 261922
rect 495808 262350 496128 262384
rect 495808 262294 495878 262350
rect 495934 262294 496002 262350
rect 496058 262294 496128 262350
rect 495808 262226 496128 262294
rect 495808 262170 495878 262226
rect 495934 262170 496002 262226
rect 496058 262170 496128 262226
rect 495808 262102 496128 262170
rect 495808 262046 495878 262102
rect 495934 262046 496002 262102
rect 496058 262046 496128 262102
rect 495808 261978 496128 262046
rect 495808 261922 495878 261978
rect 495934 261922 496002 261978
rect 496058 261922 496128 261978
rect 495808 261888 496128 261922
rect 472220 261044 472276 261054
rect 472108 260372 472164 260382
rect 472108 258778 472164 260316
rect 472220 259588 472276 260988
rect 472220 259522 472276 259532
rect 472108 258712 472164 258722
rect 480448 256350 480768 256384
rect 480448 256294 480518 256350
rect 480574 256294 480642 256350
rect 480698 256294 480768 256350
rect 480448 256226 480768 256294
rect 480448 256170 480518 256226
rect 480574 256170 480642 256226
rect 480698 256170 480768 256226
rect 480448 256102 480768 256170
rect 480448 256046 480518 256102
rect 480574 256046 480642 256102
rect 480698 256046 480768 256102
rect 480448 255978 480768 256046
rect 480448 255922 480518 255978
rect 480574 255922 480642 255978
rect 480698 255922 480768 255978
rect 480448 255888 480768 255922
rect 496938 256350 497558 262994
rect 496938 256294 497034 256350
rect 497090 256294 497158 256350
rect 497214 256294 497282 256350
rect 497338 256294 497406 256350
rect 497462 256294 497558 256350
rect 496938 256226 497558 256294
rect 496938 256170 497034 256226
rect 497090 256170 497158 256226
rect 497214 256170 497282 256226
rect 497338 256170 497406 256226
rect 497462 256170 497558 256226
rect 496938 256102 497558 256170
rect 496938 256046 497034 256102
rect 497090 256046 497158 256102
rect 497214 256046 497282 256102
rect 497338 256046 497406 256102
rect 497462 256046 497558 256102
rect 496938 255978 497558 256046
rect 496938 255922 497034 255978
rect 497090 255922 497158 255978
rect 497214 255922 497282 255978
rect 497338 255922 497406 255978
rect 497462 255922 497558 255978
rect 469938 244294 470034 244350
rect 470090 244294 470158 244350
rect 470214 244294 470282 244350
rect 470338 244294 470406 244350
rect 470462 244294 470558 244350
rect 469938 244226 470558 244294
rect 469938 244170 470034 244226
rect 470090 244170 470158 244226
rect 470214 244170 470282 244226
rect 470338 244170 470406 244226
rect 470462 244170 470558 244226
rect 469938 244102 470558 244170
rect 469938 244046 470034 244102
rect 470090 244046 470158 244102
rect 470214 244046 470282 244102
rect 470338 244046 470406 244102
rect 470462 244046 470558 244102
rect 469938 243978 470558 244046
rect 469938 243922 470034 243978
rect 470090 243922 470158 243978
rect 470214 243922 470282 243978
rect 470338 243922 470406 243978
rect 470462 243922 470558 243978
rect 469938 226350 470558 243922
rect 469938 226294 470034 226350
rect 470090 226294 470158 226350
rect 470214 226294 470282 226350
rect 470338 226294 470406 226350
rect 470462 226294 470558 226350
rect 469938 226226 470558 226294
rect 469938 226170 470034 226226
rect 470090 226170 470158 226226
rect 470214 226170 470282 226226
rect 470338 226170 470406 226226
rect 470462 226170 470558 226226
rect 469938 226102 470558 226170
rect 469938 226046 470034 226102
rect 470090 226046 470158 226102
rect 470214 226046 470282 226102
rect 470338 226046 470406 226102
rect 470462 226046 470558 226102
rect 469938 225978 470558 226046
rect 469938 225922 470034 225978
rect 470090 225922 470158 225978
rect 470214 225922 470282 225978
rect 470338 225922 470406 225978
rect 470462 225922 470558 225978
rect 469938 208350 470558 225922
rect 496938 238350 497558 255922
rect 496938 238294 497034 238350
rect 497090 238294 497158 238350
rect 497214 238294 497282 238350
rect 497338 238294 497406 238350
rect 497462 238294 497558 238350
rect 496938 238226 497558 238294
rect 496938 238170 497034 238226
rect 497090 238170 497158 238226
rect 497214 238170 497282 238226
rect 497338 238170 497406 238226
rect 497462 238170 497558 238226
rect 496938 238102 497558 238170
rect 496938 238046 497034 238102
rect 497090 238046 497158 238102
rect 497214 238046 497282 238102
rect 497338 238046 497406 238102
rect 497462 238046 497558 238102
rect 496938 237978 497558 238046
rect 496938 237922 497034 237978
rect 497090 237922 497158 237978
rect 497214 237922 497282 237978
rect 497338 237922 497406 237978
rect 497462 237922 497558 237978
rect 496938 220350 497558 237922
rect 496938 220294 497034 220350
rect 497090 220294 497158 220350
rect 497214 220294 497282 220350
rect 497338 220294 497406 220350
rect 497462 220294 497558 220350
rect 496938 220226 497558 220294
rect 496938 220170 497034 220226
rect 497090 220170 497158 220226
rect 497214 220170 497282 220226
rect 497338 220170 497406 220226
rect 497462 220170 497558 220226
rect 496938 220102 497558 220170
rect 496938 220046 497034 220102
rect 497090 220046 497158 220102
rect 497214 220046 497282 220102
rect 497338 220046 497406 220102
rect 497462 220046 497558 220102
rect 496938 219978 497558 220046
rect 496938 219922 497034 219978
rect 497090 219922 497158 219978
rect 497214 219922 497282 219978
rect 497338 219922 497406 219978
rect 497462 219922 497558 219978
rect 472108 214228 472164 214238
rect 472108 208628 472164 214172
rect 472108 208562 472164 208572
rect 469938 208294 470034 208350
rect 470090 208294 470158 208350
rect 470214 208294 470282 208350
rect 470338 208294 470406 208350
rect 470462 208294 470558 208350
rect 469938 208226 470558 208294
rect 469938 208170 470034 208226
rect 470090 208170 470158 208226
rect 470214 208170 470282 208226
rect 470338 208170 470406 208226
rect 470462 208170 470558 208226
rect 469938 208102 470558 208170
rect 469938 208046 470034 208102
rect 470090 208046 470158 208102
rect 470214 208046 470282 208102
rect 470338 208046 470406 208102
rect 470462 208046 470558 208102
rect 469938 207978 470558 208046
rect 469938 207922 470034 207978
rect 470090 207922 470158 207978
rect 470214 207922 470282 207978
rect 470338 207922 470406 207978
rect 470462 207922 470558 207978
rect 467852 200098 467908 200108
rect 467852 196532 467908 200042
rect 467852 196466 467908 196476
rect 466218 184294 466314 184350
rect 466370 184294 466438 184350
rect 466494 184294 466562 184350
rect 466618 184294 466686 184350
rect 466742 184294 466838 184350
rect 466218 184226 466838 184294
rect 466218 184170 466314 184226
rect 466370 184170 466438 184226
rect 466494 184170 466562 184226
rect 466618 184170 466686 184226
rect 466742 184170 466838 184226
rect 466218 184102 466838 184170
rect 466218 184046 466314 184102
rect 466370 184046 466438 184102
rect 466494 184046 466562 184102
rect 466618 184046 466686 184102
rect 466742 184046 466838 184102
rect 466218 183978 466838 184046
rect 466218 183922 466314 183978
rect 466370 183922 466438 183978
rect 466494 183922 466562 183978
rect 466618 183922 466686 183978
rect 466742 183922 466838 183978
rect 439218 172294 439314 172350
rect 439370 172294 439438 172350
rect 439494 172294 439562 172350
rect 439618 172294 439686 172350
rect 439742 172294 439838 172350
rect 439218 172226 439838 172294
rect 439218 172170 439314 172226
rect 439370 172170 439438 172226
rect 439494 172170 439562 172226
rect 439618 172170 439686 172226
rect 439742 172170 439838 172226
rect 439218 172102 439838 172170
rect 439218 172046 439314 172102
rect 439370 172046 439438 172102
rect 439494 172046 439562 172102
rect 439618 172046 439686 172102
rect 439742 172046 439838 172102
rect 439218 171978 439838 172046
rect 439218 171922 439314 171978
rect 439370 171922 439438 171978
rect 439494 171922 439562 171978
rect 439618 171922 439686 171978
rect 439742 171922 439838 171978
rect 439218 154350 439838 171922
rect 462812 173796 462868 173806
rect 461356 170436 461412 170446
rect 455308 165396 455364 165406
rect 439218 154294 439314 154350
rect 439370 154294 439438 154350
rect 439494 154294 439562 154350
rect 439618 154294 439686 154350
rect 439742 154294 439838 154350
rect 439218 154226 439838 154294
rect 439218 154170 439314 154226
rect 439370 154170 439438 154226
rect 439494 154170 439562 154226
rect 439618 154170 439686 154226
rect 439742 154170 439838 154226
rect 439218 154102 439838 154170
rect 439218 154046 439314 154102
rect 439370 154046 439438 154102
rect 439494 154046 439562 154102
rect 439618 154046 439686 154102
rect 439742 154046 439838 154102
rect 439218 153978 439838 154046
rect 439218 153922 439314 153978
rect 439370 153922 439438 153978
rect 439494 153922 439562 153978
rect 439618 153922 439686 153978
rect 439742 153922 439838 153978
rect 439218 136350 439838 153922
rect 452732 163156 452788 163166
rect 449372 148596 449428 148606
rect 449372 143780 449428 148540
rect 449372 143714 449428 143724
rect 452732 142100 452788 163100
rect 452732 142034 452788 142044
rect 455308 137788 455364 165340
rect 457772 162596 457828 162606
rect 456092 162036 456148 162046
rect 455308 137732 455700 137788
rect 439218 136294 439314 136350
rect 439370 136294 439438 136350
rect 439494 136294 439562 136350
rect 439618 136294 439686 136350
rect 439742 136294 439838 136350
rect 439218 136226 439838 136294
rect 439218 136170 439314 136226
rect 439370 136170 439438 136226
rect 439494 136170 439562 136226
rect 439618 136170 439686 136226
rect 439742 136170 439838 136226
rect 439218 136102 439838 136170
rect 439218 136046 439314 136102
rect 439370 136046 439438 136102
rect 439494 136046 439562 136102
rect 439618 136046 439686 136102
rect 439742 136046 439838 136102
rect 439218 135978 439838 136046
rect 439218 135922 439314 135978
rect 439370 135922 439438 135978
rect 439494 135922 439562 135978
rect 439618 135922 439686 135978
rect 439742 135922 439838 135978
rect 433808 118350 434128 118384
rect 433808 118294 433878 118350
rect 433934 118294 434002 118350
rect 434058 118294 434128 118350
rect 433808 118226 434128 118294
rect 433808 118170 433878 118226
rect 433934 118170 434002 118226
rect 434058 118170 434128 118226
rect 433808 118102 434128 118170
rect 433808 118046 433878 118102
rect 433934 118046 434002 118102
rect 434058 118046 434128 118102
rect 433808 117978 434128 118046
rect 433808 117922 433878 117978
rect 433934 117922 434002 117978
rect 434058 117922 434128 117978
rect 433808 117888 434128 117922
rect 439218 118350 439838 135922
rect 449168 130350 449488 130384
rect 449168 130294 449238 130350
rect 449294 130294 449362 130350
rect 449418 130294 449488 130350
rect 449168 130226 449488 130294
rect 449168 130170 449238 130226
rect 449294 130170 449362 130226
rect 449418 130170 449488 130226
rect 449168 130102 449488 130170
rect 449168 130046 449238 130102
rect 449294 130046 449362 130102
rect 449418 130046 449488 130102
rect 449168 129978 449488 130046
rect 449168 129922 449238 129978
rect 449294 129922 449362 129978
rect 449418 129922 449488 129978
rect 449168 129888 449488 129922
rect 455420 125758 455476 125768
rect 455420 125188 455476 125702
rect 455420 125122 455476 125132
rect 455308 123958 455364 123994
rect 455308 123890 455364 123900
rect 455308 120538 455364 120548
rect 455308 120372 455364 120482
rect 455308 120306 455364 120316
rect 439218 118294 439314 118350
rect 439370 118294 439438 118350
rect 439494 118294 439562 118350
rect 439618 118294 439686 118350
rect 439742 118294 439838 118350
rect 439218 118226 439838 118294
rect 439218 118170 439314 118226
rect 439370 118170 439438 118226
rect 439494 118170 439562 118226
rect 439618 118170 439686 118226
rect 439742 118170 439838 118226
rect 439218 118102 439838 118170
rect 439218 118046 439314 118102
rect 439370 118046 439438 118102
rect 439494 118046 439562 118102
rect 439618 118046 439686 118102
rect 439742 118046 439838 118102
rect 439218 117978 439838 118046
rect 439218 117922 439314 117978
rect 439370 117922 439438 117978
rect 439494 117922 439562 117978
rect 439618 117922 439686 117978
rect 439742 117922 439838 117978
rect 410844 116498 410900 116508
rect 418448 112350 418768 112384
rect 418448 112294 418518 112350
rect 418574 112294 418642 112350
rect 418698 112294 418768 112350
rect 418448 112226 418768 112294
rect 418448 112170 418518 112226
rect 418574 112170 418642 112226
rect 418698 112170 418768 112226
rect 418448 112102 418768 112170
rect 418448 112046 418518 112102
rect 418574 112046 418642 112102
rect 418698 112046 418768 112102
rect 418448 111978 418768 112046
rect 418448 111922 418518 111978
rect 418574 111922 418642 111978
rect 418698 111922 418768 111978
rect 418448 111888 418768 111922
rect 435498 112350 436118 114322
rect 435498 112294 435594 112350
rect 435650 112294 435718 112350
rect 435774 112294 435842 112350
rect 435898 112294 435966 112350
rect 436022 112294 436118 112350
rect 435498 112226 436118 112294
rect 435498 112170 435594 112226
rect 435650 112170 435718 112226
rect 435774 112170 435842 112226
rect 435898 112170 435966 112226
rect 436022 112170 436118 112226
rect 435498 112102 436118 112170
rect 435498 112046 435594 112102
rect 435650 112046 435718 112102
rect 435774 112046 435842 112102
rect 435898 112046 435966 112102
rect 436022 112046 436118 112102
rect 435498 111978 436118 112046
rect 435498 111922 435594 111978
rect 435650 111922 435718 111978
rect 435774 111922 435842 111978
rect 435898 111922 435966 111978
rect 436022 111922 436118 111978
rect 422044 102004 422100 102014
rect 408498 100294 408594 100350
rect 408650 100294 408718 100350
rect 408774 100294 408842 100350
rect 408898 100294 408966 100350
rect 409022 100294 409118 100350
rect 408498 100226 409118 100294
rect 408498 100170 408594 100226
rect 408650 100170 408718 100226
rect 408774 100170 408842 100226
rect 408898 100170 408966 100226
rect 409022 100170 409118 100226
rect 408498 100102 409118 100170
rect 408498 100046 408594 100102
rect 408650 100046 408718 100102
rect 408774 100046 408842 100102
rect 408898 100046 408966 100102
rect 409022 100046 409118 100102
rect 408498 99978 409118 100046
rect 408498 99922 408594 99978
rect 408650 99922 408718 99978
rect 408774 99922 408842 99978
rect 408898 99922 408966 99978
rect 409022 99922 409118 99978
rect 408498 82350 409118 99922
rect 408498 82294 408594 82350
rect 408650 82294 408718 82350
rect 408774 82294 408842 82350
rect 408898 82294 408966 82350
rect 409022 82294 409118 82350
rect 408498 82226 409118 82294
rect 408498 82170 408594 82226
rect 408650 82170 408718 82226
rect 408774 82170 408842 82226
rect 408898 82170 408966 82226
rect 409022 82170 409118 82226
rect 408498 82102 409118 82170
rect 408498 82046 408594 82102
rect 408650 82046 408718 82102
rect 408774 82046 408842 82102
rect 408898 82046 408966 82102
rect 409022 82046 409118 82102
rect 408498 81978 409118 82046
rect 408498 81922 408594 81978
rect 408650 81922 408718 81978
rect 408774 81922 408842 81978
rect 408898 81922 408966 81978
rect 409022 81922 409118 81978
rect 408498 64350 409118 81922
rect 411068 101668 411124 101678
rect 408498 64294 408594 64350
rect 408650 64294 408718 64350
rect 408774 64294 408842 64350
rect 408898 64294 408966 64350
rect 409022 64294 409118 64350
rect 408498 64226 409118 64294
rect 408498 64170 408594 64226
rect 408650 64170 408718 64226
rect 408774 64170 408842 64226
rect 408898 64170 408966 64226
rect 409022 64170 409118 64226
rect 408498 64102 409118 64170
rect 408498 64046 408594 64102
rect 408650 64046 408718 64102
rect 408774 64046 408842 64102
rect 408898 64046 408966 64102
rect 409022 64046 409118 64102
rect 408498 63978 409118 64046
rect 408498 63922 408594 63978
rect 408650 63922 408718 63978
rect 408774 63922 408842 63978
rect 408898 63922 408966 63978
rect 409022 63922 409118 63978
rect 408498 46350 409118 63922
rect 410732 73556 410788 73566
rect 410732 52164 410788 73500
rect 411068 55524 411124 101612
rect 422044 100772 422100 101948
rect 422044 100706 422100 100716
rect 429436 101892 429492 101902
rect 429436 100772 429492 101836
rect 429436 100706 429492 100716
rect 434140 101780 434196 101790
rect 434140 100772 434196 101724
rect 434140 100706 434196 100716
rect 435498 94350 436118 111922
rect 438844 101668 438900 101678
rect 438844 100772 438900 101612
rect 438844 100706 438900 100716
rect 435498 94294 435594 94350
rect 435650 94294 435718 94350
rect 435774 94294 435842 94350
rect 435898 94294 435966 94350
rect 436022 94294 436118 94350
rect 435498 94226 436118 94294
rect 435498 94170 435594 94226
rect 435650 94170 435718 94226
rect 435774 94170 435842 94226
rect 435898 94170 435966 94226
rect 436022 94170 436118 94226
rect 435498 94102 436118 94170
rect 435498 94046 435594 94102
rect 435650 94046 435718 94102
rect 435774 94046 435842 94102
rect 435898 94046 435966 94102
rect 436022 94046 436118 94102
rect 435498 93978 436118 94046
rect 435498 93922 435594 93978
rect 435650 93922 435718 93978
rect 435774 93922 435842 93978
rect 435898 93922 435966 93978
rect 436022 93922 436118 93978
rect 435498 76350 436118 93922
rect 435498 76294 435594 76350
rect 435650 76294 435718 76350
rect 435774 76294 435842 76350
rect 435898 76294 435966 76350
rect 436022 76294 436118 76350
rect 435498 76226 436118 76294
rect 435498 76170 435594 76226
rect 435650 76170 435718 76226
rect 435774 76170 435842 76226
rect 435898 76170 435966 76226
rect 436022 76170 436118 76226
rect 435498 76102 436118 76170
rect 435498 76046 435594 76102
rect 435650 76046 435718 76102
rect 435774 76046 435842 76102
rect 435898 76046 435966 76102
rect 436022 76046 436118 76102
rect 435498 75978 436118 76046
rect 435498 75922 435594 75978
rect 435650 75922 435718 75978
rect 435774 75922 435842 75978
rect 435898 75922 435966 75978
rect 436022 75922 436118 75978
rect 433808 64350 434128 64384
rect 433808 64294 433878 64350
rect 433934 64294 434002 64350
rect 434058 64294 434128 64350
rect 433808 64226 434128 64294
rect 433808 64170 433878 64226
rect 433934 64170 434002 64226
rect 434058 64170 434128 64226
rect 433808 64102 434128 64170
rect 433808 64046 433878 64102
rect 433934 64046 434002 64102
rect 434058 64046 434128 64102
rect 433808 63978 434128 64046
rect 433808 63922 433878 63978
rect 433934 63922 434002 63978
rect 434058 63922 434128 63978
rect 433808 63888 434128 63922
rect 418448 58350 418768 58384
rect 418448 58294 418518 58350
rect 418574 58294 418642 58350
rect 418698 58294 418768 58350
rect 418448 58226 418768 58294
rect 418448 58170 418518 58226
rect 418574 58170 418642 58226
rect 418698 58170 418768 58226
rect 418448 58102 418768 58170
rect 418448 58046 418518 58102
rect 418574 58046 418642 58102
rect 418698 58046 418768 58102
rect 418448 57978 418768 58046
rect 418448 57922 418518 57978
rect 418574 57922 418642 57978
rect 418698 57922 418768 57978
rect 418448 57888 418768 57922
rect 435498 58350 436118 75922
rect 435498 58294 435594 58350
rect 435650 58294 435718 58350
rect 435774 58294 435842 58350
rect 435898 58294 435966 58350
rect 436022 58294 436118 58350
rect 435498 58226 436118 58294
rect 435498 58170 435594 58226
rect 435650 58170 435718 58226
rect 435774 58170 435842 58226
rect 435898 58170 435966 58226
rect 436022 58170 436118 58226
rect 435498 58102 436118 58170
rect 435498 58046 435594 58102
rect 435650 58046 435718 58102
rect 435774 58046 435842 58102
rect 435898 58046 435966 58102
rect 436022 58046 436118 58102
rect 435498 57978 436118 58046
rect 435498 57922 435594 57978
rect 435650 57922 435718 57978
rect 435774 57922 435842 57978
rect 435898 57922 435966 57978
rect 436022 57922 436118 57978
rect 414652 56308 414708 56318
rect 414652 56212 414708 56222
rect 411068 55458 411124 55468
rect 435498 53694 436118 57922
rect 439218 100350 439838 117922
rect 455644 116564 455700 137732
rect 456092 119252 456148 161980
rect 456988 133498 457044 133508
rect 456988 120596 457044 133442
rect 457772 121156 457828 162540
rect 459004 157332 459060 157342
rect 458780 155652 458836 155662
rect 458780 121268 458836 155596
rect 458780 121202 458836 121212
rect 458892 142100 458948 142110
rect 457772 121090 457828 121100
rect 458668 121156 458724 121166
rect 456988 120530 457044 120540
rect 456092 119186 456148 119196
rect 458668 117236 458724 121100
rect 458892 117908 458948 142044
rect 459004 118580 459060 157276
rect 461356 119924 461412 170380
rect 462812 120148 462868 173740
rect 466218 166350 466838 183922
rect 466218 166294 466314 166350
rect 466370 166294 466438 166350
rect 466494 166294 466562 166350
rect 466618 166294 466686 166350
rect 466742 166294 466838 166350
rect 466218 166226 466838 166294
rect 466218 166170 466314 166226
rect 466370 166170 466438 166226
rect 466494 166170 466562 166226
rect 466618 166170 466686 166226
rect 466742 166170 466838 166226
rect 466218 166102 466838 166170
rect 466218 166046 466314 166102
rect 466370 166046 466438 166102
rect 466494 166046 466562 166102
rect 466618 166046 466686 166102
rect 466742 166046 466838 166102
rect 466218 165978 466838 166046
rect 466218 165922 466314 165978
rect 466370 165922 466438 165978
rect 466494 165922 466562 165978
rect 466618 165922 466686 165978
rect 466742 165922 466838 165978
rect 466218 148350 466838 165922
rect 466218 148294 466314 148350
rect 466370 148294 466438 148350
rect 466494 148294 466562 148350
rect 466618 148294 466686 148350
rect 466742 148294 466838 148350
rect 466218 148226 466838 148294
rect 466218 148170 466314 148226
rect 466370 148170 466438 148226
rect 466494 148170 466562 148226
rect 466618 148170 466686 148226
rect 466742 148170 466838 148226
rect 466218 148102 466838 148170
rect 466218 148046 466314 148102
rect 466370 148046 466438 148102
rect 466494 148046 466562 148102
rect 466618 148046 466686 148102
rect 466742 148046 466838 148102
rect 466218 147978 466838 148046
rect 466218 147922 466314 147978
rect 466370 147922 466438 147978
rect 466494 147922 466562 147978
rect 466618 147922 466686 147978
rect 466742 147922 466838 147978
rect 464492 140644 464548 140654
rect 464492 123956 464548 140588
rect 464492 123890 464548 123900
rect 466218 130350 466838 147922
rect 466218 130294 466314 130350
rect 466370 130294 466438 130350
rect 466494 130294 466562 130350
rect 466618 130294 466686 130350
rect 466742 130294 466838 130350
rect 466218 130226 466838 130294
rect 466218 130170 466314 130226
rect 466370 130170 466438 130226
rect 466494 130170 466562 130226
rect 466618 130170 466686 130226
rect 466742 130170 466838 130226
rect 466218 130102 466838 130170
rect 466218 130046 466314 130102
rect 466370 130046 466438 130102
rect 466494 130046 466562 130102
rect 466618 130046 466686 130102
rect 466742 130046 466838 130102
rect 466218 129978 466838 130046
rect 466218 129922 466314 129978
rect 466370 129922 466438 129978
rect 466494 129922 466562 129978
rect 466618 129922 466686 129978
rect 466742 129922 466838 129978
rect 462812 120082 462868 120092
rect 461356 119858 461412 119868
rect 459004 118514 459060 118524
rect 458892 117842 458948 117852
rect 458668 117170 458724 117180
rect 455644 116498 455700 116508
rect 449168 112350 449488 112384
rect 449168 112294 449238 112350
rect 449294 112294 449362 112350
rect 449418 112294 449488 112350
rect 449168 112226 449488 112294
rect 449168 112170 449238 112226
rect 449294 112170 449362 112226
rect 449418 112170 449488 112226
rect 449168 112102 449488 112170
rect 449168 112046 449238 112102
rect 449294 112046 449362 112102
rect 449418 112046 449488 112102
rect 449168 111978 449488 112046
rect 449168 111922 449238 111978
rect 449294 111922 449362 111978
rect 449418 111922 449488 111978
rect 449168 111888 449488 111922
rect 466218 112350 466838 129922
rect 466218 112294 466314 112350
rect 466370 112294 466438 112350
rect 466494 112294 466562 112350
rect 466618 112294 466686 112350
rect 466742 112294 466838 112350
rect 466218 112226 466838 112294
rect 466218 112170 466314 112226
rect 466370 112170 466438 112226
rect 466494 112170 466562 112226
rect 466618 112170 466686 112226
rect 466742 112170 466838 112226
rect 466218 112102 466838 112170
rect 466218 112046 466314 112102
rect 466370 112046 466438 112102
rect 466494 112046 466562 112102
rect 466618 112046 466686 112102
rect 466742 112046 466838 112102
rect 466218 111978 466838 112046
rect 466218 111922 466314 111978
rect 466370 111922 466438 111978
rect 466494 111922 466562 111978
rect 466618 111922 466686 111978
rect 466742 111922 466838 111978
rect 439218 100294 439314 100350
rect 439370 100294 439438 100350
rect 439494 100294 439562 100350
rect 439618 100294 439686 100350
rect 439742 100294 439838 100350
rect 439218 100226 439838 100294
rect 439218 100170 439314 100226
rect 439370 100170 439438 100226
rect 439494 100170 439562 100226
rect 439618 100170 439686 100226
rect 439742 100170 439838 100226
rect 439218 100102 439838 100170
rect 439218 100046 439314 100102
rect 439370 100046 439438 100102
rect 439494 100046 439562 100102
rect 439618 100046 439686 100102
rect 439742 100046 439838 100102
rect 439218 99978 439838 100046
rect 439218 99922 439314 99978
rect 439370 99922 439438 99978
rect 439494 99922 439562 99978
rect 439618 99922 439686 99978
rect 439742 99922 439838 99978
rect 439218 82350 439838 99922
rect 456988 99988 457044 99998
rect 439218 82294 439314 82350
rect 439370 82294 439438 82350
rect 439494 82294 439562 82350
rect 439618 82294 439686 82350
rect 439742 82294 439838 82350
rect 439218 82226 439838 82294
rect 439218 82170 439314 82226
rect 439370 82170 439438 82226
rect 439494 82170 439562 82226
rect 439618 82170 439686 82226
rect 439742 82170 439838 82226
rect 439218 82102 439838 82170
rect 439218 82046 439314 82102
rect 439370 82046 439438 82102
rect 439494 82046 439562 82102
rect 439618 82046 439686 82102
rect 439742 82046 439838 82102
rect 439218 81978 439838 82046
rect 439218 81922 439314 81978
rect 439370 81922 439438 81978
rect 439494 81922 439562 81978
rect 439618 81922 439686 81978
rect 439742 81922 439838 81978
rect 439218 64350 439838 81922
rect 439218 64294 439314 64350
rect 439370 64294 439438 64350
rect 439494 64294 439562 64350
rect 439618 64294 439686 64350
rect 439742 64294 439838 64350
rect 439218 64226 439838 64294
rect 439218 64170 439314 64226
rect 439370 64170 439438 64226
rect 439494 64170 439562 64226
rect 439618 64170 439686 64226
rect 439742 64170 439838 64226
rect 439218 64102 439838 64170
rect 439218 64046 439314 64102
rect 439370 64046 439438 64102
rect 439494 64046 439562 64102
rect 439618 64046 439686 64102
rect 439742 64046 439838 64102
rect 439218 63978 439838 64046
rect 439218 63922 439314 63978
rect 439370 63922 439438 63978
rect 439494 63922 439562 63978
rect 439618 63922 439686 63978
rect 439742 63922 439838 63978
rect 410732 52098 410788 52108
rect 408498 46294 408594 46350
rect 408650 46294 408718 46350
rect 408774 46294 408842 46350
rect 408898 46294 408966 46350
rect 409022 46294 409118 46350
rect 408498 46226 409118 46294
rect 408498 46170 408594 46226
rect 408650 46170 408718 46226
rect 408774 46170 408842 46226
rect 408898 46170 408966 46226
rect 409022 46170 409118 46226
rect 408498 46102 409118 46170
rect 408498 46046 408594 46102
rect 408650 46046 408718 46102
rect 408774 46046 408842 46102
rect 408898 46046 408966 46102
rect 409022 46046 409118 46102
rect 408498 45978 409118 46046
rect 408498 45922 408594 45978
rect 408650 45922 408718 45978
rect 408774 45922 408842 45978
rect 408898 45922 408966 45978
rect 409022 45922 409118 45978
rect 408498 28350 409118 45922
rect 433808 46350 434128 46384
rect 433808 46294 433878 46350
rect 433934 46294 434002 46350
rect 434058 46294 434128 46350
rect 433808 46226 434128 46294
rect 433808 46170 433878 46226
rect 433934 46170 434002 46226
rect 434058 46170 434128 46226
rect 433808 46102 434128 46170
rect 433808 46046 433878 46102
rect 433934 46046 434002 46102
rect 434058 46046 434128 46102
rect 433808 45978 434128 46046
rect 433808 45922 433878 45978
rect 433934 45922 434002 45978
rect 434058 45922 434128 45978
rect 433808 45888 434128 45922
rect 439218 46350 439838 63922
rect 455308 95060 455364 95070
rect 449168 58350 449488 58384
rect 449168 58294 449238 58350
rect 449294 58294 449362 58350
rect 449418 58294 449488 58350
rect 449168 58226 449488 58294
rect 449168 58170 449238 58226
rect 449294 58170 449362 58226
rect 449418 58170 449488 58226
rect 449168 58102 449488 58170
rect 449168 58046 449238 58102
rect 449294 58046 449362 58102
rect 449418 58046 449488 58102
rect 449168 57978 449488 58046
rect 449168 57922 449238 57978
rect 449294 57922 449362 57978
rect 449418 57922 449488 57978
rect 449168 57888 449488 57922
rect 455308 53508 455364 95004
rect 455308 53442 455364 53452
rect 455420 73444 455476 73454
rect 455420 48132 455476 73388
rect 455420 48066 455476 48076
rect 456092 72996 456148 73006
rect 456092 47572 456148 72940
rect 456988 51492 457044 99932
rect 466218 94350 466838 111922
rect 466218 94294 466314 94350
rect 466370 94294 466438 94350
rect 466494 94294 466562 94350
rect 466618 94294 466686 94350
rect 466742 94294 466838 94350
rect 466218 94226 466838 94294
rect 466218 94170 466314 94226
rect 466370 94170 466438 94226
rect 466494 94170 466562 94226
rect 466618 94170 466686 94226
rect 466742 94170 466838 94226
rect 466218 94102 466838 94170
rect 466218 94046 466314 94102
rect 466370 94046 466438 94102
rect 466494 94046 466562 94102
rect 466618 94046 466686 94102
rect 466742 94046 466838 94102
rect 466218 93978 466838 94046
rect 466218 93922 466314 93978
rect 466370 93922 466438 93978
rect 466494 93922 466562 93978
rect 466618 93922 466686 93978
rect 466742 93922 466838 93978
rect 458668 88340 458724 88350
rect 457100 84980 457156 84990
rect 457100 55524 457156 84924
rect 457772 76916 457828 76926
rect 457100 55458 457156 55468
rect 457212 71652 457268 71662
rect 456988 51426 457044 51436
rect 457212 50820 457268 71596
rect 457772 52948 457828 76860
rect 458668 54852 458724 88284
rect 458668 54786 458724 54796
rect 458780 86660 458836 86670
rect 458780 54180 458836 86604
rect 462812 84196 462868 84206
rect 458780 54114 458836 54124
rect 458892 79940 458948 79950
rect 457772 52882 457828 52892
rect 457212 50754 457268 50764
rect 458892 50148 458948 79884
rect 459116 71764 459172 71774
rect 458892 50082 458948 50092
rect 459004 68292 459060 68302
rect 459004 49476 459060 68236
rect 459116 53284 459172 71708
rect 459116 53218 459172 53228
rect 462812 52836 462868 84140
rect 462812 52770 462868 52780
rect 466218 76350 466838 93922
rect 466218 76294 466314 76350
rect 466370 76294 466438 76350
rect 466494 76294 466562 76350
rect 466618 76294 466686 76350
rect 466742 76294 466838 76350
rect 466218 76226 466838 76294
rect 466218 76170 466314 76226
rect 466370 76170 466438 76226
rect 466494 76170 466562 76226
rect 466618 76170 466686 76226
rect 466742 76170 466838 76226
rect 466218 76102 466838 76170
rect 466218 76046 466314 76102
rect 466370 76046 466438 76102
rect 466494 76046 466562 76102
rect 466618 76046 466686 76102
rect 466742 76046 466838 76102
rect 466218 75978 466838 76046
rect 466218 75922 466314 75978
rect 466370 75922 466438 75978
rect 466494 75922 466562 75978
rect 466618 75922 466686 75978
rect 466742 75922 466838 75978
rect 466218 58350 466838 75922
rect 466218 58294 466314 58350
rect 466370 58294 466438 58350
rect 466494 58294 466562 58350
rect 466618 58294 466686 58350
rect 466742 58294 466838 58350
rect 466218 58226 466838 58294
rect 466218 58170 466314 58226
rect 466370 58170 466438 58226
rect 466494 58170 466562 58226
rect 466618 58170 466686 58226
rect 466742 58170 466838 58226
rect 466218 58102 466838 58170
rect 466218 58046 466314 58102
rect 466370 58046 466438 58102
rect 466494 58046 466562 58102
rect 466618 58046 466686 58102
rect 466742 58046 466838 58102
rect 466218 57978 466838 58046
rect 466218 57922 466314 57978
rect 466370 57922 466438 57978
rect 466494 57922 466562 57978
rect 466618 57922 466686 57978
rect 466742 57922 466838 57978
rect 459004 49410 459060 49420
rect 456092 47506 456148 47516
rect 439218 46294 439314 46350
rect 439370 46294 439438 46350
rect 439494 46294 439562 46350
rect 439618 46294 439686 46350
rect 439742 46294 439838 46350
rect 439218 46226 439838 46294
rect 439218 46170 439314 46226
rect 439370 46170 439438 46226
rect 439494 46170 439562 46226
rect 439618 46170 439686 46226
rect 439742 46170 439838 46226
rect 439218 46102 439838 46170
rect 439218 46046 439314 46102
rect 439370 46046 439438 46102
rect 439494 46046 439562 46102
rect 439618 46046 439686 46102
rect 439742 46046 439838 46102
rect 439218 45978 439838 46046
rect 439218 45922 439314 45978
rect 439370 45922 439438 45978
rect 439494 45922 439562 45978
rect 439618 45922 439686 45978
rect 439742 45922 439838 45978
rect 418448 40350 418768 40384
rect 418448 40294 418518 40350
rect 418574 40294 418642 40350
rect 418698 40294 418768 40350
rect 418448 40226 418768 40294
rect 418448 40170 418518 40226
rect 418574 40170 418642 40226
rect 418698 40170 418768 40226
rect 418448 40102 418768 40170
rect 418448 40046 418518 40102
rect 418574 40046 418642 40102
rect 418698 40046 418768 40102
rect 418448 39978 418768 40046
rect 418448 39922 418518 39978
rect 418574 39922 418642 39978
rect 418698 39922 418768 39978
rect 418448 39888 418768 39922
rect 435498 40350 436118 45698
rect 435498 40294 435594 40350
rect 435650 40294 435718 40350
rect 435774 40294 435842 40350
rect 435898 40294 435966 40350
rect 436022 40294 436118 40350
rect 435498 40226 436118 40294
rect 435498 40170 435594 40226
rect 435650 40170 435718 40226
rect 435774 40170 435842 40226
rect 435898 40170 435966 40226
rect 436022 40170 436118 40226
rect 435498 40102 436118 40170
rect 435498 40046 435594 40102
rect 435650 40046 435718 40102
rect 435774 40046 435842 40102
rect 435898 40046 435966 40102
rect 436022 40046 436118 40102
rect 435498 39978 436118 40046
rect 435498 39922 435594 39978
rect 435650 39922 435718 39978
rect 435774 39922 435842 39978
rect 435898 39922 435966 39978
rect 436022 39922 436118 39978
rect 408498 28294 408594 28350
rect 408650 28294 408718 28350
rect 408774 28294 408842 28350
rect 408898 28294 408966 28350
rect 409022 28294 409118 28350
rect 408498 28226 409118 28294
rect 408498 28170 408594 28226
rect 408650 28170 408718 28226
rect 408774 28170 408842 28226
rect 408898 28170 408966 28226
rect 409022 28170 409118 28226
rect 408498 28102 409118 28170
rect 408498 28046 408594 28102
rect 408650 28046 408718 28102
rect 408774 28046 408842 28102
rect 408898 28046 408966 28102
rect 409022 28046 409118 28102
rect 408498 27978 409118 28046
rect 408498 27922 408594 27978
rect 408650 27922 408718 27978
rect 408774 27922 408842 27978
rect 408898 27922 408966 27978
rect 409022 27922 409118 27978
rect 408498 10350 409118 27922
rect 408498 10294 408594 10350
rect 408650 10294 408718 10350
rect 408774 10294 408842 10350
rect 408898 10294 408966 10350
rect 409022 10294 409118 10350
rect 408498 10226 409118 10294
rect 408498 10170 408594 10226
rect 408650 10170 408718 10226
rect 408774 10170 408842 10226
rect 408898 10170 408966 10226
rect 409022 10170 409118 10226
rect 408498 10102 409118 10170
rect 408498 10046 408594 10102
rect 408650 10046 408718 10102
rect 408774 10046 408842 10102
rect 408898 10046 408966 10102
rect 409022 10046 409118 10102
rect 408498 9978 409118 10046
rect 408498 9922 408594 9978
rect 408650 9922 408718 9978
rect 408774 9922 408842 9978
rect 408898 9922 408966 9978
rect 409022 9922 409118 9978
rect 408498 -1120 409118 9922
rect 408498 -1176 408594 -1120
rect 408650 -1176 408718 -1120
rect 408774 -1176 408842 -1120
rect 408898 -1176 408966 -1120
rect 409022 -1176 409118 -1120
rect 408498 -1244 409118 -1176
rect 408498 -1300 408594 -1244
rect 408650 -1300 408718 -1244
rect 408774 -1300 408842 -1244
rect 408898 -1300 408966 -1244
rect 409022 -1300 409118 -1244
rect 408498 -1368 409118 -1300
rect 408498 -1424 408594 -1368
rect 408650 -1424 408718 -1368
rect 408774 -1424 408842 -1368
rect 408898 -1424 408966 -1368
rect 409022 -1424 409118 -1368
rect 408498 -1492 409118 -1424
rect 408498 -1548 408594 -1492
rect 408650 -1548 408718 -1492
rect 408774 -1548 408842 -1492
rect 408898 -1548 408966 -1492
rect 409022 -1548 409118 -1492
rect 408498 -1644 409118 -1548
rect 435498 22350 436118 39922
rect 435498 22294 435594 22350
rect 435650 22294 435718 22350
rect 435774 22294 435842 22350
rect 435898 22294 435966 22350
rect 436022 22294 436118 22350
rect 435498 22226 436118 22294
rect 435498 22170 435594 22226
rect 435650 22170 435718 22226
rect 435774 22170 435842 22226
rect 435898 22170 435966 22226
rect 436022 22170 436118 22226
rect 435498 22102 436118 22170
rect 435498 22046 435594 22102
rect 435650 22046 435718 22102
rect 435774 22046 435842 22102
rect 435898 22046 435966 22102
rect 436022 22046 436118 22102
rect 435498 21978 436118 22046
rect 435498 21922 435594 21978
rect 435650 21922 435718 21978
rect 435774 21922 435842 21978
rect 435898 21922 435966 21978
rect 436022 21922 436118 21978
rect 435498 4350 436118 21922
rect 435498 4294 435594 4350
rect 435650 4294 435718 4350
rect 435774 4294 435842 4350
rect 435898 4294 435966 4350
rect 436022 4294 436118 4350
rect 435498 4226 436118 4294
rect 435498 4170 435594 4226
rect 435650 4170 435718 4226
rect 435774 4170 435842 4226
rect 435898 4170 435966 4226
rect 436022 4170 436118 4226
rect 435498 4102 436118 4170
rect 435498 4046 435594 4102
rect 435650 4046 435718 4102
rect 435774 4046 435842 4102
rect 435898 4046 435966 4102
rect 436022 4046 436118 4102
rect 435498 3978 436118 4046
rect 435498 3922 435594 3978
rect 435650 3922 435718 3978
rect 435774 3922 435842 3978
rect 435898 3922 435966 3978
rect 436022 3922 436118 3978
rect 435498 -160 436118 3922
rect 435498 -216 435594 -160
rect 435650 -216 435718 -160
rect 435774 -216 435842 -160
rect 435898 -216 435966 -160
rect 436022 -216 436118 -160
rect 435498 -284 436118 -216
rect 435498 -340 435594 -284
rect 435650 -340 435718 -284
rect 435774 -340 435842 -284
rect 435898 -340 435966 -284
rect 436022 -340 436118 -284
rect 435498 -408 436118 -340
rect 435498 -464 435594 -408
rect 435650 -464 435718 -408
rect 435774 -464 435842 -408
rect 435898 -464 435966 -408
rect 436022 -464 436118 -408
rect 435498 -532 436118 -464
rect 435498 -588 435594 -532
rect 435650 -588 435718 -532
rect 435774 -588 435842 -532
rect 435898 -588 435966 -532
rect 436022 -588 436118 -532
rect 435498 -1644 436118 -588
rect 439218 28350 439838 45922
rect 449168 40350 449488 40384
rect 449168 40294 449238 40350
rect 449294 40294 449362 40350
rect 449418 40294 449488 40350
rect 449168 40226 449488 40294
rect 449168 40170 449238 40226
rect 449294 40170 449362 40226
rect 449418 40170 449488 40226
rect 449168 40102 449488 40170
rect 449168 40046 449238 40102
rect 449294 40046 449362 40102
rect 449418 40046 449488 40102
rect 449168 39978 449488 40046
rect 449168 39922 449238 39978
rect 449294 39922 449362 39978
rect 449418 39922 449488 39978
rect 449168 39888 449488 39922
rect 466218 40350 466838 57922
rect 466218 40294 466314 40350
rect 466370 40294 466438 40350
rect 466494 40294 466562 40350
rect 466618 40294 466686 40350
rect 466742 40294 466838 40350
rect 466218 40226 466838 40294
rect 466218 40170 466314 40226
rect 466370 40170 466438 40226
rect 466494 40170 466562 40226
rect 466618 40170 466686 40226
rect 466742 40170 466838 40226
rect 466218 40102 466838 40170
rect 466218 40046 466314 40102
rect 466370 40046 466438 40102
rect 466494 40046 466562 40102
rect 466618 40046 466686 40102
rect 466742 40046 466838 40102
rect 466218 39978 466838 40046
rect 466218 39922 466314 39978
rect 466370 39922 466438 39978
rect 466494 39922 466562 39978
rect 466618 39922 466686 39978
rect 466742 39922 466838 39978
rect 439218 28294 439314 28350
rect 439370 28294 439438 28350
rect 439494 28294 439562 28350
rect 439618 28294 439686 28350
rect 439742 28294 439838 28350
rect 439218 28226 439838 28294
rect 439218 28170 439314 28226
rect 439370 28170 439438 28226
rect 439494 28170 439562 28226
rect 439618 28170 439686 28226
rect 439742 28170 439838 28226
rect 439218 28102 439838 28170
rect 439218 28046 439314 28102
rect 439370 28046 439438 28102
rect 439494 28046 439562 28102
rect 439618 28046 439686 28102
rect 439742 28046 439838 28102
rect 439218 27978 439838 28046
rect 439218 27922 439314 27978
rect 439370 27922 439438 27978
rect 439494 27922 439562 27978
rect 439618 27922 439686 27978
rect 439742 27922 439838 27978
rect 439218 10350 439838 27922
rect 439218 10294 439314 10350
rect 439370 10294 439438 10350
rect 439494 10294 439562 10350
rect 439618 10294 439686 10350
rect 439742 10294 439838 10350
rect 439218 10226 439838 10294
rect 439218 10170 439314 10226
rect 439370 10170 439438 10226
rect 439494 10170 439562 10226
rect 439618 10170 439686 10226
rect 439742 10170 439838 10226
rect 439218 10102 439838 10170
rect 439218 10046 439314 10102
rect 439370 10046 439438 10102
rect 439494 10046 439562 10102
rect 439618 10046 439686 10102
rect 439742 10046 439838 10102
rect 439218 9978 439838 10046
rect 439218 9922 439314 9978
rect 439370 9922 439438 9978
rect 439494 9922 439562 9978
rect 439618 9922 439686 9978
rect 439742 9922 439838 9978
rect 439218 -1120 439838 9922
rect 439218 -1176 439314 -1120
rect 439370 -1176 439438 -1120
rect 439494 -1176 439562 -1120
rect 439618 -1176 439686 -1120
rect 439742 -1176 439838 -1120
rect 439218 -1244 439838 -1176
rect 439218 -1300 439314 -1244
rect 439370 -1300 439438 -1244
rect 439494 -1300 439562 -1244
rect 439618 -1300 439686 -1244
rect 439742 -1300 439838 -1244
rect 439218 -1368 439838 -1300
rect 439218 -1424 439314 -1368
rect 439370 -1424 439438 -1368
rect 439494 -1424 439562 -1368
rect 439618 -1424 439686 -1368
rect 439742 -1424 439838 -1368
rect 439218 -1492 439838 -1424
rect 439218 -1548 439314 -1492
rect 439370 -1548 439438 -1492
rect 439494 -1548 439562 -1492
rect 439618 -1548 439686 -1492
rect 439742 -1548 439838 -1492
rect 439218 -1644 439838 -1548
rect 466218 22350 466838 39922
rect 466218 22294 466314 22350
rect 466370 22294 466438 22350
rect 466494 22294 466562 22350
rect 466618 22294 466686 22350
rect 466742 22294 466838 22350
rect 466218 22226 466838 22294
rect 466218 22170 466314 22226
rect 466370 22170 466438 22226
rect 466494 22170 466562 22226
rect 466618 22170 466686 22226
rect 466742 22170 466838 22226
rect 466218 22102 466838 22170
rect 466218 22046 466314 22102
rect 466370 22046 466438 22102
rect 466494 22046 466562 22102
rect 466618 22046 466686 22102
rect 466742 22046 466838 22102
rect 466218 21978 466838 22046
rect 466218 21922 466314 21978
rect 466370 21922 466438 21978
rect 466494 21922 466562 21978
rect 466618 21922 466686 21978
rect 466742 21922 466838 21978
rect 466218 4350 466838 21922
rect 466218 4294 466314 4350
rect 466370 4294 466438 4350
rect 466494 4294 466562 4350
rect 466618 4294 466686 4350
rect 466742 4294 466838 4350
rect 466218 4226 466838 4294
rect 466218 4170 466314 4226
rect 466370 4170 466438 4226
rect 466494 4170 466562 4226
rect 466618 4170 466686 4226
rect 466742 4170 466838 4226
rect 466218 4102 466838 4170
rect 466218 4046 466314 4102
rect 466370 4046 466438 4102
rect 466494 4046 466562 4102
rect 466618 4046 466686 4102
rect 466742 4046 466838 4102
rect 466218 3978 466838 4046
rect 466218 3922 466314 3978
rect 466370 3922 466438 3978
rect 466494 3922 466562 3978
rect 466618 3922 466686 3978
rect 466742 3922 466838 3978
rect 466218 -160 466838 3922
rect 466218 -216 466314 -160
rect 466370 -216 466438 -160
rect 466494 -216 466562 -160
rect 466618 -216 466686 -160
rect 466742 -216 466838 -160
rect 466218 -284 466838 -216
rect 466218 -340 466314 -284
rect 466370 -340 466438 -284
rect 466494 -340 466562 -284
rect 466618 -340 466686 -284
rect 466742 -340 466838 -284
rect 466218 -408 466838 -340
rect 466218 -464 466314 -408
rect 466370 -464 466438 -408
rect 466494 -464 466562 -408
rect 466618 -464 466686 -408
rect 466742 -464 466838 -408
rect 466218 -532 466838 -464
rect 466218 -588 466314 -532
rect 466370 -588 466438 -532
rect 466494 -588 466562 -532
rect 466618 -588 466686 -532
rect 466742 -588 466838 -532
rect 466218 -1644 466838 -588
rect 469938 190350 470558 207922
rect 495808 208350 496128 208384
rect 495808 208294 495878 208350
rect 495934 208294 496002 208350
rect 496058 208294 496128 208350
rect 495808 208226 496128 208294
rect 495808 208170 495878 208226
rect 495934 208170 496002 208226
rect 496058 208170 496128 208226
rect 495808 208102 496128 208170
rect 495808 208046 495878 208102
rect 495934 208046 496002 208102
rect 496058 208046 496128 208102
rect 495808 207978 496128 208046
rect 495808 207922 495878 207978
rect 495934 207922 496002 207978
rect 496058 207922 496128 207978
rect 495808 207888 496128 207922
rect 480448 202350 480768 202384
rect 480448 202294 480518 202350
rect 480574 202294 480642 202350
rect 480698 202294 480768 202350
rect 480448 202226 480768 202294
rect 480448 202170 480518 202226
rect 480574 202170 480642 202226
rect 480698 202170 480768 202226
rect 480448 202102 480768 202170
rect 480448 202046 480518 202102
rect 480574 202046 480642 202102
rect 480698 202046 480768 202102
rect 480448 201978 480768 202046
rect 480448 201922 480518 201978
rect 480574 201922 480642 201978
rect 480698 201922 480768 201978
rect 480448 201888 480768 201922
rect 496938 202350 497558 219922
rect 496938 202294 497034 202350
rect 497090 202294 497158 202350
rect 497214 202294 497282 202350
rect 497338 202294 497406 202350
rect 497462 202294 497558 202350
rect 496938 202226 497558 202294
rect 496938 202170 497034 202226
rect 497090 202170 497158 202226
rect 497214 202170 497282 202226
rect 497338 202170 497406 202226
rect 497462 202170 497558 202226
rect 496938 202102 497558 202170
rect 496938 202046 497034 202102
rect 497090 202046 497158 202102
rect 497214 202046 497282 202102
rect 497338 202046 497406 202102
rect 497462 202046 497558 202102
rect 496938 201978 497558 202046
rect 496938 201922 497034 201978
rect 497090 201922 497158 201978
rect 497214 201922 497282 201978
rect 497338 201922 497406 201978
rect 497462 201922 497558 201978
rect 473676 198298 473732 198308
rect 473676 197876 473732 198242
rect 473676 197810 473732 197820
rect 472108 195778 472164 195788
rect 472108 193844 472164 195722
rect 472108 193778 472164 193788
rect 472108 192388 472164 192398
rect 472108 191156 472164 192332
rect 472108 191090 472164 191100
rect 469938 190294 470034 190350
rect 470090 190294 470158 190350
rect 470214 190294 470282 190350
rect 470338 190294 470406 190350
rect 470462 190294 470558 190350
rect 469938 190226 470558 190294
rect 469938 190170 470034 190226
rect 470090 190170 470158 190226
rect 470214 190170 470282 190226
rect 470338 190170 470406 190226
rect 470462 190170 470558 190226
rect 469938 190102 470558 190170
rect 469938 190046 470034 190102
rect 470090 190046 470158 190102
rect 470214 190046 470282 190102
rect 470338 190046 470406 190102
rect 470462 190046 470558 190102
rect 469938 189978 470558 190046
rect 469938 189922 470034 189978
rect 470090 189922 470158 189978
rect 470214 189922 470282 189978
rect 470338 189922 470406 189978
rect 470462 189922 470558 189978
rect 469938 172350 470558 189922
rect 495808 190350 496128 190384
rect 495808 190294 495878 190350
rect 495934 190294 496002 190350
rect 496058 190294 496128 190350
rect 495808 190226 496128 190294
rect 495808 190170 495878 190226
rect 495934 190170 496002 190226
rect 496058 190170 496128 190226
rect 495808 190102 496128 190170
rect 495808 190046 495878 190102
rect 495934 190046 496002 190102
rect 496058 190046 496128 190102
rect 495808 189978 496128 190046
rect 495808 189922 495878 189978
rect 495934 189922 496002 189978
rect 496058 189922 496128 189978
rect 495808 189888 496128 189922
rect 472108 189812 472164 189822
rect 472108 189658 472164 189756
rect 472108 189592 472164 189602
rect 472108 188038 472164 188048
rect 472108 187124 472164 187982
rect 472108 187058 472164 187068
rect 480448 184350 480768 184384
rect 480448 184294 480518 184350
rect 480574 184294 480642 184350
rect 480698 184294 480768 184350
rect 480448 184226 480768 184294
rect 480448 184170 480518 184226
rect 480574 184170 480642 184226
rect 480698 184170 480768 184226
rect 480448 184102 480768 184170
rect 480448 184046 480518 184102
rect 480574 184046 480642 184102
rect 480698 184046 480768 184102
rect 480448 183978 480768 184046
rect 480448 183922 480518 183978
rect 480574 183922 480642 183978
rect 480698 183922 480768 183978
rect 480448 183888 480768 183922
rect 496938 184350 497558 201922
rect 496938 184294 497034 184350
rect 497090 184294 497158 184350
rect 497214 184294 497282 184350
rect 497338 184294 497406 184350
rect 497462 184294 497558 184350
rect 496938 184226 497558 184294
rect 496938 184170 497034 184226
rect 497090 184170 497158 184226
rect 497214 184170 497282 184226
rect 497338 184170 497406 184226
rect 497462 184170 497558 184226
rect 496938 184102 497558 184170
rect 496938 184046 497034 184102
rect 497090 184046 497158 184102
rect 497214 184046 497282 184102
rect 497338 184046 497406 184102
rect 497462 184046 497558 184102
rect 496938 183978 497558 184046
rect 496938 183922 497034 183978
rect 497090 183922 497158 183978
rect 497214 183922 497282 183978
rect 497338 183922 497406 183978
rect 497462 183922 497558 183978
rect 469938 172294 470034 172350
rect 470090 172294 470158 172350
rect 470214 172294 470282 172350
rect 470338 172294 470406 172350
rect 470462 172294 470558 172350
rect 469938 172226 470558 172294
rect 469938 172170 470034 172226
rect 470090 172170 470158 172226
rect 470214 172170 470282 172226
rect 470338 172170 470406 172226
rect 470462 172170 470558 172226
rect 469938 172102 470558 172170
rect 469938 172046 470034 172102
rect 470090 172046 470158 172102
rect 470214 172046 470282 172102
rect 470338 172046 470406 172102
rect 470462 172046 470558 172102
rect 469938 171978 470558 172046
rect 469938 171922 470034 171978
rect 470090 171922 470158 171978
rect 470214 171922 470282 171978
rect 470338 171922 470406 171978
rect 470462 171922 470558 171978
rect 469938 154350 470558 171922
rect 469938 154294 470034 154350
rect 470090 154294 470158 154350
rect 470214 154294 470282 154350
rect 470338 154294 470406 154350
rect 470462 154294 470558 154350
rect 469938 154226 470558 154294
rect 469938 154170 470034 154226
rect 470090 154170 470158 154226
rect 470214 154170 470282 154226
rect 470338 154170 470406 154226
rect 470462 154170 470558 154226
rect 469938 154102 470558 154170
rect 469938 154046 470034 154102
rect 470090 154046 470158 154102
rect 470214 154046 470282 154102
rect 470338 154046 470406 154102
rect 470462 154046 470558 154102
rect 469938 153978 470558 154046
rect 469938 153922 470034 153978
rect 470090 153922 470158 153978
rect 470214 153922 470282 153978
rect 470338 153922 470406 153978
rect 470462 153922 470558 153978
rect 469938 136350 470558 153922
rect 496938 166350 497558 183922
rect 496938 166294 497034 166350
rect 497090 166294 497158 166350
rect 497214 166294 497282 166350
rect 497338 166294 497406 166350
rect 497462 166294 497558 166350
rect 496938 166226 497558 166294
rect 496938 166170 497034 166226
rect 497090 166170 497158 166226
rect 497214 166170 497282 166226
rect 497338 166170 497406 166226
rect 497462 166170 497558 166226
rect 496938 166102 497558 166170
rect 496938 166046 497034 166102
rect 497090 166046 497158 166102
rect 497214 166046 497282 166102
rect 497338 166046 497406 166102
rect 497462 166046 497558 166102
rect 496938 165978 497558 166046
rect 496938 165922 497034 165978
rect 497090 165922 497158 165978
rect 497214 165922 497282 165978
rect 497338 165922 497406 165978
rect 497462 165922 497558 165978
rect 473004 152180 473060 152190
rect 469938 136294 470034 136350
rect 470090 136294 470158 136350
rect 470214 136294 470282 136350
rect 470338 136294 470406 136350
rect 470462 136294 470558 136350
rect 469938 136226 470558 136294
rect 469938 136170 470034 136226
rect 470090 136170 470158 136226
rect 470214 136170 470282 136226
rect 470338 136170 470406 136226
rect 470462 136170 470558 136226
rect 469938 136102 470558 136170
rect 469938 136046 470034 136102
rect 470090 136046 470158 136102
rect 470214 136046 470282 136102
rect 470338 136046 470406 136102
rect 470462 136046 470558 136102
rect 469938 135978 470558 136046
rect 469938 135922 470034 135978
rect 470090 135922 470158 135978
rect 470214 135922 470282 135978
rect 470338 135922 470406 135978
rect 470462 135922 470558 135978
rect 469938 118350 470558 135922
rect 472892 143668 472948 143678
rect 469938 118294 470034 118350
rect 470090 118294 470158 118350
rect 470214 118294 470282 118350
rect 470338 118294 470406 118350
rect 470462 118294 470558 118350
rect 469938 118226 470558 118294
rect 469938 118170 470034 118226
rect 470090 118170 470158 118226
rect 470214 118170 470282 118226
rect 470338 118170 470406 118226
rect 470462 118170 470558 118226
rect 469938 118102 470558 118170
rect 469938 118046 470034 118102
rect 470090 118046 470158 118102
rect 470214 118046 470282 118102
rect 470338 118046 470406 118102
rect 470462 118046 470558 118102
rect 469938 117978 470558 118046
rect 469938 117922 470034 117978
rect 470090 117922 470158 117978
rect 470214 117922 470282 117978
rect 470338 117922 470406 117978
rect 470462 117922 470558 117978
rect 469938 100350 470558 117922
rect 472108 120148 472164 120158
rect 472108 117908 472164 120092
rect 472108 117842 472164 117852
rect 472892 117236 472948 143612
rect 473004 126644 473060 152124
rect 496938 148350 497558 165922
rect 496938 148294 497034 148350
rect 497090 148294 497158 148350
rect 497214 148294 497282 148350
rect 497338 148294 497406 148350
rect 497462 148294 497558 148350
rect 496938 148226 497558 148294
rect 496938 148170 497034 148226
rect 497090 148170 497158 148226
rect 497214 148170 497282 148226
rect 497338 148170 497406 148226
rect 497462 148170 497558 148226
rect 496938 148102 497558 148170
rect 496938 148046 497034 148102
rect 497090 148046 497158 148102
rect 497214 148046 497282 148102
rect 497338 148046 497406 148102
rect 497462 148046 497558 148102
rect 496938 147978 497558 148046
rect 496938 147922 497034 147978
rect 497090 147922 497158 147978
rect 497214 147922 497282 147978
rect 497338 147922 497406 147978
rect 497462 147922 497558 147978
rect 495808 136350 496128 136384
rect 495808 136294 495878 136350
rect 495934 136294 496002 136350
rect 496058 136294 496128 136350
rect 495808 136226 496128 136294
rect 495808 136170 495878 136226
rect 495934 136170 496002 136226
rect 496058 136170 496128 136226
rect 495808 136102 496128 136170
rect 495808 136046 495878 136102
rect 495934 136046 496002 136102
rect 496058 136046 496128 136102
rect 495808 135978 496128 136046
rect 495808 135922 495878 135978
rect 495934 135922 496002 135978
rect 496058 135922 496128 135978
rect 495808 135888 496128 135922
rect 480448 130350 480768 130384
rect 480448 130294 480518 130350
rect 480574 130294 480642 130350
rect 480698 130294 480768 130350
rect 480448 130226 480768 130294
rect 480448 130170 480518 130226
rect 480574 130170 480642 130226
rect 480698 130170 480768 130226
rect 480448 130102 480768 130170
rect 480448 130046 480518 130102
rect 480574 130046 480642 130102
rect 480698 130046 480768 130102
rect 480448 129978 480768 130046
rect 480448 129922 480518 129978
rect 480574 129922 480642 129978
rect 480698 129922 480768 129978
rect 480448 129888 480768 129922
rect 496938 130350 497558 147922
rect 496938 130294 497034 130350
rect 497090 130294 497158 130350
rect 497214 130294 497282 130350
rect 497338 130294 497406 130350
rect 497462 130294 497558 130350
rect 496938 130226 497558 130294
rect 496938 130170 497034 130226
rect 497090 130170 497158 130226
rect 497214 130170 497282 130226
rect 497338 130170 497406 130226
rect 497462 130170 497558 130226
rect 496938 130102 497558 130170
rect 496938 130046 497034 130102
rect 497090 130046 497158 130102
rect 497214 130046 497282 130102
rect 497338 130046 497406 130102
rect 497462 130046 497558 130102
rect 496938 129978 497558 130046
rect 496938 129922 497034 129978
rect 497090 129922 497158 129978
rect 497214 129922 497282 129978
rect 497338 129922 497406 129978
rect 497462 129922 497558 129978
rect 473676 128458 473732 128468
rect 473676 127988 473732 128402
rect 473676 127922 473732 127932
rect 476028 127988 476084 127998
rect 476028 127918 476084 127932
rect 476028 127852 476084 127862
rect 473004 126578 473060 126588
rect 496938 125454 497558 129922
rect 500658 262350 501278 262994
rect 500658 262294 500754 262350
rect 500810 262294 500878 262350
rect 500934 262294 501002 262350
rect 501058 262294 501126 262350
rect 501182 262294 501278 262350
rect 500658 262226 501278 262294
rect 500658 262170 500754 262226
rect 500810 262170 500878 262226
rect 500934 262170 501002 262226
rect 501058 262170 501126 262226
rect 501182 262170 501278 262226
rect 500658 262102 501278 262170
rect 500658 262046 500754 262102
rect 500810 262046 500878 262102
rect 500934 262046 501002 262102
rect 501058 262046 501126 262102
rect 501182 262046 501278 262102
rect 500658 261978 501278 262046
rect 500658 261922 500754 261978
rect 500810 261922 500878 261978
rect 500934 261922 501002 261978
rect 501058 261922 501126 261978
rect 501182 261922 501278 261978
rect 500658 244350 501278 261922
rect 517692 258356 517748 273662
rect 517804 265748 517860 273812
rect 517804 265682 517860 265692
rect 519148 260372 519204 289100
rect 521052 284900 521108 284910
rect 520828 283220 520884 283230
rect 520828 278516 520884 283164
rect 520828 278450 520884 278460
rect 520940 283108 520996 283118
rect 520940 264404 520996 283052
rect 520940 264338 520996 264348
rect 521052 262388 521108 284844
rect 523292 283108 523348 293020
rect 523292 283042 523348 283052
rect 527658 292350 528278 309922
rect 527658 292294 527754 292350
rect 527810 292294 527878 292350
rect 527934 292294 528002 292350
rect 528058 292294 528126 292350
rect 528182 292294 528278 292350
rect 527658 292226 528278 292294
rect 527658 292170 527754 292226
rect 527810 292170 527878 292226
rect 527934 292170 528002 292226
rect 528058 292170 528126 292226
rect 528182 292170 528278 292226
rect 527658 292102 528278 292170
rect 527658 292046 527754 292102
rect 527810 292046 527878 292102
rect 527934 292046 528002 292102
rect 528058 292046 528126 292102
rect 528182 292046 528278 292102
rect 527658 291978 528278 292046
rect 527658 291922 527754 291978
rect 527810 291922 527878 291978
rect 527934 291922 528002 291978
rect 528058 291922 528126 291978
rect 528182 291922 528278 291978
rect 521052 262322 521108 262332
rect 527658 274350 528278 291922
rect 527658 274294 527754 274350
rect 527810 274294 527878 274350
rect 527934 274294 528002 274350
rect 528058 274294 528126 274350
rect 528182 274294 528278 274350
rect 527658 274226 528278 274294
rect 527658 274170 527754 274226
rect 527810 274170 527878 274226
rect 527934 274170 528002 274226
rect 528058 274170 528126 274226
rect 528182 274170 528278 274226
rect 527658 274102 528278 274170
rect 527658 274046 527754 274102
rect 527810 274046 527878 274102
rect 527934 274046 528002 274102
rect 528058 274046 528126 274102
rect 528182 274046 528278 274102
rect 527658 273978 528278 274046
rect 527658 273922 527754 273978
rect 527810 273922 527878 273978
rect 527934 273922 528002 273978
rect 528058 273922 528126 273978
rect 528182 273922 528278 273978
rect 519148 260306 519204 260316
rect 517692 258290 517748 258300
rect 517468 258238 517524 258248
rect 517468 258132 517524 258182
rect 517468 258066 517524 258076
rect 511168 256350 511488 256384
rect 511168 256294 511238 256350
rect 511294 256294 511362 256350
rect 511418 256294 511488 256350
rect 511168 256226 511488 256294
rect 511168 256170 511238 256226
rect 511294 256170 511362 256226
rect 511418 256170 511488 256226
rect 511168 256102 511488 256170
rect 511168 256046 511238 256102
rect 511294 256046 511362 256102
rect 511418 256046 511488 256102
rect 511168 255978 511488 256046
rect 511168 255922 511238 255978
rect 511294 255922 511362 255978
rect 511418 255922 511488 255978
rect 511168 255888 511488 255922
rect 527658 256350 528278 273922
rect 527658 256294 527754 256350
rect 527810 256294 527878 256350
rect 527934 256294 528002 256350
rect 528058 256294 528126 256350
rect 528182 256294 528278 256350
rect 527658 256226 528278 256294
rect 527658 256170 527754 256226
rect 527810 256170 527878 256226
rect 527934 256170 528002 256226
rect 528058 256170 528126 256226
rect 528182 256170 528278 256226
rect 527658 256102 528278 256170
rect 527658 256046 527754 256102
rect 527810 256046 527878 256102
rect 527934 256046 528002 256102
rect 528058 256046 528126 256102
rect 528182 256046 528278 256102
rect 527658 255978 528278 256046
rect 527658 255922 527754 255978
rect 527810 255922 527878 255978
rect 527934 255922 528002 255978
rect 528058 255922 528126 255978
rect 528182 255922 528278 255978
rect 500658 244294 500754 244350
rect 500810 244294 500878 244350
rect 500934 244294 501002 244350
rect 501058 244294 501126 244350
rect 501182 244294 501278 244350
rect 500658 244226 501278 244294
rect 500658 244170 500754 244226
rect 500810 244170 500878 244226
rect 500934 244170 501002 244226
rect 501058 244170 501126 244226
rect 501182 244170 501278 244226
rect 500658 244102 501278 244170
rect 500658 244046 500754 244102
rect 500810 244046 500878 244102
rect 500934 244046 501002 244102
rect 501058 244046 501126 244102
rect 501182 244046 501278 244102
rect 500658 243978 501278 244046
rect 500658 243922 500754 243978
rect 500810 243922 500878 243978
rect 500934 243922 501002 243978
rect 501058 243922 501126 243978
rect 501182 243922 501278 243978
rect 500658 226350 501278 243922
rect 527658 238350 528278 255922
rect 527658 238294 527754 238350
rect 527810 238294 527878 238350
rect 527934 238294 528002 238350
rect 528058 238294 528126 238350
rect 528182 238294 528278 238350
rect 527658 238226 528278 238294
rect 527658 238170 527754 238226
rect 527810 238170 527878 238226
rect 527934 238170 528002 238226
rect 528058 238170 528126 238226
rect 528182 238170 528278 238226
rect 527658 238102 528278 238170
rect 527658 238046 527754 238102
rect 527810 238046 527878 238102
rect 527934 238046 528002 238102
rect 528058 238046 528126 238102
rect 528182 238046 528278 238102
rect 527658 237978 528278 238046
rect 527658 237922 527754 237978
rect 527810 237922 527878 237978
rect 527934 237922 528002 237978
rect 528058 237922 528126 237978
rect 528182 237922 528278 237978
rect 518364 231476 518420 231486
rect 500658 226294 500754 226350
rect 500810 226294 500878 226350
rect 500934 226294 501002 226350
rect 501058 226294 501126 226350
rect 501182 226294 501278 226350
rect 500658 226226 501278 226294
rect 500658 226170 500754 226226
rect 500810 226170 500878 226226
rect 500934 226170 501002 226226
rect 501058 226170 501126 226226
rect 501182 226170 501278 226226
rect 500658 226102 501278 226170
rect 500658 226046 500754 226102
rect 500810 226046 500878 226102
rect 500934 226046 501002 226102
rect 501058 226046 501126 226102
rect 501182 226046 501278 226102
rect 500658 225978 501278 226046
rect 500658 225922 500754 225978
rect 500810 225922 500878 225978
rect 500934 225922 501002 225978
rect 501058 225922 501126 225978
rect 501182 225922 501278 225978
rect 500658 208350 501278 225922
rect 500658 208294 500754 208350
rect 500810 208294 500878 208350
rect 500934 208294 501002 208350
rect 501058 208294 501126 208350
rect 501182 208294 501278 208350
rect 500658 208226 501278 208294
rect 500658 208170 500754 208226
rect 500810 208170 500878 208226
rect 500934 208170 501002 208226
rect 501058 208170 501126 208226
rect 501182 208170 501278 208226
rect 500658 208102 501278 208170
rect 500658 208046 500754 208102
rect 500810 208046 500878 208102
rect 500934 208046 501002 208102
rect 501058 208046 501126 208102
rect 501182 208046 501278 208102
rect 500658 207978 501278 208046
rect 500658 207922 500754 207978
rect 500810 207922 500878 207978
rect 500934 207922 501002 207978
rect 501058 207922 501126 207978
rect 501182 207922 501278 207978
rect 500658 190350 501278 207922
rect 518252 226996 518308 227006
rect 511168 202350 511488 202384
rect 511168 202294 511238 202350
rect 511294 202294 511362 202350
rect 511418 202294 511488 202350
rect 511168 202226 511488 202294
rect 511168 202170 511238 202226
rect 511294 202170 511362 202226
rect 511418 202170 511488 202226
rect 511168 202102 511488 202170
rect 511168 202046 511238 202102
rect 511294 202046 511362 202102
rect 511418 202046 511488 202102
rect 511168 201978 511488 202046
rect 511168 201922 511238 201978
rect 511294 201922 511362 201978
rect 511418 201922 511488 201978
rect 511168 201888 511488 201922
rect 500658 190294 500754 190350
rect 500810 190294 500878 190350
rect 500934 190294 501002 190350
rect 501058 190294 501126 190350
rect 501182 190294 501278 190350
rect 500658 190226 501278 190294
rect 500658 190170 500754 190226
rect 500810 190170 500878 190226
rect 500934 190170 501002 190226
rect 501058 190170 501126 190226
rect 501182 190170 501278 190226
rect 500658 190102 501278 190170
rect 500658 190046 500754 190102
rect 500810 190046 500878 190102
rect 500934 190046 501002 190102
rect 501058 190046 501126 190102
rect 501182 190046 501278 190102
rect 500658 189978 501278 190046
rect 500658 189922 500754 189978
rect 500810 189922 500878 189978
rect 500934 189922 501002 189978
rect 501058 189922 501126 189978
rect 501182 189922 501278 189978
rect 500658 172350 501278 189922
rect 511168 184350 511488 184384
rect 511168 184294 511238 184350
rect 511294 184294 511362 184350
rect 511418 184294 511488 184350
rect 511168 184226 511488 184294
rect 511168 184170 511238 184226
rect 511294 184170 511362 184226
rect 511418 184170 511488 184226
rect 511168 184102 511488 184170
rect 511168 184046 511238 184102
rect 511294 184046 511362 184102
rect 511418 184046 511488 184102
rect 511168 183978 511488 184046
rect 511168 183922 511238 183978
rect 511294 183922 511362 183978
rect 511418 183922 511488 183978
rect 511168 183888 511488 183922
rect 518252 176372 518308 226940
rect 518364 191492 518420 231420
rect 519932 229796 519988 229806
rect 518364 191426 518420 191436
rect 519148 200818 519204 200828
rect 519148 189812 519204 200762
rect 519932 193284 519988 229740
rect 520156 228676 520212 228686
rect 520156 196420 520212 228620
rect 520940 224420 520996 224430
rect 520940 196532 520996 224364
rect 527658 220350 528278 237922
rect 527658 220294 527754 220350
rect 527810 220294 527878 220350
rect 527934 220294 528002 220350
rect 528058 220294 528126 220350
rect 528182 220294 528278 220350
rect 527658 220226 528278 220294
rect 527658 220170 527754 220226
rect 527810 220170 527878 220226
rect 527934 220170 528002 220226
rect 528058 220170 528126 220226
rect 528182 220170 528278 220226
rect 527658 220102 528278 220170
rect 527658 220046 527754 220102
rect 527810 220046 527878 220102
rect 527934 220046 528002 220102
rect 528058 220046 528126 220102
rect 528182 220046 528278 220102
rect 527658 219978 528278 220046
rect 527658 219922 527754 219978
rect 527810 219922 527878 219978
rect 527934 219922 528002 219978
rect 528058 219922 528126 219978
rect 528182 219922 528278 219978
rect 521164 213108 521220 213118
rect 520940 196466 520996 196476
rect 521052 211204 521108 211214
rect 520156 196354 520212 196364
rect 519932 193218 519988 193228
rect 521052 192500 521108 211148
rect 521052 192434 521108 192444
rect 519148 189746 519204 189756
rect 521164 181748 521220 213052
rect 526652 205138 526708 205148
rect 524972 203338 525028 203348
rect 524972 196532 525028 203282
rect 524972 196466 525028 196476
rect 526652 192358 526708 205082
rect 526652 192292 526708 192302
rect 527658 202350 528278 219922
rect 527658 202294 527754 202350
rect 527810 202294 527878 202350
rect 527934 202294 528002 202350
rect 528058 202294 528126 202350
rect 528182 202294 528278 202350
rect 527658 202226 528278 202294
rect 527658 202170 527754 202226
rect 527810 202170 527878 202226
rect 527934 202170 528002 202226
rect 528058 202170 528126 202226
rect 528182 202170 528278 202226
rect 527658 202102 528278 202170
rect 527658 202046 527754 202102
rect 527810 202046 527878 202102
rect 527934 202046 528002 202102
rect 528058 202046 528126 202102
rect 528182 202046 528278 202102
rect 527658 201978 528278 202046
rect 527658 201922 527754 201978
rect 527810 201922 527878 201978
rect 527934 201922 528002 201978
rect 528058 201922 528126 201978
rect 528182 201922 528278 201978
rect 521164 181682 521220 181692
rect 527658 184350 528278 201922
rect 527658 184294 527754 184350
rect 527810 184294 527878 184350
rect 527934 184294 528002 184350
rect 528058 184294 528126 184350
rect 528182 184294 528278 184350
rect 527658 184226 528278 184294
rect 527658 184170 527754 184226
rect 527810 184170 527878 184226
rect 527934 184170 528002 184226
rect 528058 184170 528126 184226
rect 528182 184170 528278 184226
rect 527658 184102 528278 184170
rect 527658 184046 527754 184102
rect 527810 184046 527878 184102
rect 527934 184046 528002 184102
rect 528058 184046 528126 184102
rect 528182 184046 528278 184102
rect 527658 183978 528278 184046
rect 527658 183922 527754 183978
rect 527810 183922 527878 183978
rect 527934 183922 528002 183978
rect 528058 183922 528126 183978
rect 528182 183922 528278 183978
rect 518252 176306 518308 176316
rect 500658 172294 500754 172350
rect 500810 172294 500878 172350
rect 500934 172294 501002 172350
rect 501058 172294 501126 172350
rect 501182 172294 501278 172350
rect 500658 172226 501278 172294
rect 500658 172170 500754 172226
rect 500810 172170 500878 172226
rect 500934 172170 501002 172226
rect 501058 172170 501126 172226
rect 501182 172170 501278 172226
rect 500658 172102 501278 172170
rect 500658 172046 500754 172102
rect 500810 172046 500878 172102
rect 500934 172046 501002 172102
rect 501058 172046 501126 172102
rect 501182 172046 501278 172102
rect 500658 171978 501278 172046
rect 500658 171922 500754 171978
rect 500810 171922 500878 171978
rect 500934 171922 501002 171978
rect 501058 171922 501126 171978
rect 501182 171922 501278 171978
rect 500658 154350 501278 171922
rect 500658 154294 500754 154350
rect 500810 154294 500878 154350
rect 500934 154294 501002 154350
rect 501058 154294 501126 154350
rect 501182 154294 501278 154350
rect 500658 154226 501278 154294
rect 500658 154170 500754 154226
rect 500810 154170 500878 154226
rect 500934 154170 501002 154226
rect 501058 154170 501126 154226
rect 501182 154170 501278 154226
rect 500658 154102 501278 154170
rect 500658 154046 500754 154102
rect 500810 154046 500878 154102
rect 500934 154046 501002 154102
rect 501058 154046 501126 154102
rect 501182 154046 501278 154102
rect 500658 153978 501278 154046
rect 500658 153922 500754 153978
rect 500810 153922 500878 153978
rect 500934 153922 501002 153978
rect 501058 153922 501126 153978
rect 501182 153922 501278 153978
rect 500658 136350 501278 153922
rect 500658 136294 500754 136350
rect 500810 136294 500878 136350
rect 500934 136294 501002 136350
rect 501058 136294 501126 136350
rect 501182 136294 501278 136350
rect 500658 136226 501278 136294
rect 500658 136170 500754 136226
rect 500810 136170 500878 136226
rect 500934 136170 501002 136226
rect 501058 136170 501126 136226
rect 501182 136170 501278 136226
rect 500658 136102 501278 136170
rect 500658 136046 500754 136102
rect 500810 136046 500878 136102
rect 500934 136046 501002 136102
rect 501058 136046 501126 136102
rect 501182 136046 501278 136102
rect 500658 135978 501278 136046
rect 500658 135922 500754 135978
rect 500810 135922 500878 135978
rect 500934 135922 501002 135978
rect 501058 135922 501126 135978
rect 501182 135922 501278 135978
rect 495808 118350 496128 118384
rect 495808 118294 495878 118350
rect 495934 118294 496002 118350
rect 496058 118294 496128 118350
rect 495808 118226 496128 118294
rect 495808 118170 495878 118226
rect 495934 118170 496002 118226
rect 496058 118170 496128 118226
rect 495808 118102 496128 118170
rect 495808 118046 495878 118102
rect 495934 118046 496002 118102
rect 496058 118046 496128 118102
rect 495808 117978 496128 118046
rect 495808 117922 495878 117978
rect 495934 117922 496002 117978
rect 496058 117922 496128 117978
rect 495808 117888 496128 117922
rect 500658 118350 501278 135922
rect 517468 173236 517524 173246
rect 511168 130350 511488 130384
rect 511168 130294 511238 130350
rect 511294 130294 511362 130350
rect 511418 130294 511488 130350
rect 511168 130226 511488 130294
rect 511168 130170 511238 130226
rect 511294 130170 511362 130226
rect 511418 130170 511488 130226
rect 511168 130102 511488 130170
rect 511168 130046 511238 130102
rect 511294 130046 511362 130102
rect 511418 130046 511488 130102
rect 511168 129978 511488 130046
rect 511168 129922 511238 129978
rect 511294 129922 511362 129978
rect 511418 129922 511488 129978
rect 511168 129888 511488 129922
rect 517468 126644 517524 173180
rect 520828 170548 520884 170558
rect 519148 167636 519204 167646
rect 517692 142548 517748 142558
rect 517468 126578 517524 126588
rect 517580 141876 517636 141886
rect 500658 118294 500754 118350
rect 500810 118294 500878 118350
rect 500934 118294 501002 118350
rect 501058 118294 501126 118350
rect 501182 118294 501278 118350
rect 500658 118226 501278 118294
rect 500658 118170 500754 118226
rect 500810 118170 500878 118226
rect 500934 118170 501002 118226
rect 501058 118170 501126 118226
rect 501182 118170 501278 118226
rect 500658 118102 501278 118170
rect 500658 118046 500754 118102
rect 500810 118046 500878 118102
rect 500934 118046 501002 118102
rect 501058 118046 501126 118102
rect 501182 118046 501278 118102
rect 500658 117978 501278 118046
rect 500658 117922 500754 117978
rect 500810 117922 500878 117978
rect 500934 117922 501002 117978
rect 501058 117922 501126 117978
rect 501182 117922 501278 117978
rect 472892 117170 472948 117180
rect 480448 112350 480768 112384
rect 480448 112294 480518 112350
rect 480574 112294 480642 112350
rect 480698 112294 480768 112350
rect 480448 112226 480768 112294
rect 480448 112170 480518 112226
rect 480574 112170 480642 112226
rect 480698 112170 480768 112226
rect 480448 112102 480768 112170
rect 480448 112046 480518 112102
rect 480574 112046 480642 112102
rect 480698 112046 480768 112102
rect 480448 111978 480768 112046
rect 480448 111922 480518 111978
rect 480574 111922 480642 111978
rect 480698 111922 480768 111978
rect 480448 111888 480768 111922
rect 496938 112350 497558 115106
rect 496938 112294 497034 112350
rect 497090 112294 497158 112350
rect 497214 112294 497282 112350
rect 497338 112294 497406 112350
rect 497462 112294 497558 112350
rect 496938 112226 497558 112294
rect 496938 112170 497034 112226
rect 497090 112170 497158 112226
rect 497214 112170 497282 112226
rect 497338 112170 497406 112226
rect 497462 112170 497558 112226
rect 496938 112102 497558 112170
rect 496938 112046 497034 112102
rect 497090 112046 497158 112102
rect 497214 112046 497282 112102
rect 497338 112046 497406 112102
rect 497462 112046 497558 112102
rect 496938 111978 497558 112046
rect 496938 111922 497034 111978
rect 497090 111922 497158 111978
rect 497214 111922 497282 111978
rect 497338 111922 497406 111978
rect 497462 111922 497558 111978
rect 469938 100294 470034 100350
rect 470090 100294 470158 100350
rect 470214 100294 470282 100350
rect 470338 100294 470406 100350
rect 470462 100294 470558 100350
rect 469938 100226 470558 100294
rect 469938 100170 470034 100226
rect 470090 100170 470158 100226
rect 470214 100170 470282 100226
rect 470338 100170 470406 100226
rect 470462 100170 470558 100226
rect 469938 100102 470558 100170
rect 469938 100046 470034 100102
rect 470090 100046 470158 100102
rect 470214 100046 470282 100102
rect 470338 100046 470406 100102
rect 470462 100046 470558 100102
rect 469938 99978 470558 100046
rect 469938 99922 470034 99978
rect 470090 99922 470158 99978
rect 470214 99922 470282 99978
rect 470338 99922 470406 99978
rect 470462 99922 470558 99978
rect 469938 82350 470558 99922
rect 496938 94350 497558 111922
rect 496938 94294 497034 94350
rect 497090 94294 497158 94350
rect 497214 94294 497282 94350
rect 497338 94294 497406 94350
rect 497462 94294 497558 94350
rect 496938 94226 497558 94294
rect 496938 94170 497034 94226
rect 497090 94170 497158 94226
rect 497214 94170 497282 94226
rect 497338 94170 497406 94226
rect 497462 94170 497558 94226
rect 496938 94102 497558 94170
rect 496938 94046 497034 94102
rect 497090 94046 497158 94102
rect 497214 94046 497282 94102
rect 497338 94046 497406 94102
rect 497462 94046 497558 94102
rect 496938 93978 497558 94046
rect 496938 93922 497034 93978
rect 497090 93922 497158 93978
rect 497214 93922 497282 93978
rect 497338 93922 497406 93978
rect 497462 93922 497558 93978
rect 469938 82294 470034 82350
rect 470090 82294 470158 82350
rect 470214 82294 470282 82350
rect 470338 82294 470406 82350
rect 470462 82294 470558 82350
rect 469938 82226 470558 82294
rect 469938 82170 470034 82226
rect 470090 82170 470158 82226
rect 470214 82170 470282 82226
rect 470338 82170 470406 82226
rect 470462 82170 470558 82226
rect 469938 82102 470558 82170
rect 469938 82046 470034 82102
rect 470090 82046 470158 82102
rect 470214 82046 470282 82102
rect 470338 82046 470406 82102
rect 470462 82046 470558 82102
rect 469938 81978 470558 82046
rect 469938 81922 470034 81978
rect 470090 81922 470158 81978
rect 470214 81922 470282 81978
rect 470338 81922 470406 81978
rect 470462 81922 470558 81978
rect 469938 64350 470558 81922
rect 469938 64294 470034 64350
rect 470090 64294 470158 64350
rect 470214 64294 470282 64350
rect 470338 64294 470406 64350
rect 470462 64294 470558 64350
rect 469938 64226 470558 64294
rect 469938 64170 470034 64226
rect 470090 64170 470158 64226
rect 470214 64170 470282 64226
rect 470338 64170 470406 64226
rect 470462 64170 470558 64226
rect 469938 64102 470558 64170
rect 469938 64046 470034 64102
rect 470090 64046 470158 64102
rect 470214 64046 470282 64102
rect 470338 64046 470406 64102
rect 470462 64046 470558 64102
rect 469938 63978 470558 64046
rect 469938 63922 470034 63978
rect 470090 63922 470158 63978
rect 470214 63922 470282 63978
rect 470338 63922 470406 63978
rect 470462 63922 470558 63978
rect 469938 46350 470558 63922
rect 469938 46294 470034 46350
rect 470090 46294 470158 46350
rect 470214 46294 470282 46350
rect 470338 46294 470406 46350
rect 470462 46294 470558 46350
rect 469938 46226 470558 46294
rect 469938 46170 470034 46226
rect 470090 46170 470158 46226
rect 470214 46170 470282 46226
rect 470338 46170 470406 46226
rect 470462 46170 470558 46226
rect 469938 46102 470558 46170
rect 469938 46046 470034 46102
rect 470090 46046 470158 46102
rect 470214 46046 470282 46102
rect 470338 46046 470406 46102
rect 470462 46046 470558 46102
rect 469938 45978 470558 46046
rect 469938 45922 470034 45978
rect 470090 45922 470158 45978
rect 470214 45922 470282 45978
rect 470338 45922 470406 45978
rect 470462 45922 470558 45978
rect 469938 28350 470558 45922
rect 472892 84868 472948 84878
rect 472892 44772 472948 84812
rect 496938 76350 497558 93922
rect 496938 76294 497034 76350
rect 497090 76294 497158 76350
rect 497214 76294 497282 76350
rect 497338 76294 497406 76350
rect 497462 76294 497558 76350
rect 496938 76226 497558 76294
rect 496938 76170 497034 76226
rect 497090 76170 497158 76226
rect 497214 76170 497282 76226
rect 497338 76170 497406 76226
rect 497462 76170 497558 76226
rect 496938 76102 497558 76170
rect 496938 76046 497034 76102
rect 497090 76046 497158 76102
rect 497214 76046 497282 76102
rect 497338 76046 497406 76102
rect 497462 76046 497558 76102
rect 496938 75978 497558 76046
rect 496938 75922 497034 75978
rect 497090 75922 497158 75978
rect 497214 75922 497282 75978
rect 497338 75922 497406 75978
rect 497462 75922 497558 75978
rect 495808 64350 496128 64384
rect 495808 64294 495878 64350
rect 495934 64294 496002 64350
rect 496058 64294 496128 64350
rect 495808 64226 496128 64294
rect 495808 64170 495878 64226
rect 495934 64170 496002 64226
rect 496058 64170 496128 64226
rect 495808 64102 496128 64170
rect 495808 64046 495878 64102
rect 495934 64046 496002 64102
rect 496058 64046 496128 64102
rect 495808 63978 496128 64046
rect 495808 63922 495878 63978
rect 495934 63922 496002 63978
rect 496058 63922 496128 63978
rect 495808 63888 496128 63922
rect 480448 58350 480768 58384
rect 480448 58294 480518 58350
rect 480574 58294 480642 58350
rect 480698 58294 480768 58350
rect 480448 58226 480768 58294
rect 480448 58170 480518 58226
rect 480574 58170 480642 58226
rect 480698 58170 480768 58226
rect 480448 58102 480768 58170
rect 480448 58046 480518 58102
rect 480574 58046 480642 58102
rect 480698 58046 480768 58102
rect 480448 57978 480768 58046
rect 480448 57922 480518 57978
rect 480574 57922 480642 57978
rect 480698 57922 480768 57978
rect 480448 57888 480768 57922
rect 496938 58350 497558 75922
rect 496938 58294 497034 58350
rect 497090 58294 497158 58350
rect 497214 58294 497282 58350
rect 497338 58294 497406 58350
rect 497462 58294 497558 58350
rect 496938 58226 497558 58294
rect 496938 58170 497034 58226
rect 497090 58170 497158 58226
rect 497214 58170 497282 58226
rect 497338 58170 497406 58226
rect 497462 58170 497558 58226
rect 496938 58102 497558 58170
rect 496938 58046 497034 58102
rect 497090 58046 497158 58102
rect 497214 58046 497282 58102
rect 497338 58046 497406 58102
rect 497462 58046 497558 58102
rect 496938 57978 497558 58046
rect 496938 57922 497034 57978
rect 497090 57922 497158 57978
rect 497214 57922 497282 57978
rect 497338 57922 497406 57978
rect 497462 57922 497558 57978
rect 473676 56278 473732 56288
rect 473676 56196 473732 56222
rect 473676 56130 473732 56140
rect 495808 46350 496128 46384
rect 495808 46294 495878 46350
rect 495934 46294 496002 46350
rect 496058 46294 496128 46350
rect 495808 46226 496128 46294
rect 495808 46170 495878 46226
rect 495934 46170 496002 46226
rect 496058 46170 496128 46226
rect 495808 46102 496128 46170
rect 495808 46046 495878 46102
rect 495934 46046 496002 46102
rect 496058 46046 496128 46102
rect 495808 45978 496128 46046
rect 495808 45922 495878 45978
rect 495934 45922 496002 45978
rect 496058 45922 496128 45978
rect 495808 45888 496128 45922
rect 472892 44706 472948 44716
rect 480448 40350 480768 40384
rect 480448 40294 480518 40350
rect 480574 40294 480642 40350
rect 480698 40294 480768 40350
rect 480448 40226 480768 40294
rect 480448 40170 480518 40226
rect 480574 40170 480642 40226
rect 480698 40170 480768 40226
rect 480448 40102 480768 40170
rect 480448 40046 480518 40102
rect 480574 40046 480642 40102
rect 480698 40046 480768 40102
rect 480448 39978 480768 40046
rect 480448 39922 480518 39978
rect 480574 39922 480642 39978
rect 480698 39922 480768 39978
rect 480448 39888 480768 39922
rect 496938 40350 497558 57922
rect 496938 40294 497034 40350
rect 497090 40294 497158 40350
rect 497214 40294 497282 40350
rect 497338 40294 497406 40350
rect 497462 40294 497558 40350
rect 496938 40226 497558 40294
rect 496938 40170 497034 40226
rect 497090 40170 497158 40226
rect 497214 40170 497282 40226
rect 497338 40170 497406 40226
rect 497462 40170 497558 40226
rect 496938 40102 497558 40170
rect 496938 40046 497034 40102
rect 497090 40046 497158 40102
rect 497214 40046 497282 40102
rect 497338 40046 497406 40102
rect 497462 40046 497558 40102
rect 496938 39978 497558 40046
rect 496938 39922 497034 39978
rect 497090 39922 497158 39978
rect 497214 39922 497282 39978
rect 497338 39922 497406 39978
rect 497462 39922 497558 39978
rect 469938 28294 470034 28350
rect 470090 28294 470158 28350
rect 470214 28294 470282 28350
rect 470338 28294 470406 28350
rect 470462 28294 470558 28350
rect 469938 28226 470558 28294
rect 469938 28170 470034 28226
rect 470090 28170 470158 28226
rect 470214 28170 470282 28226
rect 470338 28170 470406 28226
rect 470462 28170 470558 28226
rect 469938 28102 470558 28170
rect 469938 28046 470034 28102
rect 470090 28046 470158 28102
rect 470214 28046 470282 28102
rect 470338 28046 470406 28102
rect 470462 28046 470558 28102
rect 469938 27978 470558 28046
rect 469938 27922 470034 27978
rect 470090 27922 470158 27978
rect 470214 27922 470282 27978
rect 470338 27922 470406 27978
rect 470462 27922 470558 27978
rect 469938 10350 470558 27922
rect 469938 10294 470034 10350
rect 470090 10294 470158 10350
rect 470214 10294 470282 10350
rect 470338 10294 470406 10350
rect 470462 10294 470558 10350
rect 469938 10226 470558 10294
rect 469938 10170 470034 10226
rect 470090 10170 470158 10226
rect 470214 10170 470282 10226
rect 470338 10170 470406 10226
rect 470462 10170 470558 10226
rect 469938 10102 470558 10170
rect 469938 10046 470034 10102
rect 470090 10046 470158 10102
rect 470214 10046 470282 10102
rect 470338 10046 470406 10102
rect 470462 10046 470558 10102
rect 469938 9978 470558 10046
rect 469938 9922 470034 9978
rect 470090 9922 470158 9978
rect 470214 9922 470282 9978
rect 470338 9922 470406 9978
rect 470462 9922 470558 9978
rect 469938 -1120 470558 9922
rect 469938 -1176 470034 -1120
rect 470090 -1176 470158 -1120
rect 470214 -1176 470282 -1120
rect 470338 -1176 470406 -1120
rect 470462 -1176 470558 -1120
rect 469938 -1244 470558 -1176
rect 469938 -1300 470034 -1244
rect 470090 -1300 470158 -1244
rect 470214 -1300 470282 -1244
rect 470338 -1300 470406 -1244
rect 470462 -1300 470558 -1244
rect 469938 -1368 470558 -1300
rect 469938 -1424 470034 -1368
rect 470090 -1424 470158 -1368
rect 470214 -1424 470282 -1368
rect 470338 -1424 470406 -1368
rect 470462 -1424 470558 -1368
rect 469938 -1492 470558 -1424
rect 469938 -1548 470034 -1492
rect 470090 -1548 470158 -1492
rect 470214 -1548 470282 -1492
rect 470338 -1548 470406 -1492
rect 470462 -1548 470558 -1492
rect 469938 -1644 470558 -1548
rect 496938 22350 497558 39922
rect 496938 22294 497034 22350
rect 497090 22294 497158 22350
rect 497214 22294 497282 22350
rect 497338 22294 497406 22350
rect 497462 22294 497558 22350
rect 496938 22226 497558 22294
rect 496938 22170 497034 22226
rect 497090 22170 497158 22226
rect 497214 22170 497282 22226
rect 497338 22170 497406 22226
rect 497462 22170 497558 22226
rect 496938 22102 497558 22170
rect 496938 22046 497034 22102
rect 497090 22046 497158 22102
rect 497214 22046 497282 22102
rect 497338 22046 497406 22102
rect 497462 22046 497558 22102
rect 496938 21978 497558 22046
rect 496938 21922 497034 21978
rect 497090 21922 497158 21978
rect 497214 21922 497282 21978
rect 497338 21922 497406 21978
rect 497462 21922 497558 21978
rect 496938 4350 497558 21922
rect 496938 4294 497034 4350
rect 497090 4294 497158 4350
rect 497214 4294 497282 4350
rect 497338 4294 497406 4350
rect 497462 4294 497558 4350
rect 496938 4226 497558 4294
rect 496938 4170 497034 4226
rect 497090 4170 497158 4226
rect 497214 4170 497282 4226
rect 497338 4170 497406 4226
rect 497462 4170 497558 4226
rect 496938 4102 497558 4170
rect 496938 4046 497034 4102
rect 497090 4046 497158 4102
rect 497214 4046 497282 4102
rect 497338 4046 497406 4102
rect 497462 4046 497558 4102
rect 496938 3978 497558 4046
rect 496938 3922 497034 3978
rect 497090 3922 497158 3978
rect 497214 3922 497282 3978
rect 497338 3922 497406 3978
rect 497462 3922 497558 3978
rect 496938 -160 497558 3922
rect 496938 -216 497034 -160
rect 497090 -216 497158 -160
rect 497214 -216 497282 -160
rect 497338 -216 497406 -160
rect 497462 -216 497558 -160
rect 496938 -284 497558 -216
rect 496938 -340 497034 -284
rect 497090 -340 497158 -284
rect 497214 -340 497282 -284
rect 497338 -340 497406 -284
rect 497462 -340 497558 -284
rect 496938 -408 497558 -340
rect 496938 -464 497034 -408
rect 497090 -464 497158 -408
rect 497214 -464 497282 -408
rect 497338 -464 497406 -408
rect 497462 -464 497558 -408
rect 496938 -532 497558 -464
rect 496938 -588 497034 -532
rect 497090 -588 497158 -532
rect 497214 -588 497282 -532
rect 497338 -588 497406 -532
rect 497462 -588 497558 -532
rect 496938 -1644 497558 -588
rect 500658 100350 501278 117922
rect 517580 116564 517636 141820
rect 517692 119812 517748 142492
rect 517692 119746 517748 119756
rect 517580 116498 517636 116508
rect 519148 115892 519204 167580
rect 519260 144116 519316 144126
rect 519260 122612 519316 144060
rect 519372 140196 519428 140206
rect 519372 125972 519428 140140
rect 519372 125906 519428 125916
rect 519260 122546 519316 122556
rect 520828 120596 520884 170492
rect 527658 166350 528278 183922
rect 527658 166294 527754 166350
rect 527810 166294 527878 166350
rect 527934 166294 528002 166350
rect 528058 166294 528126 166350
rect 528182 166294 528278 166350
rect 527658 166226 528278 166294
rect 527658 166170 527754 166226
rect 527810 166170 527878 166226
rect 527934 166170 528002 166226
rect 528058 166170 528126 166226
rect 528182 166170 528278 166226
rect 527658 166102 528278 166170
rect 527658 166046 527754 166102
rect 527810 166046 527878 166102
rect 527934 166046 528002 166102
rect 528058 166046 528126 166102
rect 528182 166046 528278 166102
rect 527658 165978 528278 166046
rect 527658 165922 527754 165978
rect 527810 165922 527878 165978
rect 527934 165922 528002 165978
rect 528058 165922 528126 165978
rect 528182 165922 528278 165978
rect 520828 120530 520884 120540
rect 520940 160580 520996 160590
rect 520940 117236 520996 160524
rect 526652 150276 526708 150286
rect 524972 149716 525028 149726
rect 523292 149156 523348 149166
rect 521052 140420 521108 140430
rect 521052 119924 521108 140364
rect 523292 124628 523348 149100
rect 524972 125300 525028 149660
rect 524972 125234 525028 125244
rect 523292 124562 523348 124572
rect 526652 123284 526708 150220
rect 526652 123218 526708 123228
rect 527658 148350 528278 165922
rect 527658 148294 527754 148350
rect 527810 148294 527878 148350
rect 527934 148294 528002 148350
rect 528058 148294 528126 148350
rect 528182 148294 528278 148350
rect 527658 148226 528278 148294
rect 527658 148170 527754 148226
rect 527810 148170 527878 148226
rect 527934 148170 528002 148226
rect 528058 148170 528126 148226
rect 528182 148170 528278 148226
rect 527658 148102 528278 148170
rect 527658 148046 527754 148102
rect 527810 148046 527878 148102
rect 527934 148046 528002 148102
rect 528058 148046 528126 148102
rect 528182 148046 528278 148102
rect 527658 147978 528278 148046
rect 527658 147922 527754 147978
rect 527810 147922 527878 147978
rect 527934 147922 528002 147978
rect 528058 147922 528126 147978
rect 528182 147922 528278 147978
rect 527658 130350 528278 147922
rect 527658 130294 527754 130350
rect 527810 130294 527878 130350
rect 527934 130294 528002 130350
rect 528058 130294 528126 130350
rect 528182 130294 528278 130350
rect 527658 130226 528278 130294
rect 527658 130170 527754 130226
rect 527810 130170 527878 130226
rect 527934 130170 528002 130226
rect 528058 130170 528126 130226
rect 528182 130170 528278 130226
rect 527658 130102 528278 130170
rect 527658 130046 527754 130102
rect 527810 130046 527878 130102
rect 527934 130046 528002 130102
rect 528058 130046 528126 130102
rect 528182 130046 528278 130102
rect 527658 129978 528278 130046
rect 527658 129922 527754 129978
rect 527810 129922 527878 129978
rect 527934 129922 528002 129978
rect 528058 129922 528126 129978
rect 528182 129922 528278 129978
rect 521052 119858 521108 119868
rect 520940 117170 520996 117180
rect 519148 115826 519204 115836
rect 511168 112350 511488 112384
rect 511168 112294 511238 112350
rect 511294 112294 511362 112350
rect 511418 112294 511488 112350
rect 511168 112226 511488 112294
rect 511168 112170 511238 112226
rect 511294 112170 511362 112226
rect 511418 112170 511488 112226
rect 511168 112102 511488 112170
rect 511168 112046 511238 112102
rect 511294 112046 511362 112102
rect 511418 112046 511488 112102
rect 511168 111978 511488 112046
rect 511168 111922 511238 111978
rect 511294 111922 511362 111978
rect 511418 111922 511488 111978
rect 511168 111888 511488 111922
rect 527658 112350 528278 129922
rect 531378 370350 531998 387922
rect 533372 409444 533428 409454
rect 533372 379876 533428 409388
rect 535052 408100 535108 408110
rect 534268 402958 534324 402968
rect 534268 402052 534324 402902
rect 534268 401986 534324 401996
rect 533372 379810 533428 379820
rect 533484 398580 533540 398590
rect 533484 377636 533540 398524
rect 535052 385700 535108 408044
rect 557808 406350 558128 406384
rect 557808 406294 557878 406350
rect 557934 406294 558002 406350
rect 558058 406294 558128 406350
rect 557808 406226 558128 406294
rect 557808 406170 557878 406226
rect 557934 406170 558002 406226
rect 558058 406170 558128 406226
rect 557808 406102 558128 406170
rect 557808 406046 557878 406102
rect 557934 406046 558002 406102
rect 558058 406046 558128 406102
rect 557808 405978 558128 406046
rect 557808 405922 557878 405978
rect 557934 405922 558002 405978
rect 558058 405922 558128 405978
rect 557808 405888 558128 405922
rect 535612 400708 535668 400718
rect 535612 398580 535668 400652
rect 542448 400350 542768 400384
rect 542448 400294 542518 400350
rect 542574 400294 542642 400350
rect 542698 400294 542768 400350
rect 542448 400226 542768 400294
rect 542448 400170 542518 400226
rect 542574 400170 542642 400226
rect 542698 400170 542768 400226
rect 542448 400102 542768 400170
rect 542448 400046 542518 400102
rect 542574 400046 542642 400102
rect 542698 400046 542768 400102
rect 542448 399978 542768 400046
rect 542448 399922 542518 399978
rect 542574 399922 542642 399978
rect 542698 399922 542768 399978
rect 542448 399888 542768 399922
rect 558378 400350 558998 417922
rect 558378 400294 558474 400350
rect 558530 400294 558598 400350
rect 558654 400294 558722 400350
rect 558778 400294 558846 400350
rect 558902 400294 558998 400350
rect 558378 400226 558998 400294
rect 558378 400170 558474 400226
rect 558530 400170 558598 400226
rect 558654 400170 558722 400226
rect 558778 400170 558846 400226
rect 558902 400170 558998 400226
rect 558378 400102 558998 400170
rect 558378 400046 558474 400102
rect 558530 400046 558598 400102
rect 558654 400046 558722 400102
rect 558778 400046 558846 400102
rect 558902 400046 558998 400102
rect 558378 399978 558998 400046
rect 558378 399922 558474 399978
rect 558530 399922 558598 399978
rect 558654 399922 558722 399978
rect 558778 399922 558846 399978
rect 558902 399922 558998 399978
rect 535612 398514 535668 398524
rect 557808 388389 558128 388446
rect 557808 388333 557836 388389
rect 557892 388333 557940 388389
rect 557996 388333 558044 388389
rect 558100 388333 558128 388389
rect 557808 388276 558128 388333
rect 535052 385634 535108 385644
rect 533484 377570 533540 377580
rect 558378 382350 558998 399922
rect 558378 382294 558474 382350
rect 558530 382294 558598 382350
rect 558654 382294 558722 382350
rect 558778 382294 558846 382350
rect 558902 382294 558998 382350
rect 558378 382226 558998 382294
rect 558378 382170 558474 382226
rect 558530 382170 558598 382226
rect 558654 382170 558722 382226
rect 558778 382170 558846 382226
rect 558902 382170 558998 382226
rect 558378 382102 558998 382170
rect 558378 382046 558474 382102
rect 558530 382046 558598 382102
rect 558654 382046 558722 382102
rect 558778 382046 558846 382102
rect 558902 382046 558998 382102
rect 558378 381978 558998 382046
rect 558378 381922 558474 381978
rect 558530 381922 558598 381978
rect 558654 381922 558722 381978
rect 558778 381922 558846 381978
rect 558902 381922 558998 381978
rect 531378 370294 531474 370350
rect 531530 370294 531598 370350
rect 531654 370294 531722 370350
rect 531778 370294 531846 370350
rect 531902 370294 531998 370350
rect 531378 370226 531998 370294
rect 531378 370170 531474 370226
rect 531530 370170 531598 370226
rect 531654 370170 531722 370226
rect 531778 370170 531846 370226
rect 531902 370170 531998 370226
rect 531378 370102 531998 370170
rect 531378 370046 531474 370102
rect 531530 370046 531598 370102
rect 531654 370046 531722 370102
rect 531778 370046 531846 370102
rect 531902 370046 531998 370102
rect 531378 369978 531998 370046
rect 531378 369922 531474 369978
rect 531530 369922 531598 369978
rect 531654 369922 531722 369978
rect 531778 369922 531846 369978
rect 531902 369922 531998 369978
rect 531378 352350 531998 369922
rect 558378 364350 558998 381922
rect 558378 364294 558474 364350
rect 558530 364294 558598 364350
rect 558654 364294 558722 364350
rect 558778 364294 558846 364350
rect 558902 364294 558998 364350
rect 558378 364226 558998 364294
rect 558378 364170 558474 364226
rect 558530 364170 558598 364226
rect 558654 364170 558722 364226
rect 558778 364170 558846 364226
rect 558902 364170 558998 364226
rect 558378 364102 558998 364170
rect 558378 364046 558474 364102
rect 558530 364046 558598 364102
rect 558654 364046 558722 364102
rect 558778 364046 558846 364102
rect 558902 364046 558998 364102
rect 558378 363978 558998 364046
rect 558378 363922 558474 363978
rect 558530 363922 558598 363978
rect 558654 363922 558722 363978
rect 558778 363922 558846 363978
rect 558902 363922 558998 363978
rect 531378 352294 531474 352350
rect 531530 352294 531598 352350
rect 531654 352294 531722 352350
rect 531778 352294 531846 352350
rect 531902 352294 531998 352350
rect 531378 352226 531998 352294
rect 531378 352170 531474 352226
rect 531530 352170 531598 352226
rect 531654 352170 531722 352226
rect 531778 352170 531846 352226
rect 531902 352170 531998 352226
rect 531378 352102 531998 352170
rect 531378 352046 531474 352102
rect 531530 352046 531598 352102
rect 531654 352046 531722 352102
rect 531778 352046 531846 352102
rect 531902 352046 531998 352102
rect 531378 351978 531998 352046
rect 531378 351922 531474 351978
rect 531530 351922 531598 351978
rect 531654 351922 531722 351978
rect 531778 351922 531846 351978
rect 531902 351922 531998 351978
rect 531378 334350 531998 351922
rect 535164 353108 535220 353118
rect 534268 341938 534324 341948
rect 534268 341684 534324 341882
rect 534268 341618 534324 341628
rect 531378 334294 531474 334350
rect 531530 334294 531598 334350
rect 531654 334294 531722 334350
rect 531778 334294 531846 334350
rect 531902 334294 531998 334350
rect 531378 334226 531998 334294
rect 535164 334292 535220 353052
rect 557808 352350 558128 352384
rect 557808 352294 557878 352350
rect 557934 352294 558002 352350
rect 558058 352294 558128 352350
rect 557808 352226 558128 352294
rect 557808 352170 557878 352226
rect 557934 352170 558002 352226
rect 558058 352170 558128 352226
rect 557808 352102 558128 352170
rect 557808 352046 557878 352102
rect 557934 352046 558002 352102
rect 558058 352046 558128 352102
rect 557808 351978 558128 352046
rect 557808 351922 557878 351978
rect 557934 351922 558002 351978
rect 558058 351922 558128 351978
rect 557808 351888 558128 351922
rect 542448 346350 542768 346384
rect 542448 346294 542518 346350
rect 542574 346294 542642 346350
rect 542698 346294 542768 346350
rect 542448 346226 542768 346294
rect 542448 346170 542518 346226
rect 542574 346170 542642 346226
rect 542698 346170 542768 346226
rect 542448 346102 542768 346170
rect 542448 346046 542518 346102
rect 542574 346046 542642 346102
rect 542698 346046 542768 346102
rect 542448 345978 542768 346046
rect 542448 345922 542518 345978
rect 542574 345922 542642 345978
rect 542698 345922 542768 345978
rect 542448 345888 542768 345922
rect 558378 346350 558998 363922
rect 558378 346294 558474 346350
rect 558530 346294 558598 346350
rect 558654 346294 558722 346350
rect 558778 346294 558846 346350
rect 558902 346294 558998 346350
rect 558378 346226 558998 346294
rect 558378 346170 558474 346226
rect 558530 346170 558598 346226
rect 558654 346170 558722 346226
rect 558778 346170 558846 346226
rect 558902 346170 558998 346226
rect 558378 346102 558998 346170
rect 558378 346046 558474 346102
rect 558530 346046 558598 346102
rect 558654 346046 558722 346102
rect 558778 346046 558846 346102
rect 558902 346046 558998 346102
rect 558378 345978 558998 346046
rect 558378 345922 558474 345978
rect 558530 345922 558598 345978
rect 558654 345922 558722 345978
rect 558778 345922 558846 345978
rect 558902 345922 558998 345978
rect 535164 334226 535220 334236
rect 557808 334350 558128 334384
rect 557808 334294 557878 334350
rect 557934 334294 558002 334350
rect 558058 334294 558128 334350
rect 557808 334226 558128 334294
rect 531378 334170 531474 334226
rect 531530 334170 531598 334226
rect 531654 334170 531722 334226
rect 531778 334170 531846 334226
rect 531902 334170 531998 334226
rect 531378 334102 531998 334170
rect 531378 334046 531474 334102
rect 531530 334046 531598 334102
rect 531654 334046 531722 334102
rect 531778 334046 531846 334102
rect 531902 334046 531998 334102
rect 531378 333978 531998 334046
rect 531378 333922 531474 333978
rect 531530 333922 531598 333978
rect 531654 333922 531722 333978
rect 531778 333922 531846 333978
rect 531902 333922 531998 333978
rect 531378 316350 531998 333922
rect 557808 334170 557878 334226
rect 557934 334170 558002 334226
rect 558058 334170 558128 334226
rect 557808 334102 558128 334170
rect 557808 334046 557878 334102
rect 557934 334046 558002 334102
rect 558058 334046 558128 334102
rect 557808 333978 558128 334046
rect 557808 333922 557878 333978
rect 557934 333922 558002 333978
rect 558058 333922 558128 333978
rect 557808 333888 558128 333922
rect 534268 333620 534324 333630
rect 534268 330058 534324 333564
rect 534268 329992 534324 330002
rect 535052 330932 535108 330942
rect 535052 325018 535108 330876
rect 542448 328350 542768 328384
rect 542448 328294 542518 328350
rect 542574 328294 542642 328350
rect 542698 328294 542768 328350
rect 542448 328226 542768 328294
rect 542448 328170 542518 328226
rect 542574 328170 542642 328226
rect 542698 328170 542768 328226
rect 542448 328102 542768 328170
rect 542448 328046 542518 328102
rect 542574 328046 542642 328102
rect 542698 328046 542768 328102
rect 542448 327978 542768 328046
rect 542448 327922 542518 327978
rect 542574 327922 542642 327978
rect 542698 327922 542768 327978
rect 542448 327888 542768 327922
rect 558378 328350 558998 345922
rect 562098 460350 562718 477922
rect 579404 475972 579460 475982
rect 573168 472350 573488 472384
rect 573168 472294 573238 472350
rect 573294 472294 573362 472350
rect 573418 472294 573488 472350
rect 573168 472226 573488 472294
rect 573168 472170 573238 472226
rect 573294 472170 573362 472226
rect 573418 472170 573488 472226
rect 573168 472102 573488 472170
rect 573168 472046 573238 472102
rect 573294 472046 573362 472102
rect 573418 472046 573488 472102
rect 573168 471978 573488 472046
rect 573168 471922 573238 471978
rect 573294 471922 573362 471978
rect 573418 471922 573488 471978
rect 573168 471888 573488 471922
rect 579292 469924 579348 469934
rect 579292 469830 579348 469862
rect 579404 468658 579460 475916
rect 579404 468592 579460 468602
rect 579628 474628 579684 474638
rect 579628 468658 579684 474572
rect 579628 468592 579684 468602
rect 562098 460294 562194 460350
rect 562250 460294 562318 460350
rect 562374 460294 562442 460350
rect 562498 460294 562566 460350
rect 562622 460294 562718 460350
rect 562098 460226 562718 460294
rect 562098 460170 562194 460226
rect 562250 460170 562318 460226
rect 562374 460170 562442 460226
rect 562498 460170 562566 460226
rect 562622 460170 562718 460226
rect 562098 460102 562718 460170
rect 562098 460046 562194 460102
rect 562250 460046 562318 460102
rect 562374 460046 562442 460102
rect 562498 460046 562566 460102
rect 562622 460046 562718 460102
rect 562098 459978 562718 460046
rect 562098 459922 562194 459978
rect 562250 459922 562318 459978
rect 562374 459922 562442 459978
rect 562498 459922 562566 459978
rect 562622 459922 562718 459978
rect 562098 442350 562718 459922
rect 562098 442294 562194 442350
rect 562250 442294 562318 442350
rect 562374 442294 562442 442350
rect 562498 442294 562566 442350
rect 562622 442294 562718 442350
rect 562098 442226 562718 442294
rect 562098 442170 562194 442226
rect 562250 442170 562318 442226
rect 562374 442170 562442 442226
rect 562498 442170 562566 442226
rect 562622 442170 562718 442226
rect 562098 442102 562718 442170
rect 562098 442046 562194 442102
rect 562250 442046 562318 442102
rect 562374 442046 562442 442102
rect 562498 442046 562566 442102
rect 562622 442046 562718 442102
rect 562098 441978 562718 442046
rect 562098 441922 562194 441978
rect 562250 441922 562318 441978
rect 562374 441922 562442 441978
rect 562498 441922 562566 441978
rect 562622 441922 562718 441978
rect 562098 424350 562718 441922
rect 581308 441476 581364 482636
rect 583324 480676 583380 480686
rect 581308 441410 581364 441420
rect 581420 479332 581476 479342
rect 581420 439236 581476 479276
rect 582988 478660 583044 478670
rect 582988 470278 583044 478604
rect 582988 470212 583044 470222
rect 583324 446068 583380 480620
rect 583324 446002 583380 446012
rect 581420 439170 581476 439180
rect 562098 424294 562194 424350
rect 562250 424294 562318 424350
rect 562374 424294 562442 424350
rect 562498 424294 562566 424350
rect 562622 424294 562718 424350
rect 562098 424226 562718 424294
rect 562098 424170 562194 424226
rect 562250 424170 562318 424226
rect 562374 424170 562442 424226
rect 562498 424170 562566 424226
rect 562622 424170 562718 424226
rect 562098 424102 562718 424170
rect 562098 424046 562194 424102
rect 562250 424046 562318 424102
rect 562374 424046 562442 424102
rect 562498 424046 562566 424102
rect 562622 424046 562718 424102
rect 562098 423978 562718 424046
rect 562098 423922 562194 423978
rect 562250 423922 562318 423978
rect 562374 423922 562442 423978
rect 562498 423922 562566 423978
rect 562622 423922 562718 423978
rect 562098 406350 562718 423922
rect 573168 418350 573488 418384
rect 573168 418294 573238 418350
rect 573294 418294 573362 418350
rect 573418 418294 573488 418350
rect 573168 418226 573488 418294
rect 573168 418170 573238 418226
rect 573294 418170 573362 418226
rect 573418 418170 573488 418226
rect 573168 418102 573488 418170
rect 573168 418046 573238 418102
rect 573294 418046 573362 418102
rect 573418 418046 573488 418102
rect 573168 417978 573488 418046
rect 573168 417922 573238 417978
rect 573294 417922 573362 417978
rect 573418 417922 573488 417978
rect 573168 417888 573488 417922
rect 579628 411778 579684 411788
rect 579292 410788 579348 410798
rect 579292 410698 579348 410732
rect 579292 410632 579348 410642
rect 579628 410676 579684 411722
rect 579628 410610 579684 410620
rect 579292 409444 579348 409454
rect 579292 409350 579348 409382
rect 581308 407428 581364 407438
rect 579852 407098 579908 407108
rect 562098 406294 562194 406350
rect 562250 406294 562318 406350
rect 562374 406294 562442 406350
rect 562498 406294 562566 406350
rect 562622 406294 562718 406350
rect 562098 406226 562718 406294
rect 562098 406170 562194 406226
rect 562250 406170 562318 406226
rect 562374 406170 562442 406226
rect 562498 406170 562566 406226
rect 562622 406170 562718 406226
rect 562098 406102 562718 406170
rect 562098 406046 562194 406102
rect 562250 406046 562318 406102
rect 562374 406046 562442 406102
rect 562498 406046 562566 406102
rect 562622 406046 562718 406102
rect 562098 405978 562718 406046
rect 562098 405922 562194 405978
rect 562250 405922 562318 405978
rect 562374 405922 562442 405978
rect 562498 405922 562566 405978
rect 562622 405922 562718 405978
rect 562098 388350 562718 405922
rect 579628 406756 579684 406766
rect 579628 402778 579684 406700
rect 579852 406532 579908 407042
rect 579852 406466 579908 406476
rect 579740 403858 579796 403868
rect 579740 403172 579796 403802
rect 579740 403106 579796 403116
rect 579628 402722 579796 402778
rect 579628 402612 579684 402622
rect 579628 402518 579684 402542
rect 573168 400350 573488 400384
rect 573168 400294 573238 400350
rect 573294 400294 573362 400350
rect 573418 400294 573488 400350
rect 573168 400226 573488 400294
rect 573168 400170 573238 400226
rect 573294 400170 573362 400226
rect 573418 400170 573488 400226
rect 573168 400102 573488 400170
rect 573168 400046 573238 400102
rect 573294 400046 573362 400102
rect 573418 400046 573488 400102
rect 573168 399978 573488 400046
rect 573168 399922 573238 399978
rect 573294 399922 573362 399978
rect 573418 399922 573488 399978
rect 573168 399888 573488 399922
rect 579628 391078 579684 391114
rect 579628 391010 579684 391020
rect 562098 388294 562194 388350
rect 562250 388294 562318 388350
rect 562374 388294 562442 388350
rect 562498 388294 562566 388350
rect 562622 388294 562718 388350
rect 562098 388226 562718 388294
rect 562098 388170 562194 388226
rect 562250 388170 562318 388226
rect 562374 388170 562442 388226
rect 562498 388170 562566 388226
rect 562622 388170 562718 388226
rect 562098 388102 562718 388170
rect 562098 388046 562194 388102
rect 562250 388046 562318 388102
rect 562374 388046 562442 388102
rect 562498 388046 562566 388102
rect 562622 388046 562718 388102
rect 562098 387978 562718 388046
rect 562098 387922 562194 387978
rect 562250 387922 562318 387978
rect 562374 387922 562442 387978
rect 562498 387922 562566 387978
rect 562622 387922 562718 387978
rect 562098 370350 562718 387922
rect 579740 384748 579796 402722
rect 579628 384692 579796 384748
rect 579628 380996 579684 384692
rect 581308 383796 581364 407372
rect 583100 405412 583156 405422
rect 583100 387268 583156 405356
rect 583100 387202 583156 387212
rect 581308 383730 581364 383740
rect 579628 380930 579684 380940
rect 562098 370294 562194 370350
rect 562250 370294 562318 370350
rect 562374 370294 562442 370350
rect 562498 370294 562566 370350
rect 562622 370294 562718 370350
rect 562098 370226 562718 370294
rect 562098 370170 562194 370226
rect 562250 370170 562318 370226
rect 562374 370170 562442 370226
rect 562498 370170 562566 370226
rect 562622 370170 562718 370226
rect 562098 370102 562718 370170
rect 562098 370046 562194 370102
rect 562250 370046 562318 370102
rect 562374 370046 562442 370102
rect 562498 370046 562566 370102
rect 562622 370046 562718 370102
rect 562098 369978 562718 370046
rect 562098 369922 562194 369978
rect 562250 369922 562318 369978
rect 562374 369922 562442 369978
rect 562498 369922 562566 369978
rect 562622 369922 562718 369978
rect 562098 352350 562718 369922
rect 581308 356356 581364 356366
rect 580412 354116 580468 354126
rect 562098 352294 562194 352350
rect 562250 352294 562318 352350
rect 562374 352294 562442 352350
rect 562498 352294 562566 352350
rect 562622 352294 562718 352350
rect 562098 352226 562718 352294
rect 562098 352170 562194 352226
rect 562250 352170 562318 352226
rect 562374 352170 562442 352226
rect 562498 352170 562566 352226
rect 562622 352170 562718 352226
rect 562098 352102 562718 352170
rect 562098 352046 562194 352102
rect 562250 352046 562318 352102
rect 562374 352046 562442 352102
rect 562498 352046 562566 352102
rect 562622 352046 562718 352102
rect 562098 351978 562718 352046
rect 562098 351922 562194 351978
rect 562250 351922 562318 351978
rect 562374 351922 562442 351978
rect 562498 351922 562566 351978
rect 562622 351922 562718 351978
rect 562098 338830 562718 351922
rect 579628 352996 579684 353006
rect 573168 346350 573488 346384
rect 573168 346294 573238 346350
rect 573294 346294 573362 346350
rect 573418 346294 573488 346350
rect 573168 346226 573488 346294
rect 573168 346170 573238 346226
rect 573294 346170 573362 346226
rect 573418 346170 573488 346226
rect 573168 346102 573488 346170
rect 573168 346046 573238 346102
rect 573294 346046 573362 346102
rect 573418 346046 573488 346102
rect 573168 345978 573488 346046
rect 573168 345922 573238 345978
rect 573294 345922 573362 345978
rect 573418 345922 573488 345978
rect 573168 345888 573488 345922
rect 579628 333620 579684 352940
rect 580412 341796 580468 354060
rect 580412 341730 580468 341740
rect 581308 336980 581364 356300
rect 581420 355908 581476 355918
rect 581420 340340 581476 355852
rect 581420 340274 581476 340284
rect 583100 355796 583156 355806
rect 583100 337652 583156 355740
rect 583100 337586 583156 337596
rect 583212 352884 583268 352894
rect 581308 336914 581364 336924
rect 579628 333554 579684 333564
rect 582988 334964 583044 334974
rect 558378 328294 558474 328350
rect 558530 328294 558598 328350
rect 558654 328294 558722 328350
rect 558778 328294 558846 328350
rect 558902 328294 558998 328350
rect 558378 328226 558998 328294
rect 558378 328170 558474 328226
rect 558530 328170 558598 328226
rect 558654 328170 558722 328226
rect 558778 328170 558846 328226
rect 558902 328170 558998 328226
rect 558378 328102 558998 328170
rect 558378 328046 558474 328102
rect 558530 328046 558598 328102
rect 558654 328046 558722 328102
rect 558778 328046 558846 328102
rect 558902 328046 558998 328102
rect 558378 327978 558998 328046
rect 558378 327922 558474 327978
rect 558530 327922 558598 327978
rect 558654 327922 558722 327978
rect 558778 327922 558846 327978
rect 558902 327922 558998 327978
rect 535052 324952 535108 324962
rect 531378 316294 531474 316350
rect 531530 316294 531598 316350
rect 531654 316294 531722 316350
rect 531778 316294 531846 316350
rect 531902 316294 531998 316350
rect 531378 316226 531998 316294
rect 531378 316170 531474 316226
rect 531530 316170 531598 316226
rect 531654 316170 531722 316226
rect 531778 316170 531846 316226
rect 531902 316170 531998 316226
rect 531378 316102 531998 316170
rect 531378 316046 531474 316102
rect 531530 316046 531598 316102
rect 531654 316046 531722 316102
rect 531778 316046 531846 316102
rect 531902 316046 531998 316102
rect 531378 315978 531998 316046
rect 531378 315922 531474 315978
rect 531530 315922 531598 315978
rect 531654 315922 531722 315978
rect 531778 315922 531846 315978
rect 531902 315922 531998 315978
rect 531378 298350 531998 315922
rect 531378 298294 531474 298350
rect 531530 298294 531598 298350
rect 531654 298294 531722 298350
rect 531778 298294 531846 298350
rect 531902 298294 531998 298350
rect 531378 298226 531998 298294
rect 531378 298170 531474 298226
rect 531530 298170 531598 298226
rect 531654 298170 531722 298226
rect 531778 298170 531846 298226
rect 531902 298170 531998 298226
rect 531378 298102 531998 298170
rect 531378 298046 531474 298102
rect 531530 298046 531598 298102
rect 531654 298046 531722 298102
rect 531778 298046 531846 298102
rect 531902 298046 531998 298102
rect 531378 297978 531998 298046
rect 531378 297922 531474 297978
rect 531530 297922 531598 297978
rect 531654 297922 531722 297978
rect 531778 297922 531846 297978
rect 531902 297922 531998 297978
rect 531378 280350 531998 297922
rect 558378 310350 558998 327922
rect 558378 310294 558474 310350
rect 558530 310294 558598 310350
rect 558654 310294 558722 310350
rect 558778 310294 558846 310350
rect 558902 310294 558998 310350
rect 558378 310226 558998 310294
rect 558378 310170 558474 310226
rect 558530 310170 558598 310226
rect 558654 310170 558722 310226
rect 558778 310170 558846 310226
rect 558902 310170 558998 310226
rect 558378 310102 558998 310170
rect 558378 310046 558474 310102
rect 558530 310046 558598 310102
rect 558654 310046 558722 310102
rect 558778 310046 558846 310102
rect 558902 310046 558998 310102
rect 558378 309978 558998 310046
rect 558378 309922 558474 309978
rect 558530 309922 558598 309978
rect 558654 309922 558722 309978
rect 558778 309922 558846 309978
rect 558902 309922 558998 309978
rect 558378 292350 558998 309922
rect 558378 292294 558474 292350
rect 558530 292294 558598 292350
rect 558654 292294 558722 292350
rect 558778 292294 558846 292350
rect 558902 292294 558998 292350
rect 558378 292226 558998 292294
rect 558378 292170 558474 292226
rect 558530 292170 558598 292226
rect 558654 292170 558722 292226
rect 558778 292170 558846 292226
rect 558902 292170 558998 292226
rect 558378 292102 558998 292170
rect 558378 292046 558474 292102
rect 558530 292046 558598 292102
rect 558654 292046 558722 292102
rect 558778 292046 558846 292102
rect 558902 292046 558998 292102
rect 558378 291978 558998 292046
rect 558378 291922 558474 291978
rect 558530 291922 558598 291978
rect 558654 291922 558722 291978
rect 558778 291922 558846 291978
rect 558902 291922 558998 291978
rect 531378 280294 531474 280350
rect 531530 280294 531598 280350
rect 531654 280294 531722 280350
rect 531778 280294 531846 280350
rect 531902 280294 531998 280350
rect 531378 280226 531998 280294
rect 531378 280170 531474 280226
rect 531530 280170 531598 280226
rect 531654 280170 531722 280226
rect 531778 280170 531846 280226
rect 531902 280170 531998 280226
rect 531378 280102 531998 280170
rect 531378 280046 531474 280102
rect 531530 280046 531598 280102
rect 531654 280046 531722 280102
rect 531778 280046 531846 280102
rect 531902 280046 531998 280102
rect 531378 279978 531998 280046
rect 531378 279922 531474 279978
rect 531530 279922 531598 279978
rect 531654 279922 531722 279978
rect 531778 279922 531846 279978
rect 531902 279922 531998 279978
rect 531378 262350 531998 279922
rect 535164 284788 535220 284798
rect 534268 270452 534324 270462
rect 534268 269578 534324 270396
rect 534268 269512 534324 269522
rect 534268 268436 534324 268446
rect 534268 267958 534324 268380
rect 534268 267892 534324 267902
rect 531378 262294 531474 262350
rect 531530 262294 531598 262350
rect 531654 262294 531722 262350
rect 531778 262294 531846 262350
rect 531902 262294 531998 262350
rect 531378 262226 531998 262294
rect 531378 262170 531474 262226
rect 531530 262170 531598 262226
rect 531654 262170 531722 262226
rect 531778 262170 531846 262226
rect 531902 262170 531998 262226
rect 531378 262102 531998 262170
rect 531378 262046 531474 262102
rect 531530 262046 531598 262102
rect 531654 262046 531722 262102
rect 531778 262046 531846 262102
rect 531902 262046 531998 262102
rect 531378 261978 531998 262046
rect 531378 261922 531474 261978
rect 531530 261922 531598 261978
rect 531654 261922 531722 261978
rect 531778 261922 531846 261978
rect 531902 261922 531998 261978
rect 531378 244350 531998 261922
rect 534268 263060 534324 263070
rect 534268 260218 534324 263004
rect 534268 260152 534324 260162
rect 535164 258356 535220 284732
rect 557808 280350 558128 280384
rect 557808 280294 557878 280350
rect 557934 280294 558002 280350
rect 558058 280294 558128 280350
rect 557808 280226 558128 280294
rect 557808 280170 557878 280226
rect 557934 280170 558002 280226
rect 558058 280170 558128 280226
rect 557808 280102 558128 280170
rect 557808 280046 557878 280102
rect 557934 280046 558002 280102
rect 558058 280046 558128 280102
rect 557808 279978 558128 280046
rect 557808 279922 557878 279978
rect 557934 279922 558002 279978
rect 558058 279922 558128 279978
rect 557808 279888 558128 279922
rect 542448 274350 542768 274384
rect 542448 274294 542518 274350
rect 542574 274294 542642 274350
rect 542698 274294 542768 274350
rect 542448 274226 542768 274294
rect 542448 274170 542518 274226
rect 542574 274170 542642 274226
rect 542698 274170 542768 274226
rect 542448 274102 542768 274170
rect 542448 274046 542518 274102
rect 542574 274046 542642 274102
rect 542698 274046 542768 274102
rect 542448 273978 542768 274046
rect 542448 273922 542518 273978
rect 542574 273922 542642 273978
rect 542698 273922 542768 273978
rect 542448 273888 542768 273922
rect 558378 274350 558998 291922
rect 558378 274294 558474 274350
rect 558530 274294 558598 274350
rect 558654 274294 558722 274350
rect 558778 274294 558846 274350
rect 558902 274294 558998 274350
rect 558378 274226 558998 274294
rect 558378 274170 558474 274226
rect 558530 274170 558598 274226
rect 558654 274170 558722 274226
rect 558778 274170 558846 274226
rect 558902 274170 558998 274226
rect 558378 274102 558998 274170
rect 558378 274046 558474 274102
rect 558530 274046 558598 274102
rect 558654 274046 558722 274102
rect 558778 274046 558846 274102
rect 558902 274046 558998 274102
rect 558378 273978 558998 274046
rect 558378 273922 558474 273978
rect 558530 273922 558598 273978
rect 558654 273922 558722 273978
rect 558778 273922 558846 273978
rect 558902 273922 558998 273978
rect 557808 262350 558128 262384
rect 557808 262294 557878 262350
rect 557934 262294 558002 262350
rect 558058 262294 558128 262350
rect 557808 262226 558128 262294
rect 557808 262170 557878 262226
rect 557934 262170 558002 262226
rect 558058 262170 558128 262226
rect 557808 262102 558128 262170
rect 557808 262046 557878 262102
rect 557934 262046 558002 262102
rect 558058 262046 558128 262102
rect 557808 261978 558128 262046
rect 557808 261922 557878 261978
rect 557934 261922 558002 261978
rect 558058 261922 558128 261978
rect 557808 261888 558128 261922
rect 535164 258290 535220 258300
rect 542448 256350 542768 256384
rect 542448 256294 542518 256350
rect 542574 256294 542642 256350
rect 542698 256294 542768 256350
rect 542448 256226 542768 256294
rect 542448 256170 542518 256226
rect 542574 256170 542642 256226
rect 542698 256170 542768 256226
rect 542448 256102 542768 256170
rect 542448 256046 542518 256102
rect 542574 256046 542642 256102
rect 542698 256046 542768 256102
rect 542448 255978 542768 256046
rect 542448 255922 542518 255978
rect 542574 255922 542642 255978
rect 542698 255922 542768 255978
rect 542448 255888 542768 255922
rect 558378 256350 558998 273922
rect 558378 256294 558474 256350
rect 558530 256294 558598 256350
rect 558654 256294 558722 256350
rect 558778 256294 558846 256350
rect 558902 256294 558998 256350
rect 558378 256226 558998 256294
rect 558378 256170 558474 256226
rect 558530 256170 558598 256226
rect 558654 256170 558722 256226
rect 558778 256170 558846 256226
rect 558902 256170 558998 256226
rect 558378 256102 558998 256170
rect 558378 256046 558474 256102
rect 558530 256046 558598 256102
rect 558654 256046 558722 256102
rect 558778 256046 558846 256102
rect 558902 256046 558998 256102
rect 558378 255978 558998 256046
rect 558378 255922 558474 255978
rect 558530 255922 558598 255978
rect 558654 255922 558722 255978
rect 558778 255922 558846 255978
rect 558902 255922 558998 255978
rect 531378 244294 531474 244350
rect 531530 244294 531598 244350
rect 531654 244294 531722 244350
rect 531778 244294 531846 244350
rect 531902 244294 531998 244350
rect 531378 244226 531998 244294
rect 531378 244170 531474 244226
rect 531530 244170 531598 244226
rect 531654 244170 531722 244226
rect 531778 244170 531846 244226
rect 531902 244170 531998 244226
rect 531378 244102 531998 244170
rect 531378 244046 531474 244102
rect 531530 244046 531598 244102
rect 531654 244046 531722 244102
rect 531778 244046 531846 244102
rect 531902 244046 531998 244102
rect 531378 243978 531998 244046
rect 531378 243922 531474 243978
rect 531530 243922 531598 243978
rect 531654 243922 531722 243978
rect 531778 243922 531846 243978
rect 531902 243922 531998 243978
rect 531378 226350 531998 243922
rect 531378 226294 531474 226350
rect 531530 226294 531598 226350
rect 531654 226294 531722 226350
rect 531778 226294 531846 226350
rect 531902 226294 531998 226350
rect 531378 226226 531998 226294
rect 531378 226170 531474 226226
rect 531530 226170 531598 226226
rect 531654 226170 531722 226226
rect 531778 226170 531846 226226
rect 531902 226170 531998 226226
rect 531378 226102 531998 226170
rect 531378 226046 531474 226102
rect 531530 226046 531598 226102
rect 531654 226046 531722 226102
rect 531778 226046 531846 226102
rect 531902 226046 531998 226102
rect 531378 225978 531998 226046
rect 531378 225922 531474 225978
rect 531530 225922 531598 225978
rect 531654 225922 531722 225978
rect 531778 225922 531846 225978
rect 531902 225922 531998 225978
rect 531378 208350 531998 225922
rect 558378 238350 558998 255922
rect 558378 238294 558474 238350
rect 558530 238294 558598 238350
rect 558654 238294 558722 238350
rect 558778 238294 558846 238350
rect 558902 238294 558998 238350
rect 558378 238226 558998 238294
rect 558378 238170 558474 238226
rect 558530 238170 558598 238226
rect 558654 238170 558722 238226
rect 558778 238170 558846 238226
rect 558902 238170 558998 238226
rect 558378 238102 558998 238170
rect 558378 238046 558474 238102
rect 558530 238046 558598 238102
rect 558654 238046 558722 238102
rect 558778 238046 558846 238102
rect 558902 238046 558998 238102
rect 558378 237978 558998 238046
rect 558378 237922 558474 237978
rect 558530 237922 558598 237978
rect 558654 237922 558722 237978
rect 558778 237922 558846 237978
rect 558902 237922 558998 237978
rect 558378 220350 558998 237922
rect 558378 220294 558474 220350
rect 558530 220294 558598 220350
rect 558654 220294 558722 220350
rect 558778 220294 558846 220350
rect 558902 220294 558998 220350
rect 558378 220226 558998 220294
rect 558378 220170 558474 220226
rect 558530 220170 558598 220226
rect 558654 220170 558722 220226
rect 558778 220170 558846 220226
rect 558902 220170 558998 220226
rect 558378 220102 558998 220170
rect 558378 220046 558474 220102
rect 558530 220046 558598 220102
rect 558654 220046 558722 220102
rect 558778 220046 558846 220102
rect 558902 220046 558998 220102
rect 558378 219978 558998 220046
rect 558378 219922 558474 219978
rect 558530 219922 558598 219978
rect 558654 219922 558722 219978
rect 558778 219922 558846 219978
rect 558902 219922 558998 219978
rect 535276 214340 535332 214350
rect 531378 208294 531474 208350
rect 531530 208294 531598 208350
rect 531654 208294 531722 208350
rect 531778 208294 531846 208350
rect 531902 208294 531998 208350
rect 531378 208226 531998 208294
rect 531378 208170 531474 208226
rect 531530 208170 531598 208226
rect 531654 208170 531722 208226
rect 531778 208170 531846 208226
rect 531902 208170 531998 208226
rect 531378 208102 531998 208170
rect 531378 208046 531474 208102
rect 531530 208046 531598 208102
rect 531654 208046 531722 208102
rect 531778 208046 531846 208102
rect 531902 208046 531998 208102
rect 531378 207978 531998 208046
rect 531378 207922 531474 207978
rect 531530 207922 531598 207978
rect 531654 207922 531722 207978
rect 531778 207922 531846 207978
rect 531902 207922 531998 207978
rect 531378 190350 531998 207922
rect 535164 210644 535220 210654
rect 534268 199220 534324 199230
rect 534268 198298 534324 199164
rect 534268 198232 534324 198242
rect 535164 193172 535220 210588
rect 535276 195188 535332 214284
rect 535500 210532 535556 210542
rect 535500 195860 535556 210476
rect 557808 208350 558128 208384
rect 557808 208294 557878 208350
rect 557934 208294 558002 208350
rect 558058 208294 558128 208350
rect 557808 208226 558128 208294
rect 557808 208170 557878 208226
rect 557934 208170 558002 208226
rect 558058 208170 558128 208226
rect 557808 208102 558128 208170
rect 557808 208046 557878 208102
rect 557934 208046 558002 208102
rect 558058 208046 558128 208102
rect 557808 207978 558128 208046
rect 557808 207922 557878 207978
rect 557934 207922 558002 207978
rect 558058 207922 558128 207978
rect 557808 207888 558128 207922
rect 542448 202350 542768 202384
rect 542448 202294 542518 202350
rect 542574 202294 542642 202350
rect 542698 202294 542768 202350
rect 542448 202226 542768 202294
rect 542448 202170 542518 202226
rect 542574 202170 542642 202226
rect 542698 202170 542768 202226
rect 542448 202102 542768 202170
rect 542448 202046 542518 202102
rect 542574 202046 542642 202102
rect 542698 202046 542768 202102
rect 542448 201978 542768 202046
rect 542448 201922 542518 201978
rect 542574 201922 542642 201978
rect 542698 201922 542768 201978
rect 542448 201888 542768 201922
rect 558378 202350 558998 219922
rect 558378 202294 558474 202350
rect 558530 202294 558598 202350
rect 558654 202294 558722 202350
rect 558778 202294 558846 202350
rect 558902 202294 558998 202350
rect 558378 202226 558998 202294
rect 558378 202170 558474 202226
rect 558530 202170 558598 202226
rect 558654 202170 558722 202226
rect 558778 202170 558846 202226
rect 558902 202170 558998 202226
rect 558378 202102 558998 202170
rect 558378 202046 558474 202102
rect 558530 202046 558598 202102
rect 558654 202046 558722 202102
rect 558778 202046 558846 202102
rect 558902 202046 558998 202102
rect 558378 201978 558998 202046
rect 558378 201922 558474 201978
rect 558530 201922 558598 201978
rect 558654 201922 558722 201978
rect 558778 201922 558846 201978
rect 558902 201922 558998 201978
rect 535500 195794 535556 195804
rect 535276 195122 535332 195132
rect 535164 193106 535220 193116
rect 531378 190294 531474 190350
rect 531530 190294 531598 190350
rect 531654 190294 531722 190350
rect 531778 190294 531846 190350
rect 531902 190294 531998 190350
rect 531378 190226 531998 190294
rect 531378 190170 531474 190226
rect 531530 190170 531598 190226
rect 531654 190170 531722 190226
rect 531778 190170 531846 190226
rect 531902 190170 531998 190226
rect 531378 190102 531998 190170
rect 531378 190046 531474 190102
rect 531530 190046 531598 190102
rect 531654 190046 531722 190102
rect 531778 190046 531846 190102
rect 531902 190046 531998 190102
rect 531378 189978 531998 190046
rect 531378 189922 531474 189978
rect 531530 189922 531598 189978
rect 531654 189922 531722 189978
rect 531778 189922 531846 189978
rect 531902 189922 531998 189978
rect 531378 172350 531998 189922
rect 557808 190350 558128 190384
rect 557808 190294 557878 190350
rect 557934 190294 558002 190350
rect 558058 190294 558128 190350
rect 557808 190226 558128 190294
rect 557808 190170 557878 190226
rect 557934 190170 558002 190226
rect 558058 190170 558128 190226
rect 557808 190102 558128 190170
rect 557808 190046 557878 190102
rect 557934 190046 558002 190102
rect 558058 190046 558128 190102
rect 557808 189978 558128 190046
rect 557808 189922 557878 189978
rect 557934 189922 558002 189978
rect 558058 189922 558128 189978
rect 557808 189888 558128 189922
rect 542448 184350 542768 184384
rect 542448 184294 542518 184350
rect 542574 184294 542642 184350
rect 542698 184294 542768 184350
rect 542448 184226 542768 184294
rect 542448 184170 542518 184226
rect 542574 184170 542642 184226
rect 542698 184170 542768 184226
rect 542448 184102 542768 184170
rect 542448 184046 542518 184102
rect 542574 184046 542642 184102
rect 542698 184046 542768 184102
rect 542448 183978 542768 184046
rect 542448 183922 542518 183978
rect 542574 183922 542642 183978
rect 542698 183922 542768 183978
rect 542448 183888 542768 183922
rect 558378 184350 558998 201922
rect 558378 184294 558474 184350
rect 558530 184294 558598 184350
rect 558654 184294 558722 184350
rect 558778 184294 558846 184350
rect 558902 184294 558998 184350
rect 558378 184226 558998 184294
rect 558378 184170 558474 184226
rect 558530 184170 558598 184226
rect 558654 184170 558722 184226
rect 558778 184170 558846 184226
rect 558902 184170 558998 184226
rect 558378 184102 558998 184170
rect 558378 184046 558474 184102
rect 558530 184046 558598 184102
rect 558654 184046 558722 184102
rect 558778 184046 558846 184102
rect 558902 184046 558998 184102
rect 558378 183978 558998 184046
rect 558378 183922 558474 183978
rect 558530 183922 558598 183978
rect 558654 183922 558722 183978
rect 558778 183922 558846 183978
rect 558902 183922 558998 183978
rect 531378 172294 531474 172350
rect 531530 172294 531598 172350
rect 531654 172294 531722 172350
rect 531778 172294 531846 172350
rect 531902 172294 531998 172350
rect 531378 172226 531998 172294
rect 531378 172170 531474 172226
rect 531530 172170 531598 172226
rect 531654 172170 531722 172226
rect 531778 172170 531846 172226
rect 531902 172170 531998 172226
rect 531378 172102 531998 172170
rect 531378 172046 531474 172102
rect 531530 172046 531598 172102
rect 531654 172046 531722 172102
rect 531778 172046 531846 172102
rect 531902 172046 531998 172102
rect 531378 171978 531998 172046
rect 531378 171922 531474 171978
rect 531530 171922 531598 171978
rect 531654 171922 531722 171978
rect 531778 171922 531846 171978
rect 531902 171922 531998 171978
rect 531378 154350 531998 171922
rect 558378 166350 558998 183922
rect 558378 166294 558474 166350
rect 558530 166294 558598 166350
rect 558654 166294 558722 166350
rect 558778 166294 558846 166350
rect 558902 166294 558998 166350
rect 558378 166226 558998 166294
rect 558378 166170 558474 166226
rect 558530 166170 558598 166226
rect 558654 166170 558722 166226
rect 558778 166170 558846 166226
rect 558902 166170 558998 166226
rect 558378 166102 558998 166170
rect 558378 166046 558474 166102
rect 558530 166046 558598 166102
rect 558654 166046 558722 166102
rect 558778 166046 558846 166102
rect 558902 166046 558998 166102
rect 558378 165978 558998 166046
rect 558378 165922 558474 165978
rect 558530 165922 558598 165978
rect 558654 165922 558722 165978
rect 558778 165922 558846 165978
rect 558902 165922 558998 165978
rect 531378 154294 531474 154350
rect 531530 154294 531598 154350
rect 531654 154294 531722 154350
rect 531778 154294 531846 154350
rect 531902 154294 531998 154350
rect 531378 154226 531998 154294
rect 531378 154170 531474 154226
rect 531530 154170 531598 154226
rect 531654 154170 531722 154226
rect 531778 154170 531846 154226
rect 531902 154170 531998 154226
rect 531378 154102 531998 154170
rect 531378 154046 531474 154102
rect 531530 154046 531598 154102
rect 531654 154046 531722 154102
rect 531778 154046 531846 154102
rect 531902 154046 531998 154102
rect 531378 153978 531998 154046
rect 531378 153922 531474 153978
rect 531530 153922 531598 153978
rect 531654 153922 531722 153978
rect 531778 153922 531846 153978
rect 531902 153922 531998 153978
rect 531378 136350 531998 153922
rect 531378 136294 531474 136350
rect 531530 136294 531598 136350
rect 531654 136294 531722 136350
rect 531778 136294 531846 136350
rect 531902 136294 531998 136350
rect 531378 136226 531998 136294
rect 531378 136170 531474 136226
rect 531530 136170 531598 136226
rect 531654 136170 531722 136226
rect 531778 136170 531846 136226
rect 531902 136170 531998 136226
rect 531378 136102 531998 136170
rect 531378 136046 531474 136102
rect 531530 136046 531598 136102
rect 531654 136046 531722 136102
rect 531778 136046 531846 136102
rect 531902 136046 531998 136102
rect 531378 135978 531998 136046
rect 531378 135922 531474 135978
rect 531530 135922 531598 135978
rect 531654 135922 531722 135978
rect 531778 135922 531846 135978
rect 531902 135922 531998 135978
rect 530796 127738 530852 127748
rect 530796 127316 530852 127682
rect 530796 127250 530852 127260
rect 527658 112294 527754 112350
rect 527810 112294 527878 112350
rect 527934 112294 528002 112350
rect 528058 112294 528126 112350
rect 528182 112294 528278 112350
rect 527658 112226 528278 112294
rect 527658 112170 527754 112226
rect 527810 112170 527878 112226
rect 527934 112170 528002 112226
rect 528058 112170 528126 112226
rect 528182 112170 528278 112226
rect 527658 112102 528278 112170
rect 527658 112046 527754 112102
rect 527810 112046 527878 112102
rect 527934 112046 528002 112102
rect 528058 112046 528126 112102
rect 528182 112046 528278 112102
rect 527658 111978 528278 112046
rect 527658 111922 527754 111978
rect 527810 111922 527878 111978
rect 527934 111922 528002 111978
rect 528058 111922 528126 111978
rect 528182 111922 528278 111978
rect 500658 100294 500754 100350
rect 500810 100294 500878 100350
rect 500934 100294 501002 100350
rect 501058 100294 501126 100350
rect 501182 100294 501278 100350
rect 500658 100226 501278 100294
rect 500658 100170 500754 100226
rect 500810 100170 500878 100226
rect 500934 100170 501002 100226
rect 501058 100170 501126 100226
rect 501182 100170 501278 100226
rect 500658 100102 501278 100170
rect 500658 100046 500754 100102
rect 500810 100046 500878 100102
rect 500934 100046 501002 100102
rect 501058 100046 501126 100102
rect 501182 100046 501278 100102
rect 500658 99978 501278 100046
rect 500658 99922 500754 99978
rect 500810 99922 500878 99978
rect 500934 99922 501002 99978
rect 501058 99922 501126 99978
rect 501182 99922 501278 99978
rect 500658 82350 501278 99922
rect 500658 82294 500754 82350
rect 500810 82294 500878 82350
rect 500934 82294 501002 82350
rect 501058 82294 501126 82350
rect 501182 82294 501278 82350
rect 500658 82226 501278 82294
rect 500658 82170 500754 82226
rect 500810 82170 500878 82226
rect 500934 82170 501002 82226
rect 501058 82170 501126 82226
rect 501182 82170 501278 82226
rect 500658 82102 501278 82170
rect 500658 82046 500754 82102
rect 500810 82046 500878 82102
rect 500934 82046 501002 82102
rect 501058 82046 501126 82102
rect 501182 82046 501278 82102
rect 500658 81978 501278 82046
rect 500658 81922 500754 81978
rect 500810 81922 500878 81978
rect 500934 81922 501002 81978
rect 501058 81922 501126 81978
rect 501182 81922 501278 81978
rect 500658 64350 501278 81922
rect 500658 64294 500754 64350
rect 500810 64294 500878 64350
rect 500934 64294 501002 64350
rect 501058 64294 501126 64350
rect 501182 64294 501278 64350
rect 500658 64226 501278 64294
rect 500658 64170 500754 64226
rect 500810 64170 500878 64226
rect 500934 64170 501002 64226
rect 501058 64170 501126 64226
rect 501182 64170 501278 64226
rect 500658 64102 501278 64170
rect 500658 64046 500754 64102
rect 500810 64046 500878 64102
rect 500934 64046 501002 64102
rect 501058 64046 501126 64102
rect 501182 64046 501278 64102
rect 500658 63978 501278 64046
rect 500658 63922 500754 63978
rect 500810 63922 500878 63978
rect 500934 63922 501002 63978
rect 501058 63922 501126 63978
rect 501182 63922 501278 63978
rect 500658 46350 501278 63922
rect 517468 101108 517524 101118
rect 511168 58350 511488 58384
rect 511168 58294 511238 58350
rect 511294 58294 511362 58350
rect 511418 58294 511488 58350
rect 511168 58226 511488 58294
rect 511168 58170 511238 58226
rect 511294 58170 511362 58226
rect 511418 58170 511488 58226
rect 511168 58102 511488 58170
rect 511168 58046 511238 58102
rect 511294 58046 511362 58102
rect 511418 58046 511488 58102
rect 511168 57978 511488 58046
rect 511168 57922 511238 57978
rect 511294 57922 511362 57978
rect 511418 57922 511488 57978
rect 511168 57888 511488 57922
rect 500658 46294 500754 46350
rect 500810 46294 500878 46350
rect 500934 46294 501002 46350
rect 501058 46294 501126 46350
rect 501182 46294 501278 46350
rect 500658 46226 501278 46294
rect 500658 46170 500754 46226
rect 500810 46170 500878 46226
rect 500934 46170 501002 46226
rect 501058 46170 501126 46226
rect 501182 46170 501278 46226
rect 500658 46102 501278 46170
rect 500658 46046 500754 46102
rect 500810 46046 500878 46102
rect 500934 46046 501002 46102
rect 501058 46046 501126 46102
rect 501182 46046 501278 46102
rect 500658 45978 501278 46046
rect 500658 45922 500754 45978
rect 500810 45922 500878 45978
rect 500934 45922 501002 45978
rect 501058 45922 501126 45978
rect 501182 45922 501278 45978
rect 500658 28350 501278 45922
rect 517468 44772 517524 101052
rect 527658 94350 528278 111922
rect 531378 118350 531998 135922
rect 531378 118294 531474 118350
rect 531530 118294 531598 118350
rect 531654 118294 531722 118350
rect 531778 118294 531846 118350
rect 531902 118294 531998 118350
rect 531378 118226 531998 118294
rect 531378 118170 531474 118226
rect 531530 118170 531598 118226
rect 531654 118170 531722 118226
rect 531778 118170 531846 118226
rect 531902 118170 531998 118226
rect 531378 118102 531998 118170
rect 531378 118046 531474 118102
rect 531530 118046 531598 118102
rect 531654 118046 531722 118102
rect 531778 118046 531846 118102
rect 531902 118046 531998 118102
rect 531378 117978 531998 118046
rect 531378 117922 531474 117978
rect 531530 117922 531598 117978
rect 531654 117922 531722 117978
rect 531778 117922 531846 117978
rect 531902 117922 531998 117978
rect 527658 94294 527754 94350
rect 527810 94294 527878 94350
rect 527934 94294 528002 94350
rect 528058 94294 528126 94350
rect 528182 94294 528278 94350
rect 527658 94226 528278 94294
rect 527658 94170 527754 94226
rect 527810 94170 527878 94226
rect 527934 94170 528002 94226
rect 528058 94170 528126 94226
rect 528182 94170 528278 94226
rect 527658 94102 528278 94170
rect 527658 94046 527754 94102
rect 527810 94046 527878 94102
rect 527934 94046 528002 94102
rect 528058 94046 528126 94102
rect 528182 94046 528278 94102
rect 527658 93978 528278 94046
rect 527658 93922 527754 93978
rect 527810 93922 527878 93978
rect 527934 93922 528002 93978
rect 528058 93922 528126 93978
rect 528182 93922 528278 93978
rect 521276 93380 521332 93390
rect 519148 91588 519204 91598
rect 517580 82516 517636 82526
rect 517580 52164 517636 82460
rect 517580 52098 517636 52108
rect 518252 79716 518308 79726
rect 518252 47908 518308 79660
rect 519148 50820 519204 91532
rect 520940 89908 520996 89918
rect 519148 50754 519204 50764
rect 519260 83076 519316 83086
rect 519260 48132 519316 83020
rect 519372 80276 519428 80286
rect 519372 48804 519428 80220
rect 519372 48738 519428 48748
rect 519484 73332 519540 73342
rect 519260 48066 519316 48076
rect 518252 47842 518308 47852
rect 517468 44706 517524 44716
rect 519484 44100 519540 73276
rect 520940 51492 520996 89852
rect 521052 69972 521108 69982
rect 521052 52836 521108 69916
rect 521164 68068 521220 68078
rect 521164 53508 521220 68012
rect 521164 53442 521220 53452
rect 521052 52770 521108 52780
rect 520940 51426 520996 51436
rect 519484 44034 519540 44044
rect 521276 43428 521332 93324
rect 524972 92596 525028 92606
rect 523292 92036 523348 92046
rect 523292 52836 523348 91980
rect 523292 52770 523348 52780
rect 524972 50820 525028 92540
rect 524972 50754 525028 50764
rect 527658 76350 528278 93922
rect 527658 76294 527754 76350
rect 527810 76294 527878 76350
rect 527934 76294 528002 76350
rect 528058 76294 528126 76350
rect 528182 76294 528278 76350
rect 527658 76226 528278 76294
rect 527658 76170 527754 76226
rect 527810 76170 527878 76226
rect 527934 76170 528002 76226
rect 528058 76170 528126 76226
rect 528182 76170 528278 76226
rect 527658 76102 528278 76170
rect 527658 76046 527754 76102
rect 527810 76046 527878 76102
rect 527934 76046 528002 76102
rect 528058 76046 528126 76102
rect 528182 76046 528278 76102
rect 527658 75978 528278 76046
rect 527658 75922 527754 75978
rect 527810 75922 527878 75978
rect 527934 75922 528002 75978
rect 528058 75922 528126 75978
rect 528182 75922 528278 75978
rect 527658 58350 528278 75922
rect 527658 58294 527754 58350
rect 527810 58294 527878 58350
rect 527934 58294 528002 58350
rect 528058 58294 528126 58350
rect 528182 58294 528278 58350
rect 527658 58226 528278 58294
rect 527658 58170 527754 58226
rect 527810 58170 527878 58226
rect 527934 58170 528002 58226
rect 528058 58170 528126 58226
rect 528182 58170 528278 58226
rect 527658 58102 528278 58170
rect 527658 58046 527754 58102
rect 527810 58046 527878 58102
rect 527934 58046 528002 58102
rect 528058 58046 528126 58102
rect 528182 58046 528278 58102
rect 527658 57978 528278 58046
rect 527658 57922 527754 57978
rect 527810 57922 527878 57978
rect 527934 57922 528002 57978
rect 528058 57922 528126 57978
rect 528182 57922 528278 57978
rect 521276 43362 521332 43372
rect 511168 40350 511488 40384
rect 511168 40294 511238 40350
rect 511294 40294 511362 40350
rect 511418 40294 511488 40350
rect 511168 40226 511488 40294
rect 511168 40170 511238 40226
rect 511294 40170 511362 40226
rect 511418 40170 511488 40226
rect 511168 40102 511488 40170
rect 511168 40046 511238 40102
rect 511294 40046 511362 40102
rect 511418 40046 511488 40102
rect 511168 39978 511488 40046
rect 511168 39922 511238 39978
rect 511294 39922 511362 39978
rect 511418 39922 511488 39978
rect 511168 39888 511488 39922
rect 527658 40350 528278 57922
rect 530012 103348 530068 103358
rect 530012 48804 530068 103292
rect 530012 48738 530068 48748
rect 531378 100350 531998 117922
rect 535052 155540 535108 155550
rect 535052 117236 535108 155484
rect 558378 148350 558998 165922
rect 558378 148294 558474 148350
rect 558530 148294 558598 148350
rect 558654 148294 558722 148350
rect 558778 148294 558846 148350
rect 558902 148294 558998 148350
rect 558378 148226 558998 148294
rect 558378 148170 558474 148226
rect 558530 148170 558598 148226
rect 558654 148170 558722 148226
rect 558778 148170 558846 148226
rect 558902 148170 558998 148226
rect 558378 148102 558998 148170
rect 558378 148046 558474 148102
rect 558530 148046 558598 148102
rect 558654 148046 558722 148102
rect 558778 148046 558846 148102
rect 558902 148046 558998 148102
rect 558378 147978 558998 148046
rect 558378 147922 558474 147978
rect 558530 147922 558598 147978
rect 558654 147922 558722 147978
rect 558778 147922 558846 147978
rect 558902 147922 558998 147978
rect 535164 143780 535220 143790
rect 535164 119924 535220 143724
rect 557808 136350 558128 136384
rect 557808 136294 557878 136350
rect 557934 136294 558002 136350
rect 558058 136294 558128 136350
rect 557808 136226 558128 136294
rect 557808 136170 557878 136226
rect 557934 136170 558002 136226
rect 558058 136170 558128 136226
rect 557808 136102 558128 136170
rect 557808 136046 557878 136102
rect 557934 136046 558002 136102
rect 558058 136046 558128 136102
rect 557808 135978 558128 136046
rect 557808 135922 557878 135978
rect 557934 135922 558002 135978
rect 558058 135922 558128 135978
rect 557808 135888 558128 135922
rect 542448 130350 542768 130384
rect 542448 130294 542518 130350
rect 542574 130294 542642 130350
rect 542698 130294 542768 130350
rect 542448 130226 542768 130294
rect 542448 130170 542518 130226
rect 542574 130170 542642 130226
rect 542698 130170 542768 130226
rect 542448 130102 542768 130170
rect 542448 130046 542518 130102
rect 542574 130046 542642 130102
rect 542698 130046 542768 130102
rect 542448 129978 542768 130046
rect 542448 129922 542518 129978
rect 542574 129922 542642 129978
rect 542698 129922 542768 129978
rect 542448 129888 542768 129922
rect 558378 130350 558998 147922
rect 558378 130294 558474 130350
rect 558530 130294 558598 130350
rect 558654 130294 558722 130350
rect 558778 130294 558846 130350
rect 558902 130294 558998 130350
rect 558378 130226 558998 130294
rect 558378 130170 558474 130226
rect 558530 130170 558598 130226
rect 558654 130170 558722 130226
rect 558778 130170 558846 130226
rect 558902 130170 558998 130226
rect 558378 130102 558998 130170
rect 558378 130046 558474 130102
rect 558530 130046 558598 130102
rect 558654 130046 558722 130102
rect 558778 130046 558846 130102
rect 558902 130046 558998 130102
rect 558378 129978 558998 130046
rect 558378 129922 558474 129978
rect 558530 129922 558598 129978
rect 558654 129922 558722 129978
rect 558778 129922 558846 129978
rect 558902 129922 558998 129978
rect 535164 119858 535220 119868
rect 557808 118350 558128 118384
rect 557808 118294 557878 118350
rect 557934 118294 558002 118350
rect 558058 118294 558128 118350
rect 557808 118226 558128 118294
rect 557808 118170 557878 118226
rect 557934 118170 558002 118226
rect 558058 118170 558128 118226
rect 557808 118102 558128 118170
rect 557808 118046 557878 118102
rect 557934 118046 558002 118102
rect 558058 118046 558128 118102
rect 557808 117978 558128 118046
rect 557808 117922 557878 117978
rect 557934 117922 558002 117978
rect 558058 117922 558128 117978
rect 557808 117888 558128 117922
rect 535052 117170 535108 117180
rect 542448 112350 542768 112384
rect 542448 112294 542518 112350
rect 542574 112294 542642 112350
rect 542698 112294 542768 112350
rect 542448 112226 542768 112294
rect 542448 112170 542518 112226
rect 542574 112170 542642 112226
rect 542698 112170 542768 112226
rect 542448 112102 542768 112170
rect 542448 112046 542518 112102
rect 542574 112046 542642 112102
rect 542698 112046 542768 112102
rect 542448 111978 542768 112046
rect 542448 111922 542518 111978
rect 542574 111922 542642 111978
rect 542698 111922 542768 111978
rect 542448 111888 542768 111922
rect 558378 112350 558998 129922
rect 558378 112294 558474 112350
rect 558530 112294 558598 112350
rect 558654 112294 558722 112350
rect 558778 112294 558846 112350
rect 558902 112294 558998 112350
rect 558378 112226 558998 112294
rect 558378 112170 558474 112226
rect 558530 112170 558598 112226
rect 558654 112170 558722 112226
rect 558778 112170 558846 112226
rect 558902 112170 558998 112226
rect 558378 112102 558998 112170
rect 558378 112046 558474 112102
rect 558530 112046 558598 112102
rect 558654 112046 558722 112102
rect 558778 112046 558846 112102
rect 558902 112046 558998 112102
rect 558378 111978 558998 112046
rect 558378 111922 558474 111978
rect 558530 111922 558598 111978
rect 558654 111922 558722 111978
rect 558778 111922 558846 111978
rect 558902 111922 558998 111978
rect 531378 100294 531474 100350
rect 531530 100294 531598 100350
rect 531654 100294 531722 100350
rect 531778 100294 531846 100350
rect 531902 100294 531998 100350
rect 531378 100226 531998 100294
rect 531378 100170 531474 100226
rect 531530 100170 531598 100226
rect 531654 100170 531722 100226
rect 531778 100170 531846 100226
rect 531902 100170 531998 100226
rect 531378 100102 531998 100170
rect 531378 100046 531474 100102
rect 531530 100046 531598 100102
rect 531654 100046 531722 100102
rect 531778 100046 531846 100102
rect 531902 100046 531998 100102
rect 531378 99978 531998 100046
rect 531378 99922 531474 99978
rect 531530 99922 531598 99978
rect 531654 99922 531722 99978
rect 531778 99922 531846 99978
rect 531902 99922 531998 99978
rect 531378 82350 531998 99922
rect 531378 82294 531474 82350
rect 531530 82294 531598 82350
rect 531654 82294 531722 82350
rect 531778 82294 531846 82350
rect 531902 82294 531998 82350
rect 531378 82226 531998 82294
rect 531378 82170 531474 82226
rect 531530 82170 531598 82226
rect 531654 82170 531722 82226
rect 531778 82170 531846 82226
rect 531902 82170 531998 82226
rect 531378 82102 531998 82170
rect 531378 82046 531474 82102
rect 531530 82046 531598 82102
rect 531654 82046 531722 82102
rect 531778 82046 531846 82102
rect 531902 82046 531998 82102
rect 531378 81978 531998 82046
rect 531378 81922 531474 81978
rect 531530 81922 531598 81978
rect 531654 81922 531722 81978
rect 531778 81922 531846 81978
rect 531902 81922 531998 81978
rect 531378 64350 531998 81922
rect 531378 64294 531474 64350
rect 531530 64294 531598 64350
rect 531654 64294 531722 64350
rect 531778 64294 531846 64350
rect 531902 64294 531998 64350
rect 531378 64226 531998 64294
rect 531378 64170 531474 64226
rect 531530 64170 531598 64226
rect 531654 64170 531722 64226
rect 531778 64170 531846 64226
rect 531902 64170 531998 64226
rect 531378 64102 531998 64170
rect 531378 64046 531474 64102
rect 531530 64046 531598 64102
rect 531654 64046 531722 64102
rect 531778 64046 531846 64102
rect 531902 64046 531998 64102
rect 531378 63978 531998 64046
rect 531378 63922 531474 63978
rect 531530 63922 531598 63978
rect 531654 63922 531722 63978
rect 531778 63922 531846 63978
rect 531902 63922 531998 63978
rect 527658 40294 527754 40350
rect 527810 40294 527878 40350
rect 527934 40294 528002 40350
rect 528058 40294 528126 40350
rect 528182 40294 528278 40350
rect 527658 40226 528278 40294
rect 527658 40170 527754 40226
rect 527810 40170 527878 40226
rect 527934 40170 528002 40226
rect 528058 40170 528126 40226
rect 528182 40170 528278 40226
rect 527658 40102 528278 40170
rect 527658 40046 527754 40102
rect 527810 40046 527878 40102
rect 527934 40046 528002 40102
rect 528058 40046 528126 40102
rect 528182 40046 528278 40102
rect 527658 39978 528278 40046
rect 527658 39922 527754 39978
rect 527810 39922 527878 39978
rect 527934 39922 528002 39978
rect 528058 39922 528126 39978
rect 528182 39922 528278 39978
rect 500658 28294 500754 28350
rect 500810 28294 500878 28350
rect 500934 28294 501002 28350
rect 501058 28294 501126 28350
rect 501182 28294 501278 28350
rect 500658 28226 501278 28294
rect 500658 28170 500754 28226
rect 500810 28170 500878 28226
rect 500934 28170 501002 28226
rect 501058 28170 501126 28226
rect 501182 28170 501278 28226
rect 500658 28102 501278 28170
rect 500658 28046 500754 28102
rect 500810 28046 500878 28102
rect 500934 28046 501002 28102
rect 501058 28046 501126 28102
rect 501182 28046 501278 28102
rect 500658 27978 501278 28046
rect 500658 27922 500754 27978
rect 500810 27922 500878 27978
rect 500934 27922 501002 27978
rect 501058 27922 501126 27978
rect 501182 27922 501278 27978
rect 500658 10350 501278 27922
rect 500658 10294 500754 10350
rect 500810 10294 500878 10350
rect 500934 10294 501002 10350
rect 501058 10294 501126 10350
rect 501182 10294 501278 10350
rect 500658 10226 501278 10294
rect 500658 10170 500754 10226
rect 500810 10170 500878 10226
rect 500934 10170 501002 10226
rect 501058 10170 501126 10226
rect 501182 10170 501278 10226
rect 500658 10102 501278 10170
rect 500658 10046 500754 10102
rect 500810 10046 500878 10102
rect 500934 10046 501002 10102
rect 501058 10046 501126 10102
rect 501182 10046 501278 10102
rect 500658 9978 501278 10046
rect 500658 9922 500754 9978
rect 500810 9922 500878 9978
rect 500934 9922 501002 9978
rect 501058 9922 501126 9978
rect 501182 9922 501278 9978
rect 500658 -1120 501278 9922
rect 500658 -1176 500754 -1120
rect 500810 -1176 500878 -1120
rect 500934 -1176 501002 -1120
rect 501058 -1176 501126 -1120
rect 501182 -1176 501278 -1120
rect 500658 -1244 501278 -1176
rect 500658 -1300 500754 -1244
rect 500810 -1300 500878 -1244
rect 500934 -1300 501002 -1244
rect 501058 -1300 501126 -1244
rect 501182 -1300 501278 -1244
rect 500658 -1368 501278 -1300
rect 500658 -1424 500754 -1368
rect 500810 -1424 500878 -1368
rect 500934 -1424 501002 -1368
rect 501058 -1424 501126 -1368
rect 501182 -1424 501278 -1368
rect 500658 -1492 501278 -1424
rect 500658 -1548 500754 -1492
rect 500810 -1548 500878 -1492
rect 500934 -1548 501002 -1492
rect 501058 -1548 501126 -1492
rect 501182 -1548 501278 -1492
rect 500658 -1644 501278 -1548
rect 527658 22350 528278 39922
rect 527658 22294 527754 22350
rect 527810 22294 527878 22350
rect 527934 22294 528002 22350
rect 528058 22294 528126 22350
rect 528182 22294 528278 22350
rect 527658 22226 528278 22294
rect 527658 22170 527754 22226
rect 527810 22170 527878 22226
rect 527934 22170 528002 22226
rect 528058 22170 528126 22226
rect 528182 22170 528278 22226
rect 527658 22102 528278 22170
rect 527658 22046 527754 22102
rect 527810 22046 527878 22102
rect 527934 22046 528002 22102
rect 528058 22046 528126 22102
rect 528182 22046 528278 22102
rect 527658 21978 528278 22046
rect 527658 21922 527754 21978
rect 527810 21922 527878 21978
rect 527934 21922 528002 21978
rect 528058 21922 528126 21978
rect 528182 21922 528278 21978
rect 527658 4350 528278 21922
rect 527658 4294 527754 4350
rect 527810 4294 527878 4350
rect 527934 4294 528002 4350
rect 528058 4294 528126 4350
rect 528182 4294 528278 4350
rect 527658 4226 528278 4294
rect 527658 4170 527754 4226
rect 527810 4170 527878 4226
rect 527934 4170 528002 4226
rect 528058 4170 528126 4226
rect 528182 4170 528278 4226
rect 527658 4102 528278 4170
rect 527658 4046 527754 4102
rect 527810 4046 527878 4102
rect 527934 4046 528002 4102
rect 528058 4046 528126 4102
rect 528182 4046 528278 4102
rect 527658 3978 528278 4046
rect 527658 3922 527754 3978
rect 527810 3922 527878 3978
rect 527934 3922 528002 3978
rect 528058 3922 528126 3978
rect 528182 3922 528278 3978
rect 527658 -160 528278 3922
rect 527658 -216 527754 -160
rect 527810 -216 527878 -160
rect 527934 -216 528002 -160
rect 528058 -216 528126 -160
rect 528182 -216 528278 -160
rect 527658 -284 528278 -216
rect 527658 -340 527754 -284
rect 527810 -340 527878 -284
rect 527934 -340 528002 -284
rect 528058 -340 528126 -284
rect 528182 -340 528278 -284
rect 527658 -408 528278 -340
rect 527658 -464 527754 -408
rect 527810 -464 527878 -408
rect 527934 -464 528002 -408
rect 528058 -464 528126 -408
rect 528182 -464 528278 -408
rect 527658 -532 528278 -464
rect 527658 -588 527754 -532
rect 527810 -588 527878 -532
rect 527934 -588 528002 -532
rect 528058 -588 528126 -532
rect 528182 -588 528278 -532
rect 527658 -1644 528278 -588
rect 531378 46350 531998 63922
rect 535164 96852 535220 96862
rect 534268 56278 534324 56288
rect 534268 56196 534324 56222
rect 534268 56130 534324 56140
rect 535164 48132 535220 96796
rect 558378 94350 558998 111922
rect 558378 94294 558474 94350
rect 558530 94294 558598 94350
rect 558654 94294 558722 94350
rect 558778 94294 558846 94350
rect 558902 94294 558998 94350
rect 558378 94226 558998 94294
rect 558378 94170 558474 94226
rect 558530 94170 558598 94226
rect 558654 94170 558722 94226
rect 558778 94170 558846 94226
rect 558902 94170 558998 94226
rect 558378 94102 558998 94170
rect 558378 94046 558474 94102
rect 558530 94046 558598 94102
rect 558654 94046 558722 94102
rect 558778 94046 558846 94102
rect 558902 94046 558998 94102
rect 558378 93978 558998 94046
rect 558378 93922 558474 93978
rect 558530 93922 558598 93978
rect 558654 93922 558722 93978
rect 558778 93922 558846 93978
rect 558902 93922 558998 93978
rect 535388 78260 535444 78270
rect 535164 48066 535220 48076
rect 535276 73108 535332 73118
rect 531378 46294 531474 46350
rect 531530 46294 531598 46350
rect 531654 46294 531722 46350
rect 531778 46294 531846 46350
rect 531902 46294 531998 46350
rect 531378 46226 531998 46294
rect 531378 46170 531474 46226
rect 531530 46170 531598 46226
rect 531654 46170 531722 46226
rect 531778 46170 531846 46226
rect 531902 46170 531998 46226
rect 531378 46102 531998 46170
rect 531378 46046 531474 46102
rect 531530 46046 531598 46102
rect 531654 46046 531722 46102
rect 531778 46046 531846 46102
rect 531902 46046 531998 46102
rect 535276 46116 535332 73052
rect 535388 52164 535444 78204
rect 558378 76350 558998 93922
rect 558378 76294 558474 76350
rect 558530 76294 558598 76350
rect 558654 76294 558722 76350
rect 558778 76294 558846 76350
rect 558902 76294 558998 76350
rect 558378 76226 558998 76294
rect 558378 76170 558474 76226
rect 558530 76170 558598 76226
rect 558654 76170 558722 76226
rect 558778 76170 558846 76226
rect 558902 76170 558998 76226
rect 558378 76102 558998 76170
rect 558378 76046 558474 76102
rect 558530 76046 558598 76102
rect 558654 76046 558722 76102
rect 558778 76046 558846 76102
rect 558902 76046 558998 76102
rect 558378 75978 558998 76046
rect 558378 75922 558474 75978
rect 558530 75922 558598 75978
rect 558654 75922 558722 75978
rect 558778 75922 558846 75978
rect 558902 75922 558998 75978
rect 535388 52098 535444 52108
rect 535500 71540 535556 71550
rect 535276 46050 535332 46060
rect 531378 45978 531998 46046
rect 531378 45922 531474 45978
rect 531530 45922 531598 45978
rect 531654 45922 531722 45978
rect 531778 45922 531846 45978
rect 531902 45922 531998 45978
rect 531378 28350 531998 45922
rect 535500 45444 535556 71484
rect 535612 69860 535668 69870
rect 535612 49476 535668 69804
rect 535836 69748 535892 69758
rect 535836 54852 535892 69692
rect 557808 64350 558128 64384
rect 557808 64294 557878 64350
rect 557934 64294 558002 64350
rect 558058 64294 558128 64350
rect 557808 64226 558128 64294
rect 557808 64170 557878 64226
rect 557934 64170 558002 64226
rect 558058 64170 558128 64226
rect 557808 64102 558128 64170
rect 557808 64046 557878 64102
rect 557934 64046 558002 64102
rect 558058 64046 558128 64102
rect 557808 63978 558128 64046
rect 557808 63922 557878 63978
rect 557934 63922 558002 63978
rect 558058 63922 558128 63978
rect 557808 63888 558128 63922
rect 542448 58350 542768 58384
rect 542448 58294 542518 58350
rect 542574 58294 542642 58350
rect 542698 58294 542768 58350
rect 542448 58226 542768 58294
rect 542448 58170 542518 58226
rect 542574 58170 542642 58226
rect 542698 58170 542768 58226
rect 542448 58102 542768 58170
rect 542448 58046 542518 58102
rect 542574 58046 542642 58102
rect 542698 58046 542768 58102
rect 542448 57978 542768 58046
rect 542448 57922 542518 57978
rect 542574 57922 542642 57978
rect 542698 57922 542768 57978
rect 542448 57888 542768 57922
rect 558378 58350 558998 75922
rect 558378 58294 558474 58350
rect 558530 58294 558598 58350
rect 558654 58294 558722 58350
rect 558778 58294 558846 58350
rect 558902 58294 558998 58350
rect 558378 58226 558998 58294
rect 558378 58170 558474 58226
rect 558530 58170 558598 58226
rect 558654 58170 558722 58226
rect 558778 58170 558846 58226
rect 558902 58170 558998 58226
rect 558378 58102 558998 58170
rect 558378 58046 558474 58102
rect 558530 58046 558598 58102
rect 558654 58046 558722 58102
rect 558778 58046 558846 58102
rect 558902 58046 558998 58102
rect 558378 57978 558998 58046
rect 558378 57922 558474 57978
rect 558530 57922 558598 57978
rect 558654 57922 558722 57978
rect 558778 57922 558846 57978
rect 558902 57922 558998 57978
rect 535836 54786 535892 54796
rect 558378 52910 558998 57922
rect 562098 316350 562718 332178
rect 579628 331716 579684 331726
rect 579628 331612 579684 331622
rect 573168 328350 573488 328384
rect 573168 328294 573238 328350
rect 573294 328294 573362 328350
rect 573418 328294 573488 328350
rect 573168 328226 573488 328294
rect 573168 328170 573238 328226
rect 573294 328170 573362 328226
rect 573418 328170 573488 328226
rect 573168 328102 573488 328170
rect 573168 328046 573238 328102
rect 573294 328046 573362 328102
rect 573418 328046 573488 328102
rect 573168 327978 573488 328046
rect 573168 327922 573238 327978
rect 573294 327922 573362 327978
rect 573418 327922 573488 327978
rect 573168 327888 573488 327922
rect 582988 326818 583044 334908
rect 582988 326752 583044 326762
rect 583212 325556 583268 352828
rect 583212 325490 583268 325500
rect 562098 316294 562194 316350
rect 562250 316294 562318 316350
rect 562374 316294 562442 316350
rect 562498 316294 562566 316350
rect 562622 316294 562718 316350
rect 562098 316226 562718 316294
rect 562098 316170 562194 316226
rect 562250 316170 562318 316226
rect 562374 316170 562442 316226
rect 562498 316170 562566 316226
rect 562622 316170 562718 316226
rect 562098 316102 562718 316170
rect 562098 316046 562194 316102
rect 562250 316046 562318 316102
rect 562374 316046 562442 316102
rect 562498 316046 562566 316102
rect 562622 316046 562718 316102
rect 562098 315978 562718 316046
rect 562098 315922 562194 315978
rect 562250 315922 562318 315978
rect 562374 315922 562442 315978
rect 562498 315922 562566 315978
rect 562622 315922 562718 315978
rect 562098 298350 562718 315922
rect 562940 314132 562996 314142
rect 562940 314038 562996 314076
rect 562940 313972 562996 313982
rect 562098 298294 562194 298350
rect 562250 298294 562318 298350
rect 562374 298294 562442 298350
rect 562498 298294 562566 298350
rect 562622 298294 562718 298350
rect 562098 298226 562718 298294
rect 562098 298170 562194 298226
rect 562250 298170 562318 298226
rect 562374 298170 562442 298226
rect 562498 298170 562566 298226
rect 562622 298170 562718 298226
rect 562098 298102 562718 298170
rect 562098 298046 562194 298102
rect 562250 298046 562318 298102
rect 562374 298046 562442 298102
rect 562498 298046 562566 298102
rect 562622 298046 562718 298102
rect 562098 297978 562718 298046
rect 562098 297922 562194 297978
rect 562250 297922 562318 297978
rect 562374 297922 562442 297978
rect 562498 297922 562566 297978
rect 562622 297922 562718 297978
rect 562098 280350 562718 297922
rect 583548 295316 583604 295326
rect 582092 294756 582148 294766
rect 562098 280294 562194 280350
rect 562250 280294 562318 280350
rect 562374 280294 562442 280350
rect 562498 280294 562566 280350
rect 562622 280294 562718 280350
rect 562098 280226 562718 280294
rect 562098 280170 562194 280226
rect 562250 280170 562318 280226
rect 562374 280170 562442 280226
rect 562498 280170 562566 280226
rect 562622 280170 562718 280226
rect 562098 280102 562718 280170
rect 562098 280046 562194 280102
rect 562250 280046 562318 280102
rect 562374 280046 562442 280102
rect 562498 280046 562566 280102
rect 562622 280046 562718 280102
rect 562098 279978 562718 280046
rect 562098 279922 562194 279978
rect 562250 279922 562318 279978
rect 562374 279922 562442 279978
rect 562498 279922 562566 279978
rect 562622 279922 562718 279978
rect 562098 262350 562718 279922
rect 580412 294196 580468 294206
rect 573168 274350 573488 274384
rect 573168 274294 573238 274350
rect 573294 274294 573362 274350
rect 573418 274294 573488 274350
rect 573168 274226 573488 274294
rect 573168 274170 573238 274226
rect 573294 274170 573362 274226
rect 573418 274170 573488 274226
rect 573168 274102 573488 274170
rect 573168 274046 573238 274102
rect 573294 274046 573362 274102
rect 573418 274046 573488 274102
rect 573168 273978 573488 274046
rect 573168 273922 573238 273978
rect 573294 273922 573362 273978
rect 573418 273922 573488 273978
rect 573168 273888 573488 273922
rect 579292 267092 579348 267102
rect 579292 266992 579348 267002
rect 579068 266698 579124 266708
rect 579124 266642 579348 266698
rect 579068 266632 579124 266642
rect 579292 264404 579348 266642
rect 579292 264338 579348 264348
rect 580412 263844 580468 294140
rect 581308 293636 581364 293646
rect 580412 263778 580468 263788
rect 580524 292516 580580 292526
rect 562098 262294 562194 262350
rect 562250 262294 562318 262350
rect 562374 262294 562442 262350
rect 562498 262294 562566 262350
rect 562622 262294 562718 262350
rect 562098 262226 562718 262294
rect 562098 262170 562194 262226
rect 562250 262170 562318 262226
rect 562374 262170 562442 262226
rect 562498 262170 562566 262226
rect 562622 262170 562718 262226
rect 562098 262102 562718 262170
rect 562098 262046 562194 262102
rect 562250 262046 562318 262102
rect 562374 262046 562442 262102
rect 562498 262046 562566 262102
rect 562622 262046 562718 262102
rect 562098 261978 562718 262046
rect 562098 261922 562194 261978
rect 562250 261922 562318 261978
rect 562374 261922 562442 261978
rect 562498 261922 562566 261978
rect 562622 261922 562718 261978
rect 562098 244350 562718 261922
rect 579628 263284 579684 263294
rect 579292 261044 579348 261054
rect 579292 260938 579348 260988
rect 579292 260872 579348 260882
rect 579628 260398 579684 263228
rect 580524 262052 580580 292460
rect 580524 261986 580580 261996
rect 579628 260332 579684 260342
rect 581308 259700 581364 293580
rect 582092 266196 582148 294700
rect 583100 286468 583156 286478
rect 582092 266130 582148 266140
rect 582988 268858 583044 268868
rect 582988 262388 583044 268802
rect 583100 267764 583156 286412
rect 583212 283108 583268 283118
rect 583212 269108 583268 283052
rect 583212 269042 583268 269052
rect 583100 267698 583156 267708
rect 583548 266420 583604 295260
rect 583548 266354 583604 266364
rect 582988 262322 583044 262332
rect 581308 259634 581364 259644
rect 573168 256350 573488 256384
rect 573168 256294 573238 256350
rect 573294 256294 573362 256350
rect 573418 256294 573488 256350
rect 573168 256226 573488 256294
rect 573168 256170 573238 256226
rect 573294 256170 573362 256226
rect 573418 256170 573488 256226
rect 573168 256102 573488 256170
rect 573168 256046 573238 256102
rect 573294 256046 573362 256102
rect 573418 256046 573488 256102
rect 573168 255978 573488 256046
rect 573168 255922 573238 255978
rect 573294 255922 573362 255978
rect 573418 255922 573488 255978
rect 573168 255888 573488 255922
rect 562098 244294 562194 244350
rect 562250 244294 562318 244350
rect 562374 244294 562442 244350
rect 562498 244294 562566 244350
rect 562622 244294 562718 244350
rect 562098 244226 562718 244294
rect 562098 244170 562194 244226
rect 562250 244170 562318 244226
rect 562374 244170 562442 244226
rect 562498 244170 562566 244226
rect 562622 244170 562718 244226
rect 562098 244102 562718 244170
rect 562098 244046 562194 244102
rect 562250 244046 562318 244102
rect 562374 244046 562442 244102
rect 562498 244046 562566 244102
rect 562622 244046 562718 244102
rect 562098 243978 562718 244046
rect 562098 243922 562194 243978
rect 562250 243922 562318 243978
rect 562374 243922 562442 243978
rect 562498 243922 562566 243978
rect 562622 243922 562718 243978
rect 562098 226350 562718 243922
rect 562098 226294 562194 226350
rect 562250 226294 562318 226350
rect 562374 226294 562442 226350
rect 562498 226294 562566 226350
rect 562622 226294 562718 226350
rect 562098 226226 562718 226294
rect 562098 226170 562194 226226
rect 562250 226170 562318 226226
rect 562374 226170 562442 226226
rect 562498 226170 562566 226226
rect 562622 226170 562718 226226
rect 562098 226102 562718 226170
rect 562098 226046 562194 226102
rect 562250 226046 562318 226102
rect 562374 226046 562442 226102
rect 562498 226046 562566 226102
rect 562622 226046 562718 226102
rect 562098 225978 562718 226046
rect 562098 225922 562194 225978
rect 562250 225922 562318 225978
rect 562374 225922 562442 225978
rect 562498 225922 562566 225978
rect 562622 225922 562718 225978
rect 562098 208350 562718 225922
rect 581308 235396 581364 235406
rect 562098 208294 562194 208350
rect 562250 208294 562318 208350
rect 562374 208294 562442 208350
rect 562498 208294 562566 208350
rect 562622 208294 562718 208350
rect 562098 208226 562718 208294
rect 562098 208170 562194 208226
rect 562250 208170 562318 208226
rect 562374 208170 562442 208226
rect 562498 208170 562566 208226
rect 562622 208170 562718 208226
rect 562098 208102 562718 208170
rect 562098 208046 562194 208102
rect 562250 208046 562318 208102
rect 562374 208046 562442 208102
rect 562498 208046 562566 208102
rect 562622 208046 562718 208102
rect 562098 207978 562718 208046
rect 562098 207922 562194 207978
rect 562250 207922 562318 207978
rect 562374 207922 562442 207978
rect 562498 207922 562566 207978
rect 562622 207922 562718 207978
rect 562098 190350 562718 207922
rect 579628 219268 579684 219278
rect 573168 202350 573488 202384
rect 573168 202294 573238 202350
rect 573294 202294 573362 202350
rect 573418 202294 573488 202350
rect 573168 202226 573488 202294
rect 573168 202170 573238 202226
rect 573294 202170 573362 202226
rect 573418 202170 573488 202226
rect 573168 202102 573488 202170
rect 573168 202046 573238 202102
rect 573294 202046 573362 202102
rect 573418 202046 573488 202102
rect 573168 201978 573488 202046
rect 573168 201922 573238 201978
rect 573294 201922 573362 201978
rect 573418 201922 573488 201978
rect 573168 201888 573488 201922
rect 579628 197204 579684 219212
rect 579628 197138 579684 197148
rect 579740 192178 579796 192188
rect 579740 191044 579796 192122
rect 579740 190978 579796 190988
rect 562098 190294 562194 190350
rect 562250 190294 562318 190350
rect 562374 190294 562442 190350
rect 562498 190294 562566 190350
rect 562622 190294 562718 190350
rect 562098 190226 562718 190294
rect 562098 190170 562194 190226
rect 562250 190170 562318 190226
rect 562374 190170 562442 190226
rect 562498 190170 562566 190226
rect 562622 190170 562718 190226
rect 562098 190102 562718 190170
rect 562098 190046 562194 190102
rect 562250 190046 562318 190102
rect 562374 190046 562442 190102
rect 562498 190046 562566 190102
rect 562622 190046 562718 190102
rect 562098 189978 562718 190046
rect 562098 189922 562194 189978
rect 562250 189922 562318 189978
rect 562374 189922 562442 189978
rect 562498 189922 562566 189978
rect 562622 189922 562718 189978
rect 562098 172350 562718 189922
rect 581308 189140 581364 235340
rect 583436 233716 583492 233726
rect 583100 231028 583156 231038
rect 581420 224308 581476 224318
rect 581420 195860 581476 224252
rect 581420 195794 581476 195804
rect 583100 193172 583156 230972
rect 583324 210980 583380 210990
rect 583100 193106 583156 193116
rect 583212 210420 583268 210430
rect 581308 189074 581364 189084
rect 583212 187124 583268 210364
rect 583324 196532 583380 210924
rect 583324 196466 583380 196476
rect 583436 189812 583492 233660
rect 583436 189746 583492 189756
rect 583212 187058 583268 187068
rect 573168 184350 573488 184384
rect 573168 184294 573238 184350
rect 573294 184294 573362 184350
rect 573418 184294 573488 184350
rect 573168 184226 573488 184294
rect 573168 184170 573238 184226
rect 573294 184170 573362 184226
rect 573418 184170 573488 184226
rect 573168 184102 573488 184170
rect 573168 184046 573238 184102
rect 573294 184046 573362 184102
rect 573418 184046 573488 184102
rect 573168 183978 573488 184046
rect 573168 183922 573238 183978
rect 573294 183922 573362 183978
rect 573418 183922 573488 183978
rect 573168 183888 573488 183922
rect 562098 172294 562194 172350
rect 562250 172294 562318 172350
rect 562374 172294 562442 172350
rect 562498 172294 562566 172350
rect 562622 172294 562718 172350
rect 562098 172226 562718 172294
rect 562098 172170 562194 172226
rect 562250 172170 562318 172226
rect 562374 172170 562442 172226
rect 562498 172170 562566 172226
rect 562622 172170 562718 172226
rect 562098 172102 562718 172170
rect 562098 172046 562194 172102
rect 562250 172046 562318 172102
rect 562374 172046 562442 172102
rect 562498 172046 562566 172102
rect 562622 172046 562718 172102
rect 562098 171978 562718 172046
rect 562098 171922 562194 171978
rect 562250 171922 562318 171978
rect 562374 171922 562442 171978
rect 562498 171922 562566 171978
rect 562622 171922 562718 171978
rect 562098 154350 562718 171922
rect 562098 154294 562194 154350
rect 562250 154294 562318 154350
rect 562374 154294 562442 154350
rect 562498 154294 562566 154350
rect 562622 154294 562718 154350
rect 562098 154226 562718 154294
rect 562098 154170 562194 154226
rect 562250 154170 562318 154226
rect 562374 154170 562442 154226
rect 562498 154170 562566 154226
rect 562622 154170 562718 154226
rect 562098 154102 562718 154170
rect 562098 154046 562194 154102
rect 562250 154046 562318 154102
rect 562374 154046 562442 154102
rect 562498 154046 562566 154102
rect 562622 154046 562718 154102
rect 562098 153978 562718 154046
rect 562098 153922 562194 153978
rect 562250 153922 562318 153978
rect 562374 153922 562442 153978
rect 562498 153922 562566 153978
rect 562622 153922 562718 153978
rect 562098 136350 562718 153922
rect 562098 136294 562194 136350
rect 562250 136294 562318 136350
rect 562374 136294 562442 136350
rect 562498 136294 562566 136350
rect 562622 136294 562718 136350
rect 562098 136226 562718 136294
rect 562098 136170 562194 136226
rect 562250 136170 562318 136226
rect 562374 136170 562442 136226
rect 562498 136170 562566 136226
rect 562622 136170 562718 136226
rect 562098 136102 562718 136170
rect 562098 136046 562194 136102
rect 562250 136046 562318 136102
rect 562374 136046 562442 136102
rect 562498 136046 562566 136102
rect 562622 136046 562718 136102
rect 562098 135978 562718 136046
rect 562098 135922 562194 135978
rect 562250 135922 562318 135978
rect 562374 135922 562442 135978
rect 562498 135922 562566 135978
rect 562622 135922 562718 135978
rect 562098 118350 562718 135922
rect 579628 173908 579684 173918
rect 573168 130350 573488 130384
rect 573168 130294 573238 130350
rect 573294 130294 573362 130350
rect 573418 130294 573488 130350
rect 573168 130226 573488 130294
rect 573168 130170 573238 130226
rect 573294 130170 573362 130226
rect 573418 130170 573488 130226
rect 573168 130102 573488 130170
rect 573168 130046 573238 130102
rect 573294 130046 573362 130102
rect 573418 130046 573488 130102
rect 573168 129978 573488 130046
rect 573168 129922 573238 129978
rect 573294 129922 573362 129978
rect 573418 129922 573488 129978
rect 573168 129888 573488 129922
rect 579628 123284 579684 173852
rect 582988 163828 583044 163838
rect 581308 158788 581364 158798
rect 579628 123218 579684 123228
rect 579740 146916 579796 146926
rect 579740 119812 579796 146860
rect 579740 119746 579796 119756
rect 580412 144676 580468 144686
rect 580412 118916 580468 144620
rect 581308 123956 581364 158732
rect 581532 147476 581588 147486
rect 581308 123890 581364 123900
rect 581420 146356 581476 146366
rect 581420 121940 581476 146300
rect 581532 125300 581588 147420
rect 581644 145236 581700 145246
rect 581644 126644 581700 145180
rect 582988 127316 583044 163772
rect 583212 157108 583268 157118
rect 582988 127250 583044 127260
rect 583100 155428 583156 155438
rect 581644 126578 581700 126588
rect 581532 125234 581588 125244
rect 581420 121874 581476 121884
rect 583100 121268 583156 155372
rect 583212 124628 583268 157052
rect 583436 141988 583492 141998
rect 583212 124562 583268 124572
rect 583324 140308 583380 140318
rect 583324 122612 583380 140252
rect 583436 125972 583492 141932
rect 583436 125906 583492 125916
rect 583324 122546 583380 122556
rect 583100 121202 583156 121212
rect 580412 118850 580468 118860
rect 562098 118294 562194 118350
rect 562250 118294 562318 118350
rect 562374 118294 562442 118350
rect 562498 118294 562566 118350
rect 562622 118294 562718 118350
rect 562098 118226 562718 118294
rect 562098 118170 562194 118226
rect 562250 118170 562318 118226
rect 562374 118170 562442 118226
rect 562498 118170 562566 118226
rect 562622 118170 562718 118226
rect 562098 118102 562718 118170
rect 562098 118046 562194 118102
rect 562250 118046 562318 118102
rect 562374 118046 562442 118102
rect 562498 118046 562566 118102
rect 562622 118046 562718 118102
rect 562098 117978 562718 118046
rect 562098 117922 562194 117978
rect 562250 117922 562318 117978
rect 562374 117922 562442 117978
rect 562498 117922 562566 117978
rect 562622 117922 562718 117978
rect 562098 100350 562718 117922
rect 573168 112350 573488 112384
rect 573168 112294 573238 112350
rect 573294 112294 573362 112350
rect 573418 112294 573488 112350
rect 573168 112226 573488 112294
rect 573168 112170 573238 112226
rect 573294 112170 573362 112226
rect 573418 112170 573488 112226
rect 573168 112102 573488 112170
rect 573168 112046 573238 112102
rect 573294 112046 573362 112102
rect 573418 112046 573488 112102
rect 573168 111978 573488 112046
rect 573168 111922 573238 111978
rect 573294 111922 573362 111978
rect 573418 111922 573488 111978
rect 573168 111888 573488 111922
rect 562098 100294 562194 100350
rect 562250 100294 562318 100350
rect 562374 100294 562442 100350
rect 562498 100294 562566 100350
rect 562622 100294 562718 100350
rect 562098 100226 562718 100294
rect 562098 100170 562194 100226
rect 562250 100170 562318 100226
rect 562374 100170 562442 100226
rect 562498 100170 562566 100226
rect 562622 100170 562718 100226
rect 562098 100102 562718 100170
rect 562098 100046 562194 100102
rect 562250 100046 562318 100102
rect 562374 100046 562442 100102
rect 562498 100046 562566 100102
rect 562622 100046 562718 100102
rect 562098 99978 562718 100046
rect 562098 99922 562194 99978
rect 562250 99922 562318 99978
rect 562374 99922 562442 99978
rect 562498 99922 562566 99978
rect 562622 99922 562718 99978
rect 562098 82350 562718 99922
rect 583436 96628 583492 96638
rect 562098 82294 562194 82350
rect 562250 82294 562318 82350
rect 562374 82294 562442 82350
rect 562498 82294 562566 82350
rect 562622 82294 562718 82350
rect 562098 82226 562718 82294
rect 562098 82170 562194 82226
rect 562250 82170 562318 82226
rect 562374 82170 562442 82226
rect 562498 82170 562566 82226
rect 562622 82170 562718 82226
rect 562098 82102 562718 82170
rect 562098 82046 562194 82102
rect 562250 82046 562318 82102
rect 562374 82046 562442 82102
rect 562498 82046 562566 82102
rect 562622 82046 562718 82102
rect 562098 81978 562718 82046
rect 562098 81922 562194 81978
rect 562250 81922 562318 81978
rect 562374 81922 562442 81978
rect 562498 81922 562566 81978
rect 562622 81922 562718 81978
rect 562098 64350 562718 81922
rect 562098 64294 562194 64350
rect 562250 64294 562318 64350
rect 562374 64294 562442 64350
rect 562498 64294 562566 64350
rect 562622 64294 562718 64350
rect 562098 64226 562718 64294
rect 562098 64170 562194 64226
rect 562250 64170 562318 64226
rect 562374 64170 562442 64226
rect 562498 64170 562566 64226
rect 562622 64170 562718 64226
rect 562098 64102 562718 64170
rect 562098 64046 562194 64102
rect 562250 64046 562318 64102
rect 562374 64046 562442 64102
rect 562498 64046 562566 64102
rect 562622 64046 562718 64102
rect 562098 63978 562718 64046
rect 562098 63922 562194 63978
rect 562250 63922 562318 63978
rect 562374 63922 562442 63978
rect 562498 63922 562566 63978
rect 562622 63922 562718 63978
rect 535612 49410 535668 49420
rect 557808 46350 558128 46384
rect 557808 46294 557878 46350
rect 557934 46294 558002 46350
rect 558058 46294 558128 46350
rect 557808 46226 558128 46294
rect 557808 46170 557878 46226
rect 557934 46170 558002 46226
rect 558058 46170 558128 46226
rect 557808 46102 558128 46170
rect 557808 46046 557878 46102
rect 557934 46046 558002 46102
rect 558058 46046 558128 46102
rect 557808 45978 558128 46046
rect 557808 45922 557878 45978
rect 557934 45922 558002 45978
rect 558058 45922 558128 45978
rect 557808 45888 558128 45922
rect 562098 46350 562718 63922
rect 579628 90916 579684 90926
rect 573168 58350 573488 58384
rect 573168 58294 573238 58350
rect 573294 58294 573362 58350
rect 573418 58294 573488 58350
rect 573168 58226 573488 58294
rect 573168 58170 573238 58226
rect 573294 58170 573362 58226
rect 573418 58170 573488 58226
rect 573168 58102 573488 58170
rect 573168 58046 573238 58102
rect 573294 58046 573362 58102
rect 573418 58046 573488 58102
rect 573168 57978 573488 58046
rect 573168 57922 573238 57978
rect 573294 57922 573362 57978
rect 573418 57922 573488 57978
rect 573168 57888 573488 57922
rect 579628 52836 579684 90860
rect 581308 89796 581364 89806
rect 580412 88116 580468 88126
rect 579628 52770 579684 52780
rect 579740 86436 579796 86446
rect 579740 50820 579796 86380
rect 579740 50754 579796 50764
rect 580412 47124 580468 88060
rect 581308 47460 581364 89740
rect 581420 88676 581476 88686
rect 581420 55524 581476 88620
rect 581420 55458 581476 55468
rect 581532 86996 581588 87006
rect 581532 54852 581588 86940
rect 581532 54786 581588 54796
rect 583100 79828 583156 79838
rect 581308 47394 581364 47404
rect 580412 47058 580468 47068
rect 562098 46294 562194 46350
rect 562250 46294 562318 46350
rect 562374 46294 562442 46350
rect 562498 46294 562566 46350
rect 562622 46294 562718 46350
rect 562098 46226 562718 46294
rect 562098 46170 562194 46226
rect 562250 46170 562318 46226
rect 562374 46170 562442 46226
rect 562498 46170 562566 46226
rect 562622 46170 562718 46226
rect 562098 46102 562718 46170
rect 562098 46046 562194 46102
rect 562250 46046 562318 46102
rect 562374 46046 562442 46102
rect 562498 46046 562566 46102
rect 562622 46046 562718 46102
rect 562098 45978 562718 46046
rect 562098 45922 562194 45978
rect 562250 45922 562318 45978
rect 562374 45922 562442 45978
rect 562498 45922 562566 45978
rect 562622 45922 562718 45978
rect 535500 45378 535556 45388
rect 542448 40350 542768 40384
rect 542448 40294 542518 40350
rect 542574 40294 542642 40350
rect 542698 40294 542768 40350
rect 542448 40226 542768 40294
rect 542448 40170 542518 40226
rect 542574 40170 542642 40226
rect 542698 40170 542768 40226
rect 542448 40102 542768 40170
rect 542448 40046 542518 40102
rect 542574 40046 542642 40102
rect 542698 40046 542768 40102
rect 542448 39978 542768 40046
rect 542448 39922 542518 39978
rect 542574 39922 542642 39978
rect 542698 39922 542768 39978
rect 542448 39888 542768 39922
rect 558378 40350 558998 42338
rect 558378 40294 558474 40350
rect 558530 40294 558598 40350
rect 558654 40294 558722 40350
rect 558778 40294 558846 40350
rect 558902 40294 558998 40350
rect 558378 40226 558998 40294
rect 558378 40170 558474 40226
rect 558530 40170 558598 40226
rect 558654 40170 558722 40226
rect 558778 40170 558846 40226
rect 558902 40170 558998 40226
rect 558378 40102 558998 40170
rect 558378 40046 558474 40102
rect 558530 40046 558598 40102
rect 558654 40046 558722 40102
rect 558778 40046 558846 40102
rect 558902 40046 558998 40102
rect 558378 39978 558998 40046
rect 558378 39922 558474 39978
rect 558530 39922 558598 39978
rect 558654 39922 558722 39978
rect 558778 39922 558846 39978
rect 558902 39922 558998 39978
rect 531378 28294 531474 28350
rect 531530 28294 531598 28350
rect 531654 28294 531722 28350
rect 531778 28294 531846 28350
rect 531902 28294 531998 28350
rect 531378 28226 531998 28294
rect 531378 28170 531474 28226
rect 531530 28170 531598 28226
rect 531654 28170 531722 28226
rect 531778 28170 531846 28226
rect 531902 28170 531998 28226
rect 531378 28102 531998 28170
rect 531378 28046 531474 28102
rect 531530 28046 531598 28102
rect 531654 28046 531722 28102
rect 531778 28046 531846 28102
rect 531902 28046 531998 28102
rect 531378 27978 531998 28046
rect 531378 27922 531474 27978
rect 531530 27922 531598 27978
rect 531654 27922 531722 27978
rect 531778 27922 531846 27978
rect 531902 27922 531998 27978
rect 531378 10350 531998 27922
rect 531378 10294 531474 10350
rect 531530 10294 531598 10350
rect 531654 10294 531722 10350
rect 531778 10294 531846 10350
rect 531902 10294 531998 10350
rect 531378 10226 531998 10294
rect 531378 10170 531474 10226
rect 531530 10170 531598 10226
rect 531654 10170 531722 10226
rect 531778 10170 531846 10226
rect 531902 10170 531998 10226
rect 531378 10102 531998 10170
rect 531378 10046 531474 10102
rect 531530 10046 531598 10102
rect 531654 10046 531722 10102
rect 531778 10046 531846 10102
rect 531902 10046 531998 10102
rect 531378 9978 531998 10046
rect 531378 9922 531474 9978
rect 531530 9922 531598 9978
rect 531654 9922 531722 9978
rect 531778 9922 531846 9978
rect 531902 9922 531998 9978
rect 531378 -1120 531998 9922
rect 531378 -1176 531474 -1120
rect 531530 -1176 531598 -1120
rect 531654 -1176 531722 -1120
rect 531778 -1176 531846 -1120
rect 531902 -1176 531998 -1120
rect 531378 -1244 531998 -1176
rect 531378 -1300 531474 -1244
rect 531530 -1300 531598 -1244
rect 531654 -1300 531722 -1244
rect 531778 -1300 531846 -1244
rect 531902 -1300 531998 -1244
rect 531378 -1368 531998 -1300
rect 531378 -1424 531474 -1368
rect 531530 -1424 531598 -1368
rect 531654 -1424 531722 -1368
rect 531778 -1424 531846 -1368
rect 531902 -1424 531998 -1368
rect 531378 -1492 531998 -1424
rect 531378 -1548 531474 -1492
rect 531530 -1548 531598 -1492
rect 531654 -1548 531722 -1492
rect 531778 -1548 531846 -1492
rect 531902 -1548 531998 -1492
rect 531378 -1644 531998 -1548
rect 558378 22350 558998 39922
rect 558378 22294 558474 22350
rect 558530 22294 558598 22350
rect 558654 22294 558722 22350
rect 558778 22294 558846 22350
rect 558902 22294 558998 22350
rect 558378 22226 558998 22294
rect 558378 22170 558474 22226
rect 558530 22170 558598 22226
rect 558654 22170 558722 22226
rect 558778 22170 558846 22226
rect 558902 22170 558998 22226
rect 558378 22102 558998 22170
rect 558378 22046 558474 22102
rect 558530 22046 558598 22102
rect 558654 22046 558722 22102
rect 558778 22046 558846 22102
rect 558902 22046 558998 22102
rect 558378 21978 558998 22046
rect 558378 21922 558474 21978
rect 558530 21922 558598 21978
rect 558654 21922 558722 21978
rect 558778 21922 558846 21978
rect 558902 21922 558998 21978
rect 558378 4350 558998 21922
rect 558378 4294 558474 4350
rect 558530 4294 558598 4350
rect 558654 4294 558722 4350
rect 558778 4294 558846 4350
rect 558902 4294 558998 4350
rect 558378 4226 558998 4294
rect 558378 4170 558474 4226
rect 558530 4170 558598 4226
rect 558654 4170 558722 4226
rect 558778 4170 558846 4226
rect 558902 4170 558998 4226
rect 558378 4102 558998 4170
rect 558378 4046 558474 4102
rect 558530 4046 558598 4102
rect 558654 4046 558722 4102
rect 558778 4046 558846 4102
rect 558902 4046 558998 4102
rect 558378 3978 558998 4046
rect 558378 3922 558474 3978
rect 558530 3922 558598 3978
rect 558654 3922 558722 3978
rect 558778 3922 558846 3978
rect 558902 3922 558998 3978
rect 558378 -160 558998 3922
rect 558378 -216 558474 -160
rect 558530 -216 558598 -160
rect 558654 -216 558722 -160
rect 558778 -216 558846 -160
rect 558902 -216 558998 -160
rect 558378 -284 558998 -216
rect 558378 -340 558474 -284
rect 558530 -340 558598 -284
rect 558654 -340 558722 -284
rect 558778 -340 558846 -284
rect 558902 -340 558998 -284
rect 558378 -408 558998 -340
rect 558378 -464 558474 -408
rect 558530 -464 558598 -408
rect 558654 -464 558722 -408
rect 558778 -464 558846 -408
rect 558902 -464 558998 -408
rect 558378 -532 558998 -464
rect 558378 -588 558474 -532
rect 558530 -588 558598 -532
rect 558654 -588 558722 -532
rect 558778 -588 558846 -532
rect 558902 -588 558998 -532
rect 558378 -1644 558998 -588
rect 562098 28350 562718 45922
rect 583100 44772 583156 79772
rect 583212 71428 583268 71438
rect 583212 49476 583268 71372
rect 583324 70532 583380 70542
rect 583324 52164 583380 70476
rect 583324 52098 583380 52108
rect 583212 49410 583268 49420
rect 583436 45444 583492 96572
rect 583436 45378 583492 45388
rect 583100 44706 583156 44716
rect 573168 40350 573488 40384
rect 573168 40294 573238 40350
rect 573294 40294 573362 40350
rect 573418 40294 573488 40350
rect 573168 40226 573488 40294
rect 573168 40170 573238 40226
rect 573294 40170 573362 40226
rect 573418 40170 573488 40226
rect 573168 40102 573488 40170
rect 573168 40046 573238 40102
rect 573294 40046 573362 40102
rect 573418 40046 573488 40102
rect 573168 39978 573488 40046
rect 573168 39922 573238 39978
rect 573294 39922 573362 39978
rect 573418 39922 573488 39978
rect 573168 39888 573488 39922
rect 585452 33796 585508 566882
rect 585452 33730 585508 33740
rect 589098 562350 589718 579922
rect 589098 562294 589194 562350
rect 589250 562294 589318 562350
rect 589374 562294 589442 562350
rect 589498 562294 589566 562350
rect 589622 562294 589718 562350
rect 589098 562226 589718 562294
rect 589098 562170 589194 562226
rect 589250 562170 589318 562226
rect 589374 562170 589442 562226
rect 589498 562170 589566 562226
rect 589622 562170 589718 562226
rect 589098 562102 589718 562170
rect 589098 562046 589194 562102
rect 589250 562046 589318 562102
rect 589374 562046 589442 562102
rect 589498 562046 589566 562102
rect 589622 562046 589718 562102
rect 589098 561978 589718 562046
rect 589098 561922 589194 561978
rect 589250 561922 589318 561978
rect 589374 561922 589442 561978
rect 589498 561922 589566 561978
rect 589622 561922 589718 561978
rect 589098 544350 589718 561922
rect 589098 544294 589194 544350
rect 589250 544294 589318 544350
rect 589374 544294 589442 544350
rect 589498 544294 589566 544350
rect 589622 544294 589718 544350
rect 589098 544226 589718 544294
rect 589098 544170 589194 544226
rect 589250 544170 589318 544226
rect 589374 544170 589442 544226
rect 589498 544170 589566 544226
rect 589622 544170 589718 544226
rect 589098 544102 589718 544170
rect 589098 544046 589194 544102
rect 589250 544046 589318 544102
rect 589374 544046 589442 544102
rect 589498 544046 589566 544102
rect 589622 544046 589718 544102
rect 589098 543978 589718 544046
rect 589098 543922 589194 543978
rect 589250 543922 589318 543978
rect 589374 543922 589442 543978
rect 589498 543922 589566 543978
rect 589622 543922 589718 543978
rect 589098 526350 589718 543922
rect 589098 526294 589194 526350
rect 589250 526294 589318 526350
rect 589374 526294 589442 526350
rect 589498 526294 589566 526350
rect 589622 526294 589718 526350
rect 589098 526226 589718 526294
rect 589098 526170 589194 526226
rect 589250 526170 589318 526226
rect 589374 526170 589442 526226
rect 589498 526170 589566 526226
rect 589622 526170 589718 526226
rect 589098 526102 589718 526170
rect 589098 526046 589194 526102
rect 589250 526046 589318 526102
rect 589374 526046 589442 526102
rect 589498 526046 589566 526102
rect 589622 526046 589718 526102
rect 589098 525978 589718 526046
rect 589098 525922 589194 525978
rect 589250 525922 589318 525978
rect 589374 525922 589442 525978
rect 589498 525922 589566 525978
rect 589622 525922 589718 525978
rect 589098 508350 589718 525922
rect 589098 508294 589194 508350
rect 589250 508294 589318 508350
rect 589374 508294 589442 508350
rect 589498 508294 589566 508350
rect 589622 508294 589718 508350
rect 589098 508226 589718 508294
rect 589098 508170 589194 508226
rect 589250 508170 589318 508226
rect 589374 508170 589442 508226
rect 589498 508170 589566 508226
rect 589622 508170 589718 508226
rect 589098 508102 589718 508170
rect 589098 508046 589194 508102
rect 589250 508046 589318 508102
rect 589374 508046 589442 508102
rect 589498 508046 589566 508102
rect 589622 508046 589718 508102
rect 589098 507978 589718 508046
rect 589098 507922 589194 507978
rect 589250 507922 589318 507978
rect 589374 507922 589442 507978
rect 589498 507922 589566 507978
rect 589622 507922 589718 507978
rect 589098 490350 589718 507922
rect 589098 490294 589194 490350
rect 589250 490294 589318 490350
rect 589374 490294 589442 490350
rect 589498 490294 589566 490350
rect 589622 490294 589718 490350
rect 589098 490226 589718 490294
rect 589098 490170 589194 490226
rect 589250 490170 589318 490226
rect 589374 490170 589442 490226
rect 589498 490170 589566 490226
rect 589622 490170 589718 490226
rect 589098 490102 589718 490170
rect 589098 490046 589194 490102
rect 589250 490046 589318 490102
rect 589374 490046 589442 490102
rect 589498 490046 589566 490102
rect 589622 490046 589718 490102
rect 589098 489978 589718 490046
rect 589098 489922 589194 489978
rect 589250 489922 589318 489978
rect 589374 489922 589442 489978
rect 589498 489922 589566 489978
rect 589622 489922 589718 489978
rect 589098 472350 589718 489922
rect 589098 472294 589194 472350
rect 589250 472294 589318 472350
rect 589374 472294 589442 472350
rect 589498 472294 589566 472350
rect 589622 472294 589718 472350
rect 589098 472226 589718 472294
rect 589098 472170 589194 472226
rect 589250 472170 589318 472226
rect 589374 472170 589442 472226
rect 589498 472170 589566 472226
rect 589622 472170 589718 472226
rect 589098 472102 589718 472170
rect 589098 472046 589194 472102
rect 589250 472046 589318 472102
rect 589374 472046 589442 472102
rect 589498 472046 589566 472102
rect 589622 472046 589718 472102
rect 589098 471978 589718 472046
rect 589098 471922 589194 471978
rect 589250 471922 589318 471978
rect 589374 471922 589442 471978
rect 589498 471922 589566 471978
rect 589622 471922 589718 471978
rect 589098 454350 589718 471922
rect 589098 454294 589194 454350
rect 589250 454294 589318 454350
rect 589374 454294 589442 454350
rect 589498 454294 589566 454350
rect 589622 454294 589718 454350
rect 589098 454226 589718 454294
rect 589098 454170 589194 454226
rect 589250 454170 589318 454226
rect 589374 454170 589442 454226
rect 589498 454170 589566 454226
rect 589622 454170 589718 454226
rect 589098 454102 589718 454170
rect 589098 454046 589194 454102
rect 589250 454046 589318 454102
rect 589374 454046 589442 454102
rect 589498 454046 589566 454102
rect 589622 454046 589718 454102
rect 589098 453978 589718 454046
rect 589098 453922 589194 453978
rect 589250 453922 589318 453978
rect 589374 453922 589442 453978
rect 589498 453922 589566 453978
rect 589622 453922 589718 453978
rect 589098 436350 589718 453922
rect 589098 436294 589194 436350
rect 589250 436294 589318 436350
rect 589374 436294 589442 436350
rect 589498 436294 589566 436350
rect 589622 436294 589718 436350
rect 589098 436226 589718 436294
rect 589098 436170 589194 436226
rect 589250 436170 589318 436226
rect 589374 436170 589442 436226
rect 589498 436170 589566 436226
rect 589622 436170 589718 436226
rect 589098 436102 589718 436170
rect 589098 436046 589194 436102
rect 589250 436046 589318 436102
rect 589374 436046 589442 436102
rect 589498 436046 589566 436102
rect 589622 436046 589718 436102
rect 589098 435978 589718 436046
rect 589098 435922 589194 435978
rect 589250 435922 589318 435978
rect 589374 435922 589442 435978
rect 589498 435922 589566 435978
rect 589622 435922 589718 435978
rect 589098 418350 589718 435922
rect 589098 418294 589194 418350
rect 589250 418294 589318 418350
rect 589374 418294 589442 418350
rect 589498 418294 589566 418350
rect 589622 418294 589718 418350
rect 589098 418226 589718 418294
rect 589098 418170 589194 418226
rect 589250 418170 589318 418226
rect 589374 418170 589442 418226
rect 589498 418170 589566 418226
rect 589622 418170 589718 418226
rect 589098 418102 589718 418170
rect 589098 418046 589194 418102
rect 589250 418046 589318 418102
rect 589374 418046 589442 418102
rect 589498 418046 589566 418102
rect 589622 418046 589718 418102
rect 589098 417978 589718 418046
rect 589098 417922 589194 417978
rect 589250 417922 589318 417978
rect 589374 417922 589442 417978
rect 589498 417922 589566 417978
rect 589622 417922 589718 417978
rect 589098 400350 589718 417922
rect 589098 400294 589194 400350
rect 589250 400294 589318 400350
rect 589374 400294 589442 400350
rect 589498 400294 589566 400350
rect 589622 400294 589718 400350
rect 589098 400226 589718 400294
rect 589098 400170 589194 400226
rect 589250 400170 589318 400226
rect 589374 400170 589442 400226
rect 589498 400170 589566 400226
rect 589622 400170 589718 400226
rect 589098 400102 589718 400170
rect 589098 400046 589194 400102
rect 589250 400046 589318 400102
rect 589374 400046 589442 400102
rect 589498 400046 589566 400102
rect 589622 400046 589718 400102
rect 589098 399978 589718 400046
rect 589098 399922 589194 399978
rect 589250 399922 589318 399978
rect 589374 399922 589442 399978
rect 589498 399922 589566 399978
rect 589622 399922 589718 399978
rect 589098 382350 589718 399922
rect 589098 382294 589194 382350
rect 589250 382294 589318 382350
rect 589374 382294 589442 382350
rect 589498 382294 589566 382350
rect 589622 382294 589718 382350
rect 589098 382226 589718 382294
rect 589098 382170 589194 382226
rect 589250 382170 589318 382226
rect 589374 382170 589442 382226
rect 589498 382170 589566 382226
rect 589622 382170 589718 382226
rect 589098 382102 589718 382170
rect 589098 382046 589194 382102
rect 589250 382046 589318 382102
rect 589374 382046 589442 382102
rect 589498 382046 589566 382102
rect 589622 382046 589718 382102
rect 589098 381978 589718 382046
rect 589098 381922 589194 381978
rect 589250 381922 589318 381978
rect 589374 381922 589442 381978
rect 589498 381922 589566 381978
rect 589622 381922 589718 381978
rect 589098 364350 589718 381922
rect 589098 364294 589194 364350
rect 589250 364294 589318 364350
rect 589374 364294 589442 364350
rect 589498 364294 589566 364350
rect 589622 364294 589718 364350
rect 589098 364226 589718 364294
rect 589098 364170 589194 364226
rect 589250 364170 589318 364226
rect 589374 364170 589442 364226
rect 589498 364170 589566 364226
rect 589622 364170 589718 364226
rect 589098 364102 589718 364170
rect 589098 364046 589194 364102
rect 589250 364046 589318 364102
rect 589374 364046 589442 364102
rect 589498 364046 589566 364102
rect 589622 364046 589718 364102
rect 589098 363978 589718 364046
rect 589098 363922 589194 363978
rect 589250 363922 589318 363978
rect 589374 363922 589442 363978
rect 589498 363922 589566 363978
rect 589622 363922 589718 363978
rect 589098 346350 589718 363922
rect 589098 346294 589194 346350
rect 589250 346294 589318 346350
rect 589374 346294 589442 346350
rect 589498 346294 589566 346350
rect 589622 346294 589718 346350
rect 589098 346226 589718 346294
rect 589098 346170 589194 346226
rect 589250 346170 589318 346226
rect 589374 346170 589442 346226
rect 589498 346170 589566 346226
rect 589622 346170 589718 346226
rect 589098 346102 589718 346170
rect 589098 346046 589194 346102
rect 589250 346046 589318 346102
rect 589374 346046 589442 346102
rect 589498 346046 589566 346102
rect 589622 346046 589718 346102
rect 589098 345978 589718 346046
rect 589098 345922 589194 345978
rect 589250 345922 589318 345978
rect 589374 345922 589442 345978
rect 589498 345922 589566 345978
rect 589622 345922 589718 345978
rect 589098 328350 589718 345922
rect 589098 328294 589194 328350
rect 589250 328294 589318 328350
rect 589374 328294 589442 328350
rect 589498 328294 589566 328350
rect 589622 328294 589718 328350
rect 589098 328226 589718 328294
rect 589098 328170 589194 328226
rect 589250 328170 589318 328226
rect 589374 328170 589442 328226
rect 589498 328170 589566 328226
rect 589622 328170 589718 328226
rect 589098 328102 589718 328170
rect 589098 328046 589194 328102
rect 589250 328046 589318 328102
rect 589374 328046 589442 328102
rect 589498 328046 589566 328102
rect 589622 328046 589718 328102
rect 589098 327978 589718 328046
rect 589098 327922 589194 327978
rect 589250 327922 589318 327978
rect 589374 327922 589442 327978
rect 589498 327922 589566 327978
rect 589622 327922 589718 327978
rect 589098 310350 589718 327922
rect 589098 310294 589194 310350
rect 589250 310294 589318 310350
rect 589374 310294 589442 310350
rect 589498 310294 589566 310350
rect 589622 310294 589718 310350
rect 589098 310226 589718 310294
rect 589098 310170 589194 310226
rect 589250 310170 589318 310226
rect 589374 310170 589442 310226
rect 589498 310170 589566 310226
rect 589622 310170 589718 310226
rect 589098 310102 589718 310170
rect 589098 310046 589194 310102
rect 589250 310046 589318 310102
rect 589374 310046 589442 310102
rect 589498 310046 589566 310102
rect 589622 310046 589718 310102
rect 589098 309978 589718 310046
rect 589098 309922 589194 309978
rect 589250 309922 589318 309978
rect 589374 309922 589442 309978
rect 589498 309922 589566 309978
rect 589622 309922 589718 309978
rect 589098 292350 589718 309922
rect 589098 292294 589194 292350
rect 589250 292294 589318 292350
rect 589374 292294 589442 292350
rect 589498 292294 589566 292350
rect 589622 292294 589718 292350
rect 589098 292226 589718 292294
rect 589098 292170 589194 292226
rect 589250 292170 589318 292226
rect 589374 292170 589442 292226
rect 589498 292170 589566 292226
rect 589622 292170 589718 292226
rect 589098 292102 589718 292170
rect 589098 292046 589194 292102
rect 589250 292046 589318 292102
rect 589374 292046 589442 292102
rect 589498 292046 589566 292102
rect 589622 292046 589718 292102
rect 589098 291978 589718 292046
rect 589098 291922 589194 291978
rect 589250 291922 589318 291978
rect 589374 291922 589442 291978
rect 589498 291922 589566 291978
rect 589622 291922 589718 291978
rect 589098 274350 589718 291922
rect 589098 274294 589194 274350
rect 589250 274294 589318 274350
rect 589374 274294 589442 274350
rect 589498 274294 589566 274350
rect 589622 274294 589718 274350
rect 589098 274226 589718 274294
rect 589098 274170 589194 274226
rect 589250 274170 589318 274226
rect 589374 274170 589442 274226
rect 589498 274170 589566 274226
rect 589622 274170 589718 274226
rect 589098 274102 589718 274170
rect 589098 274046 589194 274102
rect 589250 274046 589318 274102
rect 589374 274046 589442 274102
rect 589498 274046 589566 274102
rect 589622 274046 589718 274102
rect 589098 273978 589718 274046
rect 589098 273922 589194 273978
rect 589250 273922 589318 273978
rect 589374 273922 589442 273978
rect 589498 273922 589566 273978
rect 589622 273922 589718 273978
rect 589098 256350 589718 273922
rect 589098 256294 589194 256350
rect 589250 256294 589318 256350
rect 589374 256294 589442 256350
rect 589498 256294 589566 256350
rect 589622 256294 589718 256350
rect 589098 256226 589718 256294
rect 589098 256170 589194 256226
rect 589250 256170 589318 256226
rect 589374 256170 589442 256226
rect 589498 256170 589566 256226
rect 589622 256170 589718 256226
rect 589098 256102 589718 256170
rect 589098 256046 589194 256102
rect 589250 256046 589318 256102
rect 589374 256046 589442 256102
rect 589498 256046 589566 256102
rect 589622 256046 589718 256102
rect 589098 255978 589718 256046
rect 589098 255922 589194 255978
rect 589250 255922 589318 255978
rect 589374 255922 589442 255978
rect 589498 255922 589566 255978
rect 589622 255922 589718 255978
rect 589098 238350 589718 255922
rect 589098 238294 589194 238350
rect 589250 238294 589318 238350
rect 589374 238294 589442 238350
rect 589498 238294 589566 238350
rect 589622 238294 589718 238350
rect 589098 238226 589718 238294
rect 589098 238170 589194 238226
rect 589250 238170 589318 238226
rect 589374 238170 589442 238226
rect 589498 238170 589566 238226
rect 589622 238170 589718 238226
rect 589098 238102 589718 238170
rect 589098 238046 589194 238102
rect 589250 238046 589318 238102
rect 589374 238046 589442 238102
rect 589498 238046 589566 238102
rect 589622 238046 589718 238102
rect 589098 237978 589718 238046
rect 589098 237922 589194 237978
rect 589250 237922 589318 237978
rect 589374 237922 589442 237978
rect 589498 237922 589566 237978
rect 589622 237922 589718 237978
rect 589098 220350 589718 237922
rect 589098 220294 589194 220350
rect 589250 220294 589318 220350
rect 589374 220294 589442 220350
rect 589498 220294 589566 220350
rect 589622 220294 589718 220350
rect 589098 220226 589718 220294
rect 589098 220170 589194 220226
rect 589250 220170 589318 220226
rect 589374 220170 589442 220226
rect 589498 220170 589566 220226
rect 589622 220170 589718 220226
rect 589098 220102 589718 220170
rect 589098 220046 589194 220102
rect 589250 220046 589318 220102
rect 589374 220046 589442 220102
rect 589498 220046 589566 220102
rect 589622 220046 589718 220102
rect 589098 219978 589718 220046
rect 589098 219922 589194 219978
rect 589250 219922 589318 219978
rect 589374 219922 589442 219978
rect 589498 219922 589566 219978
rect 589622 219922 589718 219978
rect 589098 202350 589718 219922
rect 589098 202294 589194 202350
rect 589250 202294 589318 202350
rect 589374 202294 589442 202350
rect 589498 202294 589566 202350
rect 589622 202294 589718 202350
rect 589098 202226 589718 202294
rect 589098 202170 589194 202226
rect 589250 202170 589318 202226
rect 589374 202170 589442 202226
rect 589498 202170 589566 202226
rect 589622 202170 589718 202226
rect 589098 202102 589718 202170
rect 589098 202046 589194 202102
rect 589250 202046 589318 202102
rect 589374 202046 589442 202102
rect 589498 202046 589566 202102
rect 589622 202046 589718 202102
rect 589098 201978 589718 202046
rect 589098 201922 589194 201978
rect 589250 201922 589318 201978
rect 589374 201922 589442 201978
rect 589498 201922 589566 201978
rect 589622 201922 589718 201978
rect 589098 184350 589718 201922
rect 589098 184294 589194 184350
rect 589250 184294 589318 184350
rect 589374 184294 589442 184350
rect 589498 184294 589566 184350
rect 589622 184294 589718 184350
rect 589098 184226 589718 184294
rect 589098 184170 589194 184226
rect 589250 184170 589318 184226
rect 589374 184170 589442 184226
rect 589498 184170 589566 184226
rect 589622 184170 589718 184226
rect 589098 184102 589718 184170
rect 589098 184046 589194 184102
rect 589250 184046 589318 184102
rect 589374 184046 589442 184102
rect 589498 184046 589566 184102
rect 589622 184046 589718 184102
rect 589098 183978 589718 184046
rect 589098 183922 589194 183978
rect 589250 183922 589318 183978
rect 589374 183922 589442 183978
rect 589498 183922 589566 183978
rect 589622 183922 589718 183978
rect 589098 166350 589718 183922
rect 589098 166294 589194 166350
rect 589250 166294 589318 166350
rect 589374 166294 589442 166350
rect 589498 166294 589566 166350
rect 589622 166294 589718 166350
rect 589098 166226 589718 166294
rect 589098 166170 589194 166226
rect 589250 166170 589318 166226
rect 589374 166170 589442 166226
rect 589498 166170 589566 166226
rect 589622 166170 589718 166226
rect 589098 166102 589718 166170
rect 589098 166046 589194 166102
rect 589250 166046 589318 166102
rect 589374 166046 589442 166102
rect 589498 166046 589566 166102
rect 589622 166046 589718 166102
rect 589098 165978 589718 166046
rect 589098 165922 589194 165978
rect 589250 165922 589318 165978
rect 589374 165922 589442 165978
rect 589498 165922 589566 165978
rect 589622 165922 589718 165978
rect 589098 148350 589718 165922
rect 589098 148294 589194 148350
rect 589250 148294 589318 148350
rect 589374 148294 589442 148350
rect 589498 148294 589566 148350
rect 589622 148294 589718 148350
rect 589098 148226 589718 148294
rect 589098 148170 589194 148226
rect 589250 148170 589318 148226
rect 589374 148170 589442 148226
rect 589498 148170 589566 148226
rect 589622 148170 589718 148226
rect 589098 148102 589718 148170
rect 589098 148046 589194 148102
rect 589250 148046 589318 148102
rect 589374 148046 589442 148102
rect 589498 148046 589566 148102
rect 589622 148046 589718 148102
rect 589098 147978 589718 148046
rect 589098 147922 589194 147978
rect 589250 147922 589318 147978
rect 589374 147922 589442 147978
rect 589498 147922 589566 147978
rect 589622 147922 589718 147978
rect 589098 130350 589718 147922
rect 589098 130294 589194 130350
rect 589250 130294 589318 130350
rect 589374 130294 589442 130350
rect 589498 130294 589566 130350
rect 589622 130294 589718 130350
rect 589098 130226 589718 130294
rect 589098 130170 589194 130226
rect 589250 130170 589318 130226
rect 589374 130170 589442 130226
rect 589498 130170 589566 130226
rect 589622 130170 589718 130226
rect 589098 130102 589718 130170
rect 589098 130046 589194 130102
rect 589250 130046 589318 130102
rect 589374 130046 589442 130102
rect 589498 130046 589566 130102
rect 589622 130046 589718 130102
rect 589098 129978 589718 130046
rect 589098 129922 589194 129978
rect 589250 129922 589318 129978
rect 589374 129922 589442 129978
rect 589498 129922 589566 129978
rect 589622 129922 589718 129978
rect 589098 112350 589718 129922
rect 589098 112294 589194 112350
rect 589250 112294 589318 112350
rect 589374 112294 589442 112350
rect 589498 112294 589566 112350
rect 589622 112294 589718 112350
rect 589098 112226 589718 112294
rect 589098 112170 589194 112226
rect 589250 112170 589318 112226
rect 589374 112170 589442 112226
rect 589498 112170 589566 112226
rect 589622 112170 589718 112226
rect 589098 112102 589718 112170
rect 589098 112046 589194 112102
rect 589250 112046 589318 112102
rect 589374 112046 589442 112102
rect 589498 112046 589566 112102
rect 589622 112046 589718 112102
rect 589098 111978 589718 112046
rect 589098 111922 589194 111978
rect 589250 111922 589318 111978
rect 589374 111922 589442 111978
rect 589498 111922 589566 111978
rect 589622 111922 589718 111978
rect 589098 94350 589718 111922
rect 589098 94294 589194 94350
rect 589250 94294 589318 94350
rect 589374 94294 589442 94350
rect 589498 94294 589566 94350
rect 589622 94294 589718 94350
rect 589098 94226 589718 94294
rect 589098 94170 589194 94226
rect 589250 94170 589318 94226
rect 589374 94170 589442 94226
rect 589498 94170 589566 94226
rect 589622 94170 589718 94226
rect 589098 94102 589718 94170
rect 589098 94046 589194 94102
rect 589250 94046 589318 94102
rect 589374 94046 589442 94102
rect 589498 94046 589566 94102
rect 589622 94046 589718 94102
rect 589098 93978 589718 94046
rect 589098 93922 589194 93978
rect 589250 93922 589318 93978
rect 589374 93922 589442 93978
rect 589498 93922 589566 93978
rect 589622 93922 589718 93978
rect 589098 76350 589718 93922
rect 589098 76294 589194 76350
rect 589250 76294 589318 76350
rect 589374 76294 589442 76350
rect 589498 76294 589566 76350
rect 589622 76294 589718 76350
rect 589098 76226 589718 76294
rect 589098 76170 589194 76226
rect 589250 76170 589318 76226
rect 589374 76170 589442 76226
rect 589498 76170 589566 76226
rect 589622 76170 589718 76226
rect 589098 76102 589718 76170
rect 589098 76046 589194 76102
rect 589250 76046 589318 76102
rect 589374 76046 589442 76102
rect 589498 76046 589566 76102
rect 589622 76046 589718 76102
rect 589098 75978 589718 76046
rect 589098 75922 589194 75978
rect 589250 75922 589318 75978
rect 589374 75922 589442 75978
rect 589498 75922 589566 75978
rect 589622 75922 589718 75978
rect 589098 58350 589718 75922
rect 589098 58294 589194 58350
rect 589250 58294 589318 58350
rect 589374 58294 589442 58350
rect 589498 58294 589566 58350
rect 589622 58294 589718 58350
rect 589098 58226 589718 58294
rect 589098 58170 589194 58226
rect 589250 58170 589318 58226
rect 589374 58170 589442 58226
rect 589498 58170 589566 58226
rect 589622 58170 589718 58226
rect 589098 58102 589718 58170
rect 589098 58046 589194 58102
rect 589250 58046 589318 58102
rect 589374 58046 589442 58102
rect 589498 58046 589566 58102
rect 589622 58046 589718 58102
rect 589098 57978 589718 58046
rect 589098 57922 589194 57978
rect 589250 57922 589318 57978
rect 589374 57922 589442 57978
rect 589498 57922 589566 57978
rect 589622 57922 589718 57978
rect 589098 40350 589718 57922
rect 589098 40294 589194 40350
rect 589250 40294 589318 40350
rect 589374 40294 589442 40350
rect 589498 40294 589566 40350
rect 589622 40294 589718 40350
rect 589098 40226 589718 40294
rect 589098 40170 589194 40226
rect 589250 40170 589318 40226
rect 589374 40170 589442 40226
rect 589498 40170 589566 40226
rect 589622 40170 589718 40226
rect 589098 40102 589718 40170
rect 589098 40046 589194 40102
rect 589250 40046 589318 40102
rect 589374 40046 589442 40102
rect 589498 40046 589566 40102
rect 589622 40046 589718 40102
rect 589098 39978 589718 40046
rect 589098 39922 589194 39978
rect 589250 39922 589318 39978
rect 589374 39922 589442 39978
rect 589498 39922 589566 39978
rect 589622 39922 589718 39978
rect 562098 28294 562194 28350
rect 562250 28294 562318 28350
rect 562374 28294 562442 28350
rect 562498 28294 562566 28350
rect 562622 28294 562718 28350
rect 562098 28226 562718 28294
rect 562098 28170 562194 28226
rect 562250 28170 562318 28226
rect 562374 28170 562442 28226
rect 562498 28170 562566 28226
rect 562622 28170 562718 28226
rect 562098 28102 562718 28170
rect 562098 28046 562194 28102
rect 562250 28046 562318 28102
rect 562374 28046 562442 28102
rect 562498 28046 562566 28102
rect 562622 28046 562718 28102
rect 562098 27978 562718 28046
rect 562098 27922 562194 27978
rect 562250 27922 562318 27978
rect 562374 27922 562442 27978
rect 562498 27922 562566 27978
rect 562622 27922 562718 27978
rect 562098 10350 562718 27922
rect 562098 10294 562194 10350
rect 562250 10294 562318 10350
rect 562374 10294 562442 10350
rect 562498 10294 562566 10350
rect 562622 10294 562718 10350
rect 562098 10226 562718 10294
rect 562098 10170 562194 10226
rect 562250 10170 562318 10226
rect 562374 10170 562442 10226
rect 562498 10170 562566 10226
rect 562622 10170 562718 10226
rect 562098 10102 562718 10170
rect 562098 10046 562194 10102
rect 562250 10046 562318 10102
rect 562374 10046 562442 10102
rect 562498 10046 562566 10102
rect 562622 10046 562718 10102
rect 562098 9978 562718 10046
rect 562098 9922 562194 9978
rect 562250 9922 562318 9978
rect 562374 9922 562442 9978
rect 562498 9922 562566 9978
rect 562622 9922 562718 9978
rect 562098 -1120 562718 9922
rect 562098 -1176 562194 -1120
rect 562250 -1176 562318 -1120
rect 562374 -1176 562442 -1120
rect 562498 -1176 562566 -1120
rect 562622 -1176 562718 -1120
rect 562098 -1244 562718 -1176
rect 562098 -1300 562194 -1244
rect 562250 -1300 562318 -1244
rect 562374 -1300 562442 -1244
rect 562498 -1300 562566 -1244
rect 562622 -1300 562718 -1244
rect 562098 -1368 562718 -1300
rect 562098 -1424 562194 -1368
rect 562250 -1424 562318 -1368
rect 562374 -1424 562442 -1368
rect 562498 -1424 562566 -1368
rect 562622 -1424 562718 -1368
rect 562098 -1492 562718 -1424
rect 562098 -1548 562194 -1492
rect 562250 -1548 562318 -1492
rect 562374 -1548 562442 -1492
rect 562498 -1548 562566 -1492
rect 562622 -1548 562718 -1492
rect 562098 -1644 562718 -1548
rect 589098 22350 589718 39922
rect 589098 22294 589194 22350
rect 589250 22294 589318 22350
rect 589374 22294 589442 22350
rect 589498 22294 589566 22350
rect 589622 22294 589718 22350
rect 589098 22226 589718 22294
rect 589098 22170 589194 22226
rect 589250 22170 589318 22226
rect 589374 22170 589442 22226
rect 589498 22170 589566 22226
rect 589622 22170 589718 22226
rect 589098 22102 589718 22170
rect 589098 22046 589194 22102
rect 589250 22046 589318 22102
rect 589374 22046 589442 22102
rect 589498 22046 589566 22102
rect 589622 22046 589718 22102
rect 589098 21978 589718 22046
rect 589098 21922 589194 21978
rect 589250 21922 589318 21978
rect 589374 21922 589442 21978
rect 589498 21922 589566 21978
rect 589622 21922 589718 21978
rect 589098 4350 589718 21922
rect 589098 4294 589194 4350
rect 589250 4294 589318 4350
rect 589374 4294 589442 4350
rect 589498 4294 589566 4350
rect 589622 4294 589718 4350
rect 589098 4226 589718 4294
rect 589098 4170 589194 4226
rect 589250 4170 589318 4226
rect 589374 4170 589442 4226
rect 589498 4170 589566 4226
rect 589622 4170 589718 4226
rect 589098 4102 589718 4170
rect 589098 4046 589194 4102
rect 589250 4046 589318 4102
rect 589374 4046 589442 4102
rect 589498 4046 589566 4102
rect 589622 4046 589718 4102
rect 589098 3978 589718 4046
rect 589098 3922 589194 3978
rect 589250 3922 589318 3978
rect 589374 3922 589442 3978
rect 589498 3922 589566 3978
rect 589622 3922 589718 3978
rect 589098 -160 589718 3922
rect 589098 -216 589194 -160
rect 589250 -216 589318 -160
rect 589374 -216 589442 -160
rect 589498 -216 589566 -160
rect 589622 -216 589718 -160
rect 589098 -284 589718 -216
rect 589098 -340 589194 -284
rect 589250 -340 589318 -284
rect 589374 -340 589442 -284
rect 589498 -340 589566 -284
rect 589622 -340 589718 -284
rect 589098 -408 589718 -340
rect 589098 -464 589194 -408
rect 589250 -464 589318 -408
rect 589374 -464 589442 -408
rect 589498 -464 589566 -408
rect 589622 -464 589718 -408
rect 589098 -532 589718 -464
rect 589098 -588 589194 -532
rect 589250 -588 589318 -532
rect 589374 -588 589442 -532
rect 589498 -588 589566 -532
rect 589622 -588 589718 -532
rect 589098 -1644 589718 -588
rect 592818 598172 593438 598268
rect 592818 598116 592914 598172
rect 592970 598116 593038 598172
rect 593094 598116 593162 598172
rect 593218 598116 593286 598172
rect 593342 598116 593438 598172
rect 592818 598048 593438 598116
rect 592818 597992 592914 598048
rect 592970 597992 593038 598048
rect 593094 597992 593162 598048
rect 593218 597992 593286 598048
rect 593342 597992 593438 598048
rect 592818 597924 593438 597992
rect 592818 597868 592914 597924
rect 592970 597868 593038 597924
rect 593094 597868 593162 597924
rect 593218 597868 593286 597924
rect 593342 597868 593438 597924
rect 592818 597800 593438 597868
rect 592818 597744 592914 597800
rect 592970 597744 593038 597800
rect 593094 597744 593162 597800
rect 593218 597744 593286 597800
rect 593342 597744 593438 597800
rect 592818 586350 593438 597744
rect 597360 598172 597980 598268
rect 597360 598116 597456 598172
rect 597512 598116 597580 598172
rect 597636 598116 597704 598172
rect 597760 598116 597828 598172
rect 597884 598116 597980 598172
rect 597360 598048 597980 598116
rect 597360 597992 597456 598048
rect 597512 597992 597580 598048
rect 597636 597992 597704 598048
rect 597760 597992 597828 598048
rect 597884 597992 597980 598048
rect 597360 597924 597980 597992
rect 597360 597868 597456 597924
rect 597512 597868 597580 597924
rect 597636 597868 597704 597924
rect 597760 597868 597828 597924
rect 597884 597868 597980 597924
rect 597360 597800 597980 597868
rect 597360 597744 597456 597800
rect 597512 597744 597580 597800
rect 597636 597744 597704 597800
rect 597760 597744 597828 597800
rect 597884 597744 597980 597800
rect 592818 586294 592914 586350
rect 592970 586294 593038 586350
rect 593094 586294 593162 586350
rect 593218 586294 593286 586350
rect 593342 586294 593438 586350
rect 592818 586226 593438 586294
rect 592818 586170 592914 586226
rect 592970 586170 593038 586226
rect 593094 586170 593162 586226
rect 593218 586170 593286 586226
rect 593342 586170 593438 586226
rect 592818 586102 593438 586170
rect 592818 586046 592914 586102
rect 592970 586046 593038 586102
rect 593094 586046 593162 586102
rect 593218 586046 593286 586102
rect 593342 586046 593438 586102
rect 592818 585978 593438 586046
rect 592818 585922 592914 585978
rect 592970 585922 593038 585978
rect 593094 585922 593162 585978
rect 593218 585922 593286 585978
rect 593342 585922 593438 585978
rect 592818 568350 593438 585922
rect 592818 568294 592914 568350
rect 592970 568294 593038 568350
rect 593094 568294 593162 568350
rect 593218 568294 593286 568350
rect 593342 568294 593438 568350
rect 592818 568226 593438 568294
rect 592818 568170 592914 568226
rect 592970 568170 593038 568226
rect 593094 568170 593162 568226
rect 593218 568170 593286 568226
rect 593342 568170 593438 568226
rect 592818 568102 593438 568170
rect 592818 568046 592914 568102
rect 592970 568046 593038 568102
rect 593094 568046 593162 568102
rect 593218 568046 593286 568102
rect 593342 568046 593438 568102
rect 592818 567978 593438 568046
rect 592818 567922 592914 567978
rect 592970 567922 593038 567978
rect 593094 567922 593162 567978
rect 593218 567922 593286 567978
rect 593342 567922 593438 567978
rect 592818 550350 593438 567922
rect 592818 550294 592914 550350
rect 592970 550294 593038 550350
rect 593094 550294 593162 550350
rect 593218 550294 593286 550350
rect 593342 550294 593438 550350
rect 592818 550226 593438 550294
rect 592818 550170 592914 550226
rect 592970 550170 593038 550226
rect 593094 550170 593162 550226
rect 593218 550170 593286 550226
rect 593342 550170 593438 550226
rect 592818 550102 593438 550170
rect 592818 550046 592914 550102
rect 592970 550046 593038 550102
rect 593094 550046 593162 550102
rect 593218 550046 593286 550102
rect 593342 550046 593438 550102
rect 592818 549978 593438 550046
rect 592818 549922 592914 549978
rect 592970 549922 593038 549978
rect 593094 549922 593162 549978
rect 593218 549922 593286 549978
rect 593342 549922 593438 549978
rect 592818 532350 593438 549922
rect 592818 532294 592914 532350
rect 592970 532294 593038 532350
rect 593094 532294 593162 532350
rect 593218 532294 593286 532350
rect 593342 532294 593438 532350
rect 592818 532226 593438 532294
rect 592818 532170 592914 532226
rect 592970 532170 593038 532226
rect 593094 532170 593162 532226
rect 593218 532170 593286 532226
rect 593342 532170 593438 532226
rect 592818 532102 593438 532170
rect 592818 532046 592914 532102
rect 592970 532046 593038 532102
rect 593094 532046 593162 532102
rect 593218 532046 593286 532102
rect 593342 532046 593438 532102
rect 592818 531978 593438 532046
rect 592818 531922 592914 531978
rect 592970 531922 593038 531978
rect 593094 531922 593162 531978
rect 593218 531922 593286 531978
rect 593342 531922 593438 531978
rect 592818 514350 593438 531922
rect 592818 514294 592914 514350
rect 592970 514294 593038 514350
rect 593094 514294 593162 514350
rect 593218 514294 593286 514350
rect 593342 514294 593438 514350
rect 592818 514226 593438 514294
rect 592818 514170 592914 514226
rect 592970 514170 593038 514226
rect 593094 514170 593162 514226
rect 593218 514170 593286 514226
rect 593342 514170 593438 514226
rect 592818 514102 593438 514170
rect 592818 514046 592914 514102
rect 592970 514046 593038 514102
rect 593094 514046 593162 514102
rect 593218 514046 593286 514102
rect 593342 514046 593438 514102
rect 592818 513978 593438 514046
rect 592818 513922 592914 513978
rect 592970 513922 593038 513978
rect 593094 513922 593162 513978
rect 593218 513922 593286 513978
rect 593342 513922 593438 513978
rect 592818 496350 593438 513922
rect 592818 496294 592914 496350
rect 592970 496294 593038 496350
rect 593094 496294 593162 496350
rect 593218 496294 593286 496350
rect 593342 496294 593438 496350
rect 592818 496226 593438 496294
rect 592818 496170 592914 496226
rect 592970 496170 593038 496226
rect 593094 496170 593162 496226
rect 593218 496170 593286 496226
rect 593342 496170 593438 496226
rect 592818 496102 593438 496170
rect 592818 496046 592914 496102
rect 592970 496046 593038 496102
rect 593094 496046 593162 496102
rect 593218 496046 593286 496102
rect 593342 496046 593438 496102
rect 592818 495978 593438 496046
rect 592818 495922 592914 495978
rect 592970 495922 593038 495978
rect 593094 495922 593162 495978
rect 593218 495922 593286 495978
rect 593342 495922 593438 495978
rect 592818 478350 593438 495922
rect 592818 478294 592914 478350
rect 592970 478294 593038 478350
rect 593094 478294 593162 478350
rect 593218 478294 593286 478350
rect 593342 478294 593438 478350
rect 592818 478226 593438 478294
rect 592818 478170 592914 478226
rect 592970 478170 593038 478226
rect 593094 478170 593162 478226
rect 593218 478170 593286 478226
rect 593342 478170 593438 478226
rect 592818 478102 593438 478170
rect 592818 478046 592914 478102
rect 592970 478046 593038 478102
rect 593094 478046 593162 478102
rect 593218 478046 593286 478102
rect 593342 478046 593438 478102
rect 592818 477978 593438 478046
rect 592818 477922 592914 477978
rect 592970 477922 593038 477978
rect 593094 477922 593162 477978
rect 593218 477922 593286 477978
rect 593342 477922 593438 477978
rect 592818 460350 593438 477922
rect 592818 460294 592914 460350
rect 592970 460294 593038 460350
rect 593094 460294 593162 460350
rect 593218 460294 593286 460350
rect 593342 460294 593438 460350
rect 592818 460226 593438 460294
rect 592818 460170 592914 460226
rect 592970 460170 593038 460226
rect 593094 460170 593162 460226
rect 593218 460170 593286 460226
rect 593342 460170 593438 460226
rect 592818 460102 593438 460170
rect 592818 460046 592914 460102
rect 592970 460046 593038 460102
rect 593094 460046 593162 460102
rect 593218 460046 593286 460102
rect 593342 460046 593438 460102
rect 592818 459978 593438 460046
rect 592818 459922 592914 459978
rect 592970 459922 593038 459978
rect 593094 459922 593162 459978
rect 593218 459922 593286 459978
rect 593342 459922 593438 459978
rect 592818 442350 593438 459922
rect 592818 442294 592914 442350
rect 592970 442294 593038 442350
rect 593094 442294 593162 442350
rect 593218 442294 593286 442350
rect 593342 442294 593438 442350
rect 592818 442226 593438 442294
rect 592818 442170 592914 442226
rect 592970 442170 593038 442226
rect 593094 442170 593162 442226
rect 593218 442170 593286 442226
rect 593342 442170 593438 442226
rect 592818 442102 593438 442170
rect 592818 442046 592914 442102
rect 592970 442046 593038 442102
rect 593094 442046 593162 442102
rect 593218 442046 593286 442102
rect 593342 442046 593438 442102
rect 592818 441978 593438 442046
rect 592818 441922 592914 441978
rect 592970 441922 593038 441978
rect 593094 441922 593162 441978
rect 593218 441922 593286 441978
rect 593342 441922 593438 441978
rect 592818 424350 593438 441922
rect 592818 424294 592914 424350
rect 592970 424294 593038 424350
rect 593094 424294 593162 424350
rect 593218 424294 593286 424350
rect 593342 424294 593438 424350
rect 592818 424226 593438 424294
rect 592818 424170 592914 424226
rect 592970 424170 593038 424226
rect 593094 424170 593162 424226
rect 593218 424170 593286 424226
rect 593342 424170 593438 424226
rect 592818 424102 593438 424170
rect 592818 424046 592914 424102
rect 592970 424046 593038 424102
rect 593094 424046 593162 424102
rect 593218 424046 593286 424102
rect 593342 424046 593438 424102
rect 592818 423978 593438 424046
rect 592818 423922 592914 423978
rect 592970 423922 593038 423978
rect 593094 423922 593162 423978
rect 593218 423922 593286 423978
rect 593342 423922 593438 423978
rect 592818 406350 593438 423922
rect 592818 406294 592914 406350
rect 592970 406294 593038 406350
rect 593094 406294 593162 406350
rect 593218 406294 593286 406350
rect 593342 406294 593438 406350
rect 592818 406226 593438 406294
rect 592818 406170 592914 406226
rect 592970 406170 593038 406226
rect 593094 406170 593162 406226
rect 593218 406170 593286 406226
rect 593342 406170 593438 406226
rect 592818 406102 593438 406170
rect 592818 406046 592914 406102
rect 592970 406046 593038 406102
rect 593094 406046 593162 406102
rect 593218 406046 593286 406102
rect 593342 406046 593438 406102
rect 592818 405978 593438 406046
rect 592818 405922 592914 405978
rect 592970 405922 593038 405978
rect 593094 405922 593162 405978
rect 593218 405922 593286 405978
rect 593342 405922 593438 405978
rect 592818 388350 593438 405922
rect 592818 388294 592914 388350
rect 592970 388294 593038 388350
rect 593094 388294 593162 388350
rect 593218 388294 593286 388350
rect 593342 388294 593438 388350
rect 592818 388226 593438 388294
rect 592818 388170 592914 388226
rect 592970 388170 593038 388226
rect 593094 388170 593162 388226
rect 593218 388170 593286 388226
rect 593342 388170 593438 388226
rect 592818 388102 593438 388170
rect 592818 388046 592914 388102
rect 592970 388046 593038 388102
rect 593094 388046 593162 388102
rect 593218 388046 593286 388102
rect 593342 388046 593438 388102
rect 592818 387978 593438 388046
rect 592818 387922 592914 387978
rect 592970 387922 593038 387978
rect 593094 387922 593162 387978
rect 593218 387922 593286 387978
rect 593342 387922 593438 387978
rect 592818 370350 593438 387922
rect 592818 370294 592914 370350
rect 592970 370294 593038 370350
rect 593094 370294 593162 370350
rect 593218 370294 593286 370350
rect 593342 370294 593438 370350
rect 592818 370226 593438 370294
rect 592818 370170 592914 370226
rect 592970 370170 593038 370226
rect 593094 370170 593162 370226
rect 593218 370170 593286 370226
rect 593342 370170 593438 370226
rect 592818 370102 593438 370170
rect 592818 370046 592914 370102
rect 592970 370046 593038 370102
rect 593094 370046 593162 370102
rect 593218 370046 593286 370102
rect 593342 370046 593438 370102
rect 592818 369978 593438 370046
rect 592818 369922 592914 369978
rect 592970 369922 593038 369978
rect 593094 369922 593162 369978
rect 593218 369922 593286 369978
rect 593342 369922 593438 369978
rect 592818 352350 593438 369922
rect 592818 352294 592914 352350
rect 592970 352294 593038 352350
rect 593094 352294 593162 352350
rect 593218 352294 593286 352350
rect 593342 352294 593438 352350
rect 592818 352226 593438 352294
rect 592818 352170 592914 352226
rect 592970 352170 593038 352226
rect 593094 352170 593162 352226
rect 593218 352170 593286 352226
rect 593342 352170 593438 352226
rect 592818 352102 593438 352170
rect 592818 352046 592914 352102
rect 592970 352046 593038 352102
rect 593094 352046 593162 352102
rect 593218 352046 593286 352102
rect 593342 352046 593438 352102
rect 592818 351978 593438 352046
rect 592818 351922 592914 351978
rect 592970 351922 593038 351978
rect 593094 351922 593162 351978
rect 593218 351922 593286 351978
rect 593342 351922 593438 351978
rect 592818 334350 593438 351922
rect 592818 334294 592914 334350
rect 592970 334294 593038 334350
rect 593094 334294 593162 334350
rect 593218 334294 593286 334350
rect 593342 334294 593438 334350
rect 592818 334226 593438 334294
rect 592818 334170 592914 334226
rect 592970 334170 593038 334226
rect 593094 334170 593162 334226
rect 593218 334170 593286 334226
rect 593342 334170 593438 334226
rect 592818 334102 593438 334170
rect 592818 334046 592914 334102
rect 592970 334046 593038 334102
rect 593094 334046 593162 334102
rect 593218 334046 593286 334102
rect 593342 334046 593438 334102
rect 592818 333978 593438 334046
rect 592818 333922 592914 333978
rect 592970 333922 593038 333978
rect 593094 333922 593162 333978
rect 593218 333922 593286 333978
rect 593342 333922 593438 333978
rect 592818 316350 593438 333922
rect 592818 316294 592914 316350
rect 592970 316294 593038 316350
rect 593094 316294 593162 316350
rect 593218 316294 593286 316350
rect 593342 316294 593438 316350
rect 592818 316226 593438 316294
rect 592818 316170 592914 316226
rect 592970 316170 593038 316226
rect 593094 316170 593162 316226
rect 593218 316170 593286 316226
rect 593342 316170 593438 316226
rect 592818 316102 593438 316170
rect 592818 316046 592914 316102
rect 592970 316046 593038 316102
rect 593094 316046 593162 316102
rect 593218 316046 593286 316102
rect 593342 316046 593438 316102
rect 592818 315978 593438 316046
rect 592818 315922 592914 315978
rect 592970 315922 593038 315978
rect 593094 315922 593162 315978
rect 593218 315922 593286 315978
rect 593342 315922 593438 315978
rect 592818 298350 593438 315922
rect 592818 298294 592914 298350
rect 592970 298294 593038 298350
rect 593094 298294 593162 298350
rect 593218 298294 593286 298350
rect 593342 298294 593438 298350
rect 592818 298226 593438 298294
rect 592818 298170 592914 298226
rect 592970 298170 593038 298226
rect 593094 298170 593162 298226
rect 593218 298170 593286 298226
rect 593342 298170 593438 298226
rect 592818 298102 593438 298170
rect 592818 298046 592914 298102
rect 592970 298046 593038 298102
rect 593094 298046 593162 298102
rect 593218 298046 593286 298102
rect 593342 298046 593438 298102
rect 592818 297978 593438 298046
rect 592818 297922 592914 297978
rect 592970 297922 593038 297978
rect 593094 297922 593162 297978
rect 593218 297922 593286 297978
rect 593342 297922 593438 297978
rect 592818 280350 593438 297922
rect 592818 280294 592914 280350
rect 592970 280294 593038 280350
rect 593094 280294 593162 280350
rect 593218 280294 593286 280350
rect 593342 280294 593438 280350
rect 592818 280226 593438 280294
rect 592818 280170 592914 280226
rect 592970 280170 593038 280226
rect 593094 280170 593162 280226
rect 593218 280170 593286 280226
rect 593342 280170 593438 280226
rect 592818 280102 593438 280170
rect 592818 280046 592914 280102
rect 592970 280046 593038 280102
rect 593094 280046 593162 280102
rect 593218 280046 593286 280102
rect 593342 280046 593438 280102
rect 592818 279978 593438 280046
rect 592818 279922 592914 279978
rect 592970 279922 593038 279978
rect 593094 279922 593162 279978
rect 593218 279922 593286 279978
rect 593342 279922 593438 279978
rect 592818 262350 593438 279922
rect 592818 262294 592914 262350
rect 592970 262294 593038 262350
rect 593094 262294 593162 262350
rect 593218 262294 593286 262350
rect 593342 262294 593438 262350
rect 592818 262226 593438 262294
rect 592818 262170 592914 262226
rect 592970 262170 593038 262226
rect 593094 262170 593162 262226
rect 593218 262170 593286 262226
rect 593342 262170 593438 262226
rect 592818 262102 593438 262170
rect 592818 262046 592914 262102
rect 592970 262046 593038 262102
rect 593094 262046 593162 262102
rect 593218 262046 593286 262102
rect 593342 262046 593438 262102
rect 592818 261978 593438 262046
rect 592818 261922 592914 261978
rect 592970 261922 593038 261978
rect 593094 261922 593162 261978
rect 593218 261922 593286 261978
rect 593342 261922 593438 261978
rect 592818 244350 593438 261922
rect 592818 244294 592914 244350
rect 592970 244294 593038 244350
rect 593094 244294 593162 244350
rect 593218 244294 593286 244350
rect 593342 244294 593438 244350
rect 592818 244226 593438 244294
rect 592818 244170 592914 244226
rect 592970 244170 593038 244226
rect 593094 244170 593162 244226
rect 593218 244170 593286 244226
rect 593342 244170 593438 244226
rect 592818 244102 593438 244170
rect 592818 244046 592914 244102
rect 592970 244046 593038 244102
rect 593094 244046 593162 244102
rect 593218 244046 593286 244102
rect 593342 244046 593438 244102
rect 592818 243978 593438 244046
rect 592818 243922 592914 243978
rect 592970 243922 593038 243978
rect 593094 243922 593162 243978
rect 593218 243922 593286 243978
rect 593342 243922 593438 243978
rect 592818 226350 593438 243922
rect 592818 226294 592914 226350
rect 592970 226294 593038 226350
rect 593094 226294 593162 226350
rect 593218 226294 593286 226350
rect 593342 226294 593438 226350
rect 592818 226226 593438 226294
rect 592818 226170 592914 226226
rect 592970 226170 593038 226226
rect 593094 226170 593162 226226
rect 593218 226170 593286 226226
rect 593342 226170 593438 226226
rect 592818 226102 593438 226170
rect 592818 226046 592914 226102
rect 592970 226046 593038 226102
rect 593094 226046 593162 226102
rect 593218 226046 593286 226102
rect 593342 226046 593438 226102
rect 592818 225978 593438 226046
rect 592818 225922 592914 225978
rect 592970 225922 593038 225978
rect 593094 225922 593162 225978
rect 593218 225922 593286 225978
rect 593342 225922 593438 225978
rect 592818 208350 593438 225922
rect 592818 208294 592914 208350
rect 592970 208294 593038 208350
rect 593094 208294 593162 208350
rect 593218 208294 593286 208350
rect 593342 208294 593438 208350
rect 592818 208226 593438 208294
rect 592818 208170 592914 208226
rect 592970 208170 593038 208226
rect 593094 208170 593162 208226
rect 593218 208170 593286 208226
rect 593342 208170 593438 208226
rect 592818 208102 593438 208170
rect 592818 208046 592914 208102
rect 592970 208046 593038 208102
rect 593094 208046 593162 208102
rect 593218 208046 593286 208102
rect 593342 208046 593438 208102
rect 592818 207978 593438 208046
rect 592818 207922 592914 207978
rect 592970 207922 593038 207978
rect 593094 207922 593162 207978
rect 593218 207922 593286 207978
rect 593342 207922 593438 207978
rect 592818 190350 593438 207922
rect 592818 190294 592914 190350
rect 592970 190294 593038 190350
rect 593094 190294 593162 190350
rect 593218 190294 593286 190350
rect 593342 190294 593438 190350
rect 592818 190226 593438 190294
rect 592818 190170 592914 190226
rect 592970 190170 593038 190226
rect 593094 190170 593162 190226
rect 593218 190170 593286 190226
rect 593342 190170 593438 190226
rect 592818 190102 593438 190170
rect 592818 190046 592914 190102
rect 592970 190046 593038 190102
rect 593094 190046 593162 190102
rect 593218 190046 593286 190102
rect 593342 190046 593438 190102
rect 592818 189978 593438 190046
rect 592818 189922 592914 189978
rect 592970 189922 593038 189978
rect 593094 189922 593162 189978
rect 593218 189922 593286 189978
rect 593342 189922 593438 189978
rect 592818 172350 593438 189922
rect 592818 172294 592914 172350
rect 592970 172294 593038 172350
rect 593094 172294 593162 172350
rect 593218 172294 593286 172350
rect 593342 172294 593438 172350
rect 592818 172226 593438 172294
rect 592818 172170 592914 172226
rect 592970 172170 593038 172226
rect 593094 172170 593162 172226
rect 593218 172170 593286 172226
rect 593342 172170 593438 172226
rect 592818 172102 593438 172170
rect 592818 172046 592914 172102
rect 592970 172046 593038 172102
rect 593094 172046 593162 172102
rect 593218 172046 593286 172102
rect 593342 172046 593438 172102
rect 592818 171978 593438 172046
rect 592818 171922 592914 171978
rect 592970 171922 593038 171978
rect 593094 171922 593162 171978
rect 593218 171922 593286 171978
rect 593342 171922 593438 171978
rect 592818 154350 593438 171922
rect 592818 154294 592914 154350
rect 592970 154294 593038 154350
rect 593094 154294 593162 154350
rect 593218 154294 593286 154350
rect 593342 154294 593438 154350
rect 592818 154226 593438 154294
rect 592818 154170 592914 154226
rect 592970 154170 593038 154226
rect 593094 154170 593162 154226
rect 593218 154170 593286 154226
rect 593342 154170 593438 154226
rect 592818 154102 593438 154170
rect 592818 154046 592914 154102
rect 592970 154046 593038 154102
rect 593094 154046 593162 154102
rect 593218 154046 593286 154102
rect 593342 154046 593438 154102
rect 592818 153978 593438 154046
rect 592818 153922 592914 153978
rect 592970 153922 593038 153978
rect 593094 153922 593162 153978
rect 593218 153922 593286 153978
rect 593342 153922 593438 153978
rect 592818 136350 593438 153922
rect 592818 136294 592914 136350
rect 592970 136294 593038 136350
rect 593094 136294 593162 136350
rect 593218 136294 593286 136350
rect 593342 136294 593438 136350
rect 592818 136226 593438 136294
rect 592818 136170 592914 136226
rect 592970 136170 593038 136226
rect 593094 136170 593162 136226
rect 593218 136170 593286 136226
rect 593342 136170 593438 136226
rect 592818 136102 593438 136170
rect 592818 136046 592914 136102
rect 592970 136046 593038 136102
rect 593094 136046 593162 136102
rect 593218 136046 593286 136102
rect 593342 136046 593438 136102
rect 592818 135978 593438 136046
rect 592818 135922 592914 135978
rect 592970 135922 593038 135978
rect 593094 135922 593162 135978
rect 593218 135922 593286 135978
rect 593342 135922 593438 135978
rect 592818 118350 593438 135922
rect 592818 118294 592914 118350
rect 592970 118294 593038 118350
rect 593094 118294 593162 118350
rect 593218 118294 593286 118350
rect 593342 118294 593438 118350
rect 592818 118226 593438 118294
rect 592818 118170 592914 118226
rect 592970 118170 593038 118226
rect 593094 118170 593162 118226
rect 593218 118170 593286 118226
rect 593342 118170 593438 118226
rect 592818 118102 593438 118170
rect 592818 118046 592914 118102
rect 592970 118046 593038 118102
rect 593094 118046 593162 118102
rect 593218 118046 593286 118102
rect 593342 118046 593438 118102
rect 592818 117978 593438 118046
rect 592818 117922 592914 117978
rect 592970 117922 593038 117978
rect 593094 117922 593162 117978
rect 593218 117922 593286 117978
rect 593342 117922 593438 117978
rect 592818 100350 593438 117922
rect 592818 100294 592914 100350
rect 592970 100294 593038 100350
rect 593094 100294 593162 100350
rect 593218 100294 593286 100350
rect 593342 100294 593438 100350
rect 592818 100226 593438 100294
rect 592818 100170 592914 100226
rect 592970 100170 593038 100226
rect 593094 100170 593162 100226
rect 593218 100170 593286 100226
rect 593342 100170 593438 100226
rect 592818 100102 593438 100170
rect 592818 100046 592914 100102
rect 592970 100046 593038 100102
rect 593094 100046 593162 100102
rect 593218 100046 593286 100102
rect 593342 100046 593438 100102
rect 592818 99978 593438 100046
rect 592818 99922 592914 99978
rect 592970 99922 593038 99978
rect 593094 99922 593162 99978
rect 593218 99922 593286 99978
rect 593342 99922 593438 99978
rect 592818 82350 593438 99922
rect 592818 82294 592914 82350
rect 592970 82294 593038 82350
rect 593094 82294 593162 82350
rect 593218 82294 593286 82350
rect 593342 82294 593438 82350
rect 592818 82226 593438 82294
rect 592818 82170 592914 82226
rect 592970 82170 593038 82226
rect 593094 82170 593162 82226
rect 593218 82170 593286 82226
rect 593342 82170 593438 82226
rect 592818 82102 593438 82170
rect 592818 82046 592914 82102
rect 592970 82046 593038 82102
rect 593094 82046 593162 82102
rect 593218 82046 593286 82102
rect 593342 82046 593438 82102
rect 592818 81978 593438 82046
rect 592818 81922 592914 81978
rect 592970 81922 593038 81978
rect 593094 81922 593162 81978
rect 593218 81922 593286 81978
rect 593342 81922 593438 81978
rect 592818 64350 593438 81922
rect 592818 64294 592914 64350
rect 592970 64294 593038 64350
rect 593094 64294 593162 64350
rect 593218 64294 593286 64350
rect 593342 64294 593438 64350
rect 592818 64226 593438 64294
rect 592818 64170 592914 64226
rect 592970 64170 593038 64226
rect 593094 64170 593162 64226
rect 593218 64170 593286 64226
rect 593342 64170 593438 64226
rect 592818 64102 593438 64170
rect 592818 64046 592914 64102
rect 592970 64046 593038 64102
rect 593094 64046 593162 64102
rect 593218 64046 593286 64102
rect 593342 64046 593438 64102
rect 592818 63978 593438 64046
rect 592818 63922 592914 63978
rect 592970 63922 593038 63978
rect 593094 63922 593162 63978
rect 593218 63922 593286 63978
rect 593342 63922 593438 63978
rect 592818 46350 593438 63922
rect 592818 46294 592914 46350
rect 592970 46294 593038 46350
rect 593094 46294 593162 46350
rect 593218 46294 593286 46350
rect 593342 46294 593438 46350
rect 592818 46226 593438 46294
rect 592818 46170 592914 46226
rect 592970 46170 593038 46226
rect 593094 46170 593162 46226
rect 593218 46170 593286 46226
rect 593342 46170 593438 46226
rect 592818 46102 593438 46170
rect 592818 46046 592914 46102
rect 592970 46046 593038 46102
rect 593094 46046 593162 46102
rect 593218 46046 593286 46102
rect 593342 46046 593438 46102
rect 592818 45978 593438 46046
rect 592818 45922 592914 45978
rect 592970 45922 593038 45978
rect 593094 45922 593162 45978
rect 593218 45922 593286 45978
rect 593342 45922 593438 45978
rect 592818 28350 593438 45922
rect 592818 28294 592914 28350
rect 592970 28294 593038 28350
rect 593094 28294 593162 28350
rect 593218 28294 593286 28350
rect 593342 28294 593438 28350
rect 592818 28226 593438 28294
rect 592818 28170 592914 28226
rect 592970 28170 593038 28226
rect 593094 28170 593162 28226
rect 593218 28170 593286 28226
rect 593342 28170 593438 28226
rect 592818 28102 593438 28170
rect 592818 28046 592914 28102
rect 592970 28046 593038 28102
rect 593094 28046 593162 28102
rect 593218 28046 593286 28102
rect 593342 28046 593438 28102
rect 592818 27978 593438 28046
rect 592818 27922 592914 27978
rect 592970 27922 593038 27978
rect 593094 27922 593162 27978
rect 593218 27922 593286 27978
rect 593342 27922 593438 27978
rect 592818 10350 593438 27922
rect 592818 10294 592914 10350
rect 592970 10294 593038 10350
rect 593094 10294 593162 10350
rect 593218 10294 593286 10350
rect 593342 10294 593438 10350
rect 592818 10226 593438 10294
rect 592818 10170 592914 10226
rect 592970 10170 593038 10226
rect 593094 10170 593162 10226
rect 593218 10170 593286 10226
rect 593342 10170 593438 10226
rect 592818 10102 593438 10170
rect 592818 10046 592914 10102
rect 592970 10046 593038 10102
rect 593094 10046 593162 10102
rect 593218 10046 593286 10102
rect 593342 10046 593438 10102
rect 592818 9978 593438 10046
rect 592818 9922 592914 9978
rect 592970 9922 593038 9978
rect 593094 9922 593162 9978
rect 593218 9922 593286 9978
rect 593342 9922 593438 9978
rect 592818 -1120 593438 9922
rect 596400 597212 597020 597308
rect 596400 597156 596496 597212
rect 596552 597156 596620 597212
rect 596676 597156 596744 597212
rect 596800 597156 596868 597212
rect 596924 597156 597020 597212
rect 596400 597088 597020 597156
rect 596400 597032 596496 597088
rect 596552 597032 596620 597088
rect 596676 597032 596744 597088
rect 596800 597032 596868 597088
rect 596924 597032 597020 597088
rect 596400 596964 597020 597032
rect 596400 596908 596496 596964
rect 596552 596908 596620 596964
rect 596676 596908 596744 596964
rect 596800 596908 596868 596964
rect 596924 596908 597020 596964
rect 596400 596840 597020 596908
rect 596400 596784 596496 596840
rect 596552 596784 596620 596840
rect 596676 596784 596744 596840
rect 596800 596784 596868 596840
rect 596924 596784 597020 596840
rect 596400 580350 597020 596784
rect 596400 580294 596496 580350
rect 596552 580294 596620 580350
rect 596676 580294 596744 580350
rect 596800 580294 596868 580350
rect 596924 580294 597020 580350
rect 596400 580226 597020 580294
rect 596400 580170 596496 580226
rect 596552 580170 596620 580226
rect 596676 580170 596744 580226
rect 596800 580170 596868 580226
rect 596924 580170 597020 580226
rect 596400 580102 597020 580170
rect 596400 580046 596496 580102
rect 596552 580046 596620 580102
rect 596676 580046 596744 580102
rect 596800 580046 596868 580102
rect 596924 580046 597020 580102
rect 596400 579978 597020 580046
rect 596400 579922 596496 579978
rect 596552 579922 596620 579978
rect 596676 579922 596744 579978
rect 596800 579922 596868 579978
rect 596924 579922 597020 579978
rect 596400 562350 597020 579922
rect 596400 562294 596496 562350
rect 596552 562294 596620 562350
rect 596676 562294 596744 562350
rect 596800 562294 596868 562350
rect 596924 562294 597020 562350
rect 596400 562226 597020 562294
rect 596400 562170 596496 562226
rect 596552 562170 596620 562226
rect 596676 562170 596744 562226
rect 596800 562170 596868 562226
rect 596924 562170 597020 562226
rect 596400 562102 597020 562170
rect 596400 562046 596496 562102
rect 596552 562046 596620 562102
rect 596676 562046 596744 562102
rect 596800 562046 596868 562102
rect 596924 562046 597020 562102
rect 596400 561978 597020 562046
rect 596400 561922 596496 561978
rect 596552 561922 596620 561978
rect 596676 561922 596744 561978
rect 596800 561922 596868 561978
rect 596924 561922 597020 561978
rect 596400 544350 597020 561922
rect 596400 544294 596496 544350
rect 596552 544294 596620 544350
rect 596676 544294 596744 544350
rect 596800 544294 596868 544350
rect 596924 544294 597020 544350
rect 596400 544226 597020 544294
rect 596400 544170 596496 544226
rect 596552 544170 596620 544226
rect 596676 544170 596744 544226
rect 596800 544170 596868 544226
rect 596924 544170 597020 544226
rect 596400 544102 597020 544170
rect 596400 544046 596496 544102
rect 596552 544046 596620 544102
rect 596676 544046 596744 544102
rect 596800 544046 596868 544102
rect 596924 544046 597020 544102
rect 596400 543978 597020 544046
rect 596400 543922 596496 543978
rect 596552 543922 596620 543978
rect 596676 543922 596744 543978
rect 596800 543922 596868 543978
rect 596924 543922 597020 543978
rect 596400 526350 597020 543922
rect 596400 526294 596496 526350
rect 596552 526294 596620 526350
rect 596676 526294 596744 526350
rect 596800 526294 596868 526350
rect 596924 526294 597020 526350
rect 596400 526226 597020 526294
rect 596400 526170 596496 526226
rect 596552 526170 596620 526226
rect 596676 526170 596744 526226
rect 596800 526170 596868 526226
rect 596924 526170 597020 526226
rect 596400 526102 597020 526170
rect 596400 526046 596496 526102
rect 596552 526046 596620 526102
rect 596676 526046 596744 526102
rect 596800 526046 596868 526102
rect 596924 526046 597020 526102
rect 596400 525978 597020 526046
rect 596400 525922 596496 525978
rect 596552 525922 596620 525978
rect 596676 525922 596744 525978
rect 596800 525922 596868 525978
rect 596924 525922 597020 525978
rect 596400 508350 597020 525922
rect 596400 508294 596496 508350
rect 596552 508294 596620 508350
rect 596676 508294 596744 508350
rect 596800 508294 596868 508350
rect 596924 508294 597020 508350
rect 596400 508226 597020 508294
rect 596400 508170 596496 508226
rect 596552 508170 596620 508226
rect 596676 508170 596744 508226
rect 596800 508170 596868 508226
rect 596924 508170 597020 508226
rect 596400 508102 597020 508170
rect 596400 508046 596496 508102
rect 596552 508046 596620 508102
rect 596676 508046 596744 508102
rect 596800 508046 596868 508102
rect 596924 508046 597020 508102
rect 596400 507978 597020 508046
rect 596400 507922 596496 507978
rect 596552 507922 596620 507978
rect 596676 507922 596744 507978
rect 596800 507922 596868 507978
rect 596924 507922 597020 507978
rect 596400 490350 597020 507922
rect 596400 490294 596496 490350
rect 596552 490294 596620 490350
rect 596676 490294 596744 490350
rect 596800 490294 596868 490350
rect 596924 490294 597020 490350
rect 596400 490226 597020 490294
rect 596400 490170 596496 490226
rect 596552 490170 596620 490226
rect 596676 490170 596744 490226
rect 596800 490170 596868 490226
rect 596924 490170 597020 490226
rect 596400 490102 597020 490170
rect 596400 490046 596496 490102
rect 596552 490046 596620 490102
rect 596676 490046 596744 490102
rect 596800 490046 596868 490102
rect 596924 490046 597020 490102
rect 596400 489978 597020 490046
rect 596400 489922 596496 489978
rect 596552 489922 596620 489978
rect 596676 489922 596744 489978
rect 596800 489922 596868 489978
rect 596924 489922 597020 489978
rect 596400 472350 597020 489922
rect 596400 472294 596496 472350
rect 596552 472294 596620 472350
rect 596676 472294 596744 472350
rect 596800 472294 596868 472350
rect 596924 472294 597020 472350
rect 596400 472226 597020 472294
rect 596400 472170 596496 472226
rect 596552 472170 596620 472226
rect 596676 472170 596744 472226
rect 596800 472170 596868 472226
rect 596924 472170 597020 472226
rect 596400 472102 597020 472170
rect 596400 472046 596496 472102
rect 596552 472046 596620 472102
rect 596676 472046 596744 472102
rect 596800 472046 596868 472102
rect 596924 472046 597020 472102
rect 596400 471978 597020 472046
rect 596400 471922 596496 471978
rect 596552 471922 596620 471978
rect 596676 471922 596744 471978
rect 596800 471922 596868 471978
rect 596924 471922 597020 471978
rect 596400 454350 597020 471922
rect 596400 454294 596496 454350
rect 596552 454294 596620 454350
rect 596676 454294 596744 454350
rect 596800 454294 596868 454350
rect 596924 454294 597020 454350
rect 596400 454226 597020 454294
rect 596400 454170 596496 454226
rect 596552 454170 596620 454226
rect 596676 454170 596744 454226
rect 596800 454170 596868 454226
rect 596924 454170 597020 454226
rect 596400 454102 597020 454170
rect 596400 454046 596496 454102
rect 596552 454046 596620 454102
rect 596676 454046 596744 454102
rect 596800 454046 596868 454102
rect 596924 454046 597020 454102
rect 596400 453978 597020 454046
rect 596400 453922 596496 453978
rect 596552 453922 596620 453978
rect 596676 453922 596744 453978
rect 596800 453922 596868 453978
rect 596924 453922 597020 453978
rect 596400 436350 597020 453922
rect 596400 436294 596496 436350
rect 596552 436294 596620 436350
rect 596676 436294 596744 436350
rect 596800 436294 596868 436350
rect 596924 436294 597020 436350
rect 596400 436226 597020 436294
rect 596400 436170 596496 436226
rect 596552 436170 596620 436226
rect 596676 436170 596744 436226
rect 596800 436170 596868 436226
rect 596924 436170 597020 436226
rect 596400 436102 597020 436170
rect 596400 436046 596496 436102
rect 596552 436046 596620 436102
rect 596676 436046 596744 436102
rect 596800 436046 596868 436102
rect 596924 436046 597020 436102
rect 596400 435978 597020 436046
rect 596400 435922 596496 435978
rect 596552 435922 596620 435978
rect 596676 435922 596744 435978
rect 596800 435922 596868 435978
rect 596924 435922 597020 435978
rect 596400 418350 597020 435922
rect 596400 418294 596496 418350
rect 596552 418294 596620 418350
rect 596676 418294 596744 418350
rect 596800 418294 596868 418350
rect 596924 418294 597020 418350
rect 596400 418226 597020 418294
rect 596400 418170 596496 418226
rect 596552 418170 596620 418226
rect 596676 418170 596744 418226
rect 596800 418170 596868 418226
rect 596924 418170 597020 418226
rect 596400 418102 597020 418170
rect 596400 418046 596496 418102
rect 596552 418046 596620 418102
rect 596676 418046 596744 418102
rect 596800 418046 596868 418102
rect 596924 418046 597020 418102
rect 596400 417978 597020 418046
rect 596400 417922 596496 417978
rect 596552 417922 596620 417978
rect 596676 417922 596744 417978
rect 596800 417922 596868 417978
rect 596924 417922 597020 417978
rect 596400 400350 597020 417922
rect 596400 400294 596496 400350
rect 596552 400294 596620 400350
rect 596676 400294 596744 400350
rect 596800 400294 596868 400350
rect 596924 400294 597020 400350
rect 596400 400226 597020 400294
rect 596400 400170 596496 400226
rect 596552 400170 596620 400226
rect 596676 400170 596744 400226
rect 596800 400170 596868 400226
rect 596924 400170 597020 400226
rect 596400 400102 597020 400170
rect 596400 400046 596496 400102
rect 596552 400046 596620 400102
rect 596676 400046 596744 400102
rect 596800 400046 596868 400102
rect 596924 400046 597020 400102
rect 596400 399978 597020 400046
rect 596400 399922 596496 399978
rect 596552 399922 596620 399978
rect 596676 399922 596744 399978
rect 596800 399922 596868 399978
rect 596924 399922 597020 399978
rect 596400 382350 597020 399922
rect 596400 382294 596496 382350
rect 596552 382294 596620 382350
rect 596676 382294 596744 382350
rect 596800 382294 596868 382350
rect 596924 382294 597020 382350
rect 596400 382226 597020 382294
rect 596400 382170 596496 382226
rect 596552 382170 596620 382226
rect 596676 382170 596744 382226
rect 596800 382170 596868 382226
rect 596924 382170 597020 382226
rect 596400 382102 597020 382170
rect 596400 382046 596496 382102
rect 596552 382046 596620 382102
rect 596676 382046 596744 382102
rect 596800 382046 596868 382102
rect 596924 382046 597020 382102
rect 596400 381978 597020 382046
rect 596400 381922 596496 381978
rect 596552 381922 596620 381978
rect 596676 381922 596744 381978
rect 596800 381922 596868 381978
rect 596924 381922 597020 381978
rect 596400 364350 597020 381922
rect 596400 364294 596496 364350
rect 596552 364294 596620 364350
rect 596676 364294 596744 364350
rect 596800 364294 596868 364350
rect 596924 364294 597020 364350
rect 596400 364226 597020 364294
rect 596400 364170 596496 364226
rect 596552 364170 596620 364226
rect 596676 364170 596744 364226
rect 596800 364170 596868 364226
rect 596924 364170 597020 364226
rect 596400 364102 597020 364170
rect 596400 364046 596496 364102
rect 596552 364046 596620 364102
rect 596676 364046 596744 364102
rect 596800 364046 596868 364102
rect 596924 364046 597020 364102
rect 596400 363978 597020 364046
rect 596400 363922 596496 363978
rect 596552 363922 596620 363978
rect 596676 363922 596744 363978
rect 596800 363922 596868 363978
rect 596924 363922 597020 363978
rect 596400 346350 597020 363922
rect 596400 346294 596496 346350
rect 596552 346294 596620 346350
rect 596676 346294 596744 346350
rect 596800 346294 596868 346350
rect 596924 346294 597020 346350
rect 596400 346226 597020 346294
rect 596400 346170 596496 346226
rect 596552 346170 596620 346226
rect 596676 346170 596744 346226
rect 596800 346170 596868 346226
rect 596924 346170 597020 346226
rect 596400 346102 597020 346170
rect 596400 346046 596496 346102
rect 596552 346046 596620 346102
rect 596676 346046 596744 346102
rect 596800 346046 596868 346102
rect 596924 346046 597020 346102
rect 596400 345978 597020 346046
rect 596400 345922 596496 345978
rect 596552 345922 596620 345978
rect 596676 345922 596744 345978
rect 596800 345922 596868 345978
rect 596924 345922 597020 345978
rect 596400 328350 597020 345922
rect 596400 328294 596496 328350
rect 596552 328294 596620 328350
rect 596676 328294 596744 328350
rect 596800 328294 596868 328350
rect 596924 328294 597020 328350
rect 596400 328226 597020 328294
rect 596400 328170 596496 328226
rect 596552 328170 596620 328226
rect 596676 328170 596744 328226
rect 596800 328170 596868 328226
rect 596924 328170 597020 328226
rect 596400 328102 597020 328170
rect 596400 328046 596496 328102
rect 596552 328046 596620 328102
rect 596676 328046 596744 328102
rect 596800 328046 596868 328102
rect 596924 328046 597020 328102
rect 596400 327978 597020 328046
rect 596400 327922 596496 327978
rect 596552 327922 596620 327978
rect 596676 327922 596744 327978
rect 596800 327922 596868 327978
rect 596924 327922 597020 327978
rect 596400 310350 597020 327922
rect 596400 310294 596496 310350
rect 596552 310294 596620 310350
rect 596676 310294 596744 310350
rect 596800 310294 596868 310350
rect 596924 310294 597020 310350
rect 596400 310226 597020 310294
rect 596400 310170 596496 310226
rect 596552 310170 596620 310226
rect 596676 310170 596744 310226
rect 596800 310170 596868 310226
rect 596924 310170 597020 310226
rect 596400 310102 597020 310170
rect 596400 310046 596496 310102
rect 596552 310046 596620 310102
rect 596676 310046 596744 310102
rect 596800 310046 596868 310102
rect 596924 310046 597020 310102
rect 596400 309978 597020 310046
rect 596400 309922 596496 309978
rect 596552 309922 596620 309978
rect 596676 309922 596744 309978
rect 596800 309922 596868 309978
rect 596924 309922 597020 309978
rect 596400 292350 597020 309922
rect 596400 292294 596496 292350
rect 596552 292294 596620 292350
rect 596676 292294 596744 292350
rect 596800 292294 596868 292350
rect 596924 292294 597020 292350
rect 596400 292226 597020 292294
rect 596400 292170 596496 292226
rect 596552 292170 596620 292226
rect 596676 292170 596744 292226
rect 596800 292170 596868 292226
rect 596924 292170 597020 292226
rect 596400 292102 597020 292170
rect 596400 292046 596496 292102
rect 596552 292046 596620 292102
rect 596676 292046 596744 292102
rect 596800 292046 596868 292102
rect 596924 292046 597020 292102
rect 596400 291978 597020 292046
rect 596400 291922 596496 291978
rect 596552 291922 596620 291978
rect 596676 291922 596744 291978
rect 596800 291922 596868 291978
rect 596924 291922 597020 291978
rect 596400 274350 597020 291922
rect 596400 274294 596496 274350
rect 596552 274294 596620 274350
rect 596676 274294 596744 274350
rect 596800 274294 596868 274350
rect 596924 274294 597020 274350
rect 596400 274226 597020 274294
rect 596400 274170 596496 274226
rect 596552 274170 596620 274226
rect 596676 274170 596744 274226
rect 596800 274170 596868 274226
rect 596924 274170 597020 274226
rect 596400 274102 597020 274170
rect 596400 274046 596496 274102
rect 596552 274046 596620 274102
rect 596676 274046 596744 274102
rect 596800 274046 596868 274102
rect 596924 274046 597020 274102
rect 596400 273978 597020 274046
rect 596400 273922 596496 273978
rect 596552 273922 596620 273978
rect 596676 273922 596744 273978
rect 596800 273922 596868 273978
rect 596924 273922 597020 273978
rect 596400 256350 597020 273922
rect 596400 256294 596496 256350
rect 596552 256294 596620 256350
rect 596676 256294 596744 256350
rect 596800 256294 596868 256350
rect 596924 256294 597020 256350
rect 596400 256226 597020 256294
rect 596400 256170 596496 256226
rect 596552 256170 596620 256226
rect 596676 256170 596744 256226
rect 596800 256170 596868 256226
rect 596924 256170 597020 256226
rect 596400 256102 597020 256170
rect 596400 256046 596496 256102
rect 596552 256046 596620 256102
rect 596676 256046 596744 256102
rect 596800 256046 596868 256102
rect 596924 256046 597020 256102
rect 596400 255978 597020 256046
rect 596400 255922 596496 255978
rect 596552 255922 596620 255978
rect 596676 255922 596744 255978
rect 596800 255922 596868 255978
rect 596924 255922 597020 255978
rect 596400 238350 597020 255922
rect 596400 238294 596496 238350
rect 596552 238294 596620 238350
rect 596676 238294 596744 238350
rect 596800 238294 596868 238350
rect 596924 238294 597020 238350
rect 596400 238226 597020 238294
rect 596400 238170 596496 238226
rect 596552 238170 596620 238226
rect 596676 238170 596744 238226
rect 596800 238170 596868 238226
rect 596924 238170 597020 238226
rect 596400 238102 597020 238170
rect 596400 238046 596496 238102
rect 596552 238046 596620 238102
rect 596676 238046 596744 238102
rect 596800 238046 596868 238102
rect 596924 238046 597020 238102
rect 596400 237978 597020 238046
rect 596400 237922 596496 237978
rect 596552 237922 596620 237978
rect 596676 237922 596744 237978
rect 596800 237922 596868 237978
rect 596924 237922 597020 237978
rect 596400 220350 597020 237922
rect 596400 220294 596496 220350
rect 596552 220294 596620 220350
rect 596676 220294 596744 220350
rect 596800 220294 596868 220350
rect 596924 220294 597020 220350
rect 596400 220226 597020 220294
rect 596400 220170 596496 220226
rect 596552 220170 596620 220226
rect 596676 220170 596744 220226
rect 596800 220170 596868 220226
rect 596924 220170 597020 220226
rect 596400 220102 597020 220170
rect 596400 220046 596496 220102
rect 596552 220046 596620 220102
rect 596676 220046 596744 220102
rect 596800 220046 596868 220102
rect 596924 220046 597020 220102
rect 596400 219978 597020 220046
rect 596400 219922 596496 219978
rect 596552 219922 596620 219978
rect 596676 219922 596744 219978
rect 596800 219922 596868 219978
rect 596924 219922 597020 219978
rect 596400 202350 597020 219922
rect 596400 202294 596496 202350
rect 596552 202294 596620 202350
rect 596676 202294 596744 202350
rect 596800 202294 596868 202350
rect 596924 202294 597020 202350
rect 596400 202226 597020 202294
rect 596400 202170 596496 202226
rect 596552 202170 596620 202226
rect 596676 202170 596744 202226
rect 596800 202170 596868 202226
rect 596924 202170 597020 202226
rect 596400 202102 597020 202170
rect 596400 202046 596496 202102
rect 596552 202046 596620 202102
rect 596676 202046 596744 202102
rect 596800 202046 596868 202102
rect 596924 202046 597020 202102
rect 596400 201978 597020 202046
rect 596400 201922 596496 201978
rect 596552 201922 596620 201978
rect 596676 201922 596744 201978
rect 596800 201922 596868 201978
rect 596924 201922 597020 201978
rect 596400 184350 597020 201922
rect 596400 184294 596496 184350
rect 596552 184294 596620 184350
rect 596676 184294 596744 184350
rect 596800 184294 596868 184350
rect 596924 184294 597020 184350
rect 596400 184226 597020 184294
rect 596400 184170 596496 184226
rect 596552 184170 596620 184226
rect 596676 184170 596744 184226
rect 596800 184170 596868 184226
rect 596924 184170 597020 184226
rect 596400 184102 597020 184170
rect 596400 184046 596496 184102
rect 596552 184046 596620 184102
rect 596676 184046 596744 184102
rect 596800 184046 596868 184102
rect 596924 184046 597020 184102
rect 596400 183978 597020 184046
rect 596400 183922 596496 183978
rect 596552 183922 596620 183978
rect 596676 183922 596744 183978
rect 596800 183922 596868 183978
rect 596924 183922 597020 183978
rect 596400 166350 597020 183922
rect 596400 166294 596496 166350
rect 596552 166294 596620 166350
rect 596676 166294 596744 166350
rect 596800 166294 596868 166350
rect 596924 166294 597020 166350
rect 596400 166226 597020 166294
rect 596400 166170 596496 166226
rect 596552 166170 596620 166226
rect 596676 166170 596744 166226
rect 596800 166170 596868 166226
rect 596924 166170 597020 166226
rect 596400 166102 597020 166170
rect 596400 166046 596496 166102
rect 596552 166046 596620 166102
rect 596676 166046 596744 166102
rect 596800 166046 596868 166102
rect 596924 166046 597020 166102
rect 596400 165978 597020 166046
rect 596400 165922 596496 165978
rect 596552 165922 596620 165978
rect 596676 165922 596744 165978
rect 596800 165922 596868 165978
rect 596924 165922 597020 165978
rect 596400 148350 597020 165922
rect 596400 148294 596496 148350
rect 596552 148294 596620 148350
rect 596676 148294 596744 148350
rect 596800 148294 596868 148350
rect 596924 148294 597020 148350
rect 596400 148226 597020 148294
rect 596400 148170 596496 148226
rect 596552 148170 596620 148226
rect 596676 148170 596744 148226
rect 596800 148170 596868 148226
rect 596924 148170 597020 148226
rect 596400 148102 597020 148170
rect 596400 148046 596496 148102
rect 596552 148046 596620 148102
rect 596676 148046 596744 148102
rect 596800 148046 596868 148102
rect 596924 148046 597020 148102
rect 596400 147978 597020 148046
rect 596400 147922 596496 147978
rect 596552 147922 596620 147978
rect 596676 147922 596744 147978
rect 596800 147922 596868 147978
rect 596924 147922 597020 147978
rect 596400 130350 597020 147922
rect 596400 130294 596496 130350
rect 596552 130294 596620 130350
rect 596676 130294 596744 130350
rect 596800 130294 596868 130350
rect 596924 130294 597020 130350
rect 596400 130226 597020 130294
rect 596400 130170 596496 130226
rect 596552 130170 596620 130226
rect 596676 130170 596744 130226
rect 596800 130170 596868 130226
rect 596924 130170 597020 130226
rect 596400 130102 597020 130170
rect 596400 130046 596496 130102
rect 596552 130046 596620 130102
rect 596676 130046 596744 130102
rect 596800 130046 596868 130102
rect 596924 130046 597020 130102
rect 596400 129978 597020 130046
rect 596400 129922 596496 129978
rect 596552 129922 596620 129978
rect 596676 129922 596744 129978
rect 596800 129922 596868 129978
rect 596924 129922 597020 129978
rect 596400 112350 597020 129922
rect 596400 112294 596496 112350
rect 596552 112294 596620 112350
rect 596676 112294 596744 112350
rect 596800 112294 596868 112350
rect 596924 112294 597020 112350
rect 596400 112226 597020 112294
rect 596400 112170 596496 112226
rect 596552 112170 596620 112226
rect 596676 112170 596744 112226
rect 596800 112170 596868 112226
rect 596924 112170 597020 112226
rect 596400 112102 597020 112170
rect 596400 112046 596496 112102
rect 596552 112046 596620 112102
rect 596676 112046 596744 112102
rect 596800 112046 596868 112102
rect 596924 112046 597020 112102
rect 596400 111978 597020 112046
rect 596400 111922 596496 111978
rect 596552 111922 596620 111978
rect 596676 111922 596744 111978
rect 596800 111922 596868 111978
rect 596924 111922 597020 111978
rect 596400 94350 597020 111922
rect 596400 94294 596496 94350
rect 596552 94294 596620 94350
rect 596676 94294 596744 94350
rect 596800 94294 596868 94350
rect 596924 94294 597020 94350
rect 596400 94226 597020 94294
rect 596400 94170 596496 94226
rect 596552 94170 596620 94226
rect 596676 94170 596744 94226
rect 596800 94170 596868 94226
rect 596924 94170 597020 94226
rect 596400 94102 597020 94170
rect 596400 94046 596496 94102
rect 596552 94046 596620 94102
rect 596676 94046 596744 94102
rect 596800 94046 596868 94102
rect 596924 94046 597020 94102
rect 596400 93978 597020 94046
rect 596400 93922 596496 93978
rect 596552 93922 596620 93978
rect 596676 93922 596744 93978
rect 596800 93922 596868 93978
rect 596924 93922 597020 93978
rect 596400 76350 597020 93922
rect 596400 76294 596496 76350
rect 596552 76294 596620 76350
rect 596676 76294 596744 76350
rect 596800 76294 596868 76350
rect 596924 76294 597020 76350
rect 596400 76226 597020 76294
rect 596400 76170 596496 76226
rect 596552 76170 596620 76226
rect 596676 76170 596744 76226
rect 596800 76170 596868 76226
rect 596924 76170 597020 76226
rect 596400 76102 597020 76170
rect 596400 76046 596496 76102
rect 596552 76046 596620 76102
rect 596676 76046 596744 76102
rect 596800 76046 596868 76102
rect 596924 76046 597020 76102
rect 596400 75978 597020 76046
rect 596400 75922 596496 75978
rect 596552 75922 596620 75978
rect 596676 75922 596744 75978
rect 596800 75922 596868 75978
rect 596924 75922 597020 75978
rect 596400 58350 597020 75922
rect 596400 58294 596496 58350
rect 596552 58294 596620 58350
rect 596676 58294 596744 58350
rect 596800 58294 596868 58350
rect 596924 58294 597020 58350
rect 596400 58226 597020 58294
rect 596400 58170 596496 58226
rect 596552 58170 596620 58226
rect 596676 58170 596744 58226
rect 596800 58170 596868 58226
rect 596924 58170 597020 58226
rect 596400 58102 597020 58170
rect 596400 58046 596496 58102
rect 596552 58046 596620 58102
rect 596676 58046 596744 58102
rect 596800 58046 596868 58102
rect 596924 58046 597020 58102
rect 596400 57978 597020 58046
rect 596400 57922 596496 57978
rect 596552 57922 596620 57978
rect 596676 57922 596744 57978
rect 596800 57922 596868 57978
rect 596924 57922 597020 57978
rect 596400 40350 597020 57922
rect 596400 40294 596496 40350
rect 596552 40294 596620 40350
rect 596676 40294 596744 40350
rect 596800 40294 596868 40350
rect 596924 40294 597020 40350
rect 596400 40226 597020 40294
rect 596400 40170 596496 40226
rect 596552 40170 596620 40226
rect 596676 40170 596744 40226
rect 596800 40170 596868 40226
rect 596924 40170 597020 40226
rect 596400 40102 597020 40170
rect 596400 40046 596496 40102
rect 596552 40046 596620 40102
rect 596676 40046 596744 40102
rect 596800 40046 596868 40102
rect 596924 40046 597020 40102
rect 596400 39978 597020 40046
rect 596400 39922 596496 39978
rect 596552 39922 596620 39978
rect 596676 39922 596744 39978
rect 596800 39922 596868 39978
rect 596924 39922 597020 39978
rect 596400 22350 597020 39922
rect 596400 22294 596496 22350
rect 596552 22294 596620 22350
rect 596676 22294 596744 22350
rect 596800 22294 596868 22350
rect 596924 22294 597020 22350
rect 596400 22226 597020 22294
rect 596400 22170 596496 22226
rect 596552 22170 596620 22226
rect 596676 22170 596744 22226
rect 596800 22170 596868 22226
rect 596924 22170 597020 22226
rect 596400 22102 597020 22170
rect 596400 22046 596496 22102
rect 596552 22046 596620 22102
rect 596676 22046 596744 22102
rect 596800 22046 596868 22102
rect 596924 22046 597020 22102
rect 596400 21978 597020 22046
rect 596400 21922 596496 21978
rect 596552 21922 596620 21978
rect 596676 21922 596744 21978
rect 596800 21922 596868 21978
rect 596924 21922 597020 21978
rect 596400 4350 597020 21922
rect 596400 4294 596496 4350
rect 596552 4294 596620 4350
rect 596676 4294 596744 4350
rect 596800 4294 596868 4350
rect 596924 4294 597020 4350
rect 596400 4226 597020 4294
rect 596400 4170 596496 4226
rect 596552 4170 596620 4226
rect 596676 4170 596744 4226
rect 596800 4170 596868 4226
rect 596924 4170 597020 4226
rect 596400 4102 597020 4170
rect 596400 4046 596496 4102
rect 596552 4046 596620 4102
rect 596676 4046 596744 4102
rect 596800 4046 596868 4102
rect 596924 4046 597020 4102
rect 596400 3978 597020 4046
rect 596400 3922 596496 3978
rect 596552 3922 596620 3978
rect 596676 3922 596744 3978
rect 596800 3922 596868 3978
rect 596924 3922 597020 3978
rect 596400 -160 597020 3922
rect 596400 -216 596496 -160
rect 596552 -216 596620 -160
rect 596676 -216 596744 -160
rect 596800 -216 596868 -160
rect 596924 -216 597020 -160
rect 596400 -284 597020 -216
rect 596400 -340 596496 -284
rect 596552 -340 596620 -284
rect 596676 -340 596744 -284
rect 596800 -340 596868 -284
rect 596924 -340 597020 -284
rect 596400 -408 597020 -340
rect 596400 -464 596496 -408
rect 596552 -464 596620 -408
rect 596676 -464 596744 -408
rect 596800 -464 596868 -408
rect 596924 -464 597020 -408
rect 596400 -532 597020 -464
rect 596400 -588 596496 -532
rect 596552 -588 596620 -532
rect 596676 -588 596744 -532
rect 596800 -588 596868 -532
rect 596924 -588 597020 -532
rect 596400 -684 597020 -588
rect 597360 586350 597980 597744
rect 597360 586294 597456 586350
rect 597512 586294 597580 586350
rect 597636 586294 597704 586350
rect 597760 586294 597828 586350
rect 597884 586294 597980 586350
rect 597360 586226 597980 586294
rect 597360 586170 597456 586226
rect 597512 586170 597580 586226
rect 597636 586170 597704 586226
rect 597760 586170 597828 586226
rect 597884 586170 597980 586226
rect 597360 586102 597980 586170
rect 597360 586046 597456 586102
rect 597512 586046 597580 586102
rect 597636 586046 597704 586102
rect 597760 586046 597828 586102
rect 597884 586046 597980 586102
rect 597360 585978 597980 586046
rect 597360 585922 597456 585978
rect 597512 585922 597580 585978
rect 597636 585922 597704 585978
rect 597760 585922 597828 585978
rect 597884 585922 597980 585978
rect 597360 568350 597980 585922
rect 597360 568294 597456 568350
rect 597512 568294 597580 568350
rect 597636 568294 597704 568350
rect 597760 568294 597828 568350
rect 597884 568294 597980 568350
rect 597360 568226 597980 568294
rect 597360 568170 597456 568226
rect 597512 568170 597580 568226
rect 597636 568170 597704 568226
rect 597760 568170 597828 568226
rect 597884 568170 597980 568226
rect 597360 568102 597980 568170
rect 597360 568046 597456 568102
rect 597512 568046 597580 568102
rect 597636 568046 597704 568102
rect 597760 568046 597828 568102
rect 597884 568046 597980 568102
rect 597360 567978 597980 568046
rect 597360 567922 597456 567978
rect 597512 567922 597580 567978
rect 597636 567922 597704 567978
rect 597760 567922 597828 567978
rect 597884 567922 597980 567978
rect 597360 550350 597980 567922
rect 597360 550294 597456 550350
rect 597512 550294 597580 550350
rect 597636 550294 597704 550350
rect 597760 550294 597828 550350
rect 597884 550294 597980 550350
rect 597360 550226 597980 550294
rect 597360 550170 597456 550226
rect 597512 550170 597580 550226
rect 597636 550170 597704 550226
rect 597760 550170 597828 550226
rect 597884 550170 597980 550226
rect 597360 550102 597980 550170
rect 597360 550046 597456 550102
rect 597512 550046 597580 550102
rect 597636 550046 597704 550102
rect 597760 550046 597828 550102
rect 597884 550046 597980 550102
rect 597360 549978 597980 550046
rect 597360 549922 597456 549978
rect 597512 549922 597580 549978
rect 597636 549922 597704 549978
rect 597760 549922 597828 549978
rect 597884 549922 597980 549978
rect 597360 532350 597980 549922
rect 597360 532294 597456 532350
rect 597512 532294 597580 532350
rect 597636 532294 597704 532350
rect 597760 532294 597828 532350
rect 597884 532294 597980 532350
rect 597360 532226 597980 532294
rect 597360 532170 597456 532226
rect 597512 532170 597580 532226
rect 597636 532170 597704 532226
rect 597760 532170 597828 532226
rect 597884 532170 597980 532226
rect 597360 532102 597980 532170
rect 597360 532046 597456 532102
rect 597512 532046 597580 532102
rect 597636 532046 597704 532102
rect 597760 532046 597828 532102
rect 597884 532046 597980 532102
rect 597360 531978 597980 532046
rect 597360 531922 597456 531978
rect 597512 531922 597580 531978
rect 597636 531922 597704 531978
rect 597760 531922 597828 531978
rect 597884 531922 597980 531978
rect 597360 514350 597980 531922
rect 597360 514294 597456 514350
rect 597512 514294 597580 514350
rect 597636 514294 597704 514350
rect 597760 514294 597828 514350
rect 597884 514294 597980 514350
rect 597360 514226 597980 514294
rect 597360 514170 597456 514226
rect 597512 514170 597580 514226
rect 597636 514170 597704 514226
rect 597760 514170 597828 514226
rect 597884 514170 597980 514226
rect 597360 514102 597980 514170
rect 597360 514046 597456 514102
rect 597512 514046 597580 514102
rect 597636 514046 597704 514102
rect 597760 514046 597828 514102
rect 597884 514046 597980 514102
rect 597360 513978 597980 514046
rect 597360 513922 597456 513978
rect 597512 513922 597580 513978
rect 597636 513922 597704 513978
rect 597760 513922 597828 513978
rect 597884 513922 597980 513978
rect 597360 496350 597980 513922
rect 597360 496294 597456 496350
rect 597512 496294 597580 496350
rect 597636 496294 597704 496350
rect 597760 496294 597828 496350
rect 597884 496294 597980 496350
rect 597360 496226 597980 496294
rect 597360 496170 597456 496226
rect 597512 496170 597580 496226
rect 597636 496170 597704 496226
rect 597760 496170 597828 496226
rect 597884 496170 597980 496226
rect 597360 496102 597980 496170
rect 597360 496046 597456 496102
rect 597512 496046 597580 496102
rect 597636 496046 597704 496102
rect 597760 496046 597828 496102
rect 597884 496046 597980 496102
rect 597360 495978 597980 496046
rect 597360 495922 597456 495978
rect 597512 495922 597580 495978
rect 597636 495922 597704 495978
rect 597760 495922 597828 495978
rect 597884 495922 597980 495978
rect 597360 478350 597980 495922
rect 597360 478294 597456 478350
rect 597512 478294 597580 478350
rect 597636 478294 597704 478350
rect 597760 478294 597828 478350
rect 597884 478294 597980 478350
rect 597360 478226 597980 478294
rect 597360 478170 597456 478226
rect 597512 478170 597580 478226
rect 597636 478170 597704 478226
rect 597760 478170 597828 478226
rect 597884 478170 597980 478226
rect 597360 478102 597980 478170
rect 597360 478046 597456 478102
rect 597512 478046 597580 478102
rect 597636 478046 597704 478102
rect 597760 478046 597828 478102
rect 597884 478046 597980 478102
rect 597360 477978 597980 478046
rect 597360 477922 597456 477978
rect 597512 477922 597580 477978
rect 597636 477922 597704 477978
rect 597760 477922 597828 477978
rect 597884 477922 597980 477978
rect 597360 460350 597980 477922
rect 597360 460294 597456 460350
rect 597512 460294 597580 460350
rect 597636 460294 597704 460350
rect 597760 460294 597828 460350
rect 597884 460294 597980 460350
rect 597360 460226 597980 460294
rect 597360 460170 597456 460226
rect 597512 460170 597580 460226
rect 597636 460170 597704 460226
rect 597760 460170 597828 460226
rect 597884 460170 597980 460226
rect 597360 460102 597980 460170
rect 597360 460046 597456 460102
rect 597512 460046 597580 460102
rect 597636 460046 597704 460102
rect 597760 460046 597828 460102
rect 597884 460046 597980 460102
rect 597360 459978 597980 460046
rect 597360 459922 597456 459978
rect 597512 459922 597580 459978
rect 597636 459922 597704 459978
rect 597760 459922 597828 459978
rect 597884 459922 597980 459978
rect 597360 442350 597980 459922
rect 597360 442294 597456 442350
rect 597512 442294 597580 442350
rect 597636 442294 597704 442350
rect 597760 442294 597828 442350
rect 597884 442294 597980 442350
rect 597360 442226 597980 442294
rect 597360 442170 597456 442226
rect 597512 442170 597580 442226
rect 597636 442170 597704 442226
rect 597760 442170 597828 442226
rect 597884 442170 597980 442226
rect 597360 442102 597980 442170
rect 597360 442046 597456 442102
rect 597512 442046 597580 442102
rect 597636 442046 597704 442102
rect 597760 442046 597828 442102
rect 597884 442046 597980 442102
rect 597360 441978 597980 442046
rect 597360 441922 597456 441978
rect 597512 441922 597580 441978
rect 597636 441922 597704 441978
rect 597760 441922 597828 441978
rect 597884 441922 597980 441978
rect 597360 424350 597980 441922
rect 597360 424294 597456 424350
rect 597512 424294 597580 424350
rect 597636 424294 597704 424350
rect 597760 424294 597828 424350
rect 597884 424294 597980 424350
rect 597360 424226 597980 424294
rect 597360 424170 597456 424226
rect 597512 424170 597580 424226
rect 597636 424170 597704 424226
rect 597760 424170 597828 424226
rect 597884 424170 597980 424226
rect 597360 424102 597980 424170
rect 597360 424046 597456 424102
rect 597512 424046 597580 424102
rect 597636 424046 597704 424102
rect 597760 424046 597828 424102
rect 597884 424046 597980 424102
rect 597360 423978 597980 424046
rect 597360 423922 597456 423978
rect 597512 423922 597580 423978
rect 597636 423922 597704 423978
rect 597760 423922 597828 423978
rect 597884 423922 597980 423978
rect 597360 406350 597980 423922
rect 597360 406294 597456 406350
rect 597512 406294 597580 406350
rect 597636 406294 597704 406350
rect 597760 406294 597828 406350
rect 597884 406294 597980 406350
rect 597360 406226 597980 406294
rect 597360 406170 597456 406226
rect 597512 406170 597580 406226
rect 597636 406170 597704 406226
rect 597760 406170 597828 406226
rect 597884 406170 597980 406226
rect 597360 406102 597980 406170
rect 597360 406046 597456 406102
rect 597512 406046 597580 406102
rect 597636 406046 597704 406102
rect 597760 406046 597828 406102
rect 597884 406046 597980 406102
rect 597360 405978 597980 406046
rect 597360 405922 597456 405978
rect 597512 405922 597580 405978
rect 597636 405922 597704 405978
rect 597760 405922 597828 405978
rect 597884 405922 597980 405978
rect 597360 388350 597980 405922
rect 597360 388294 597456 388350
rect 597512 388294 597580 388350
rect 597636 388294 597704 388350
rect 597760 388294 597828 388350
rect 597884 388294 597980 388350
rect 597360 388226 597980 388294
rect 597360 388170 597456 388226
rect 597512 388170 597580 388226
rect 597636 388170 597704 388226
rect 597760 388170 597828 388226
rect 597884 388170 597980 388226
rect 597360 388102 597980 388170
rect 597360 388046 597456 388102
rect 597512 388046 597580 388102
rect 597636 388046 597704 388102
rect 597760 388046 597828 388102
rect 597884 388046 597980 388102
rect 597360 387978 597980 388046
rect 597360 387922 597456 387978
rect 597512 387922 597580 387978
rect 597636 387922 597704 387978
rect 597760 387922 597828 387978
rect 597884 387922 597980 387978
rect 597360 370350 597980 387922
rect 597360 370294 597456 370350
rect 597512 370294 597580 370350
rect 597636 370294 597704 370350
rect 597760 370294 597828 370350
rect 597884 370294 597980 370350
rect 597360 370226 597980 370294
rect 597360 370170 597456 370226
rect 597512 370170 597580 370226
rect 597636 370170 597704 370226
rect 597760 370170 597828 370226
rect 597884 370170 597980 370226
rect 597360 370102 597980 370170
rect 597360 370046 597456 370102
rect 597512 370046 597580 370102
rect 597636 370046 597704 370102
rect 597760 370046 597828 370102
rect 597884 370046 597980 370102
rect 597360 369978 597980 370046
rect 597360 369922 597456 369978
rect 597512 369922 597580 369978
rect 597636 369922 597704 369978
rect 597760 369922 597828 369978
rect 597884 369922 597980 369978
rect 597360 352350 597980 369922
rect 597360 352294 597456 352350
rect 597512 352294 597580 352350
rect 597636 352294 597704 352350
rect 597760 352294 597828 352350
rect 597884 352294 597980 352350
rect 597360 352226 597980 352294
rect 597360 352170 597456 352226
rect 597512 352170 597580 352226
rect 597636 352170 597704 352226
rect 597760 352170 597828 352226
rect 597884 352170 597980 352226
rect 597360 352102 597980 352170
rect 597360 352046 597456 352102
rect 597512 352046 597580 352102
rect 597636 352046 597704 352102
rect 597760 352046 597828 352102
rect 597884 352046 597980 352102
rect 597360 351978 597980 352046
rect 597360 351922 597456 351978
rect 597512 351922 597580 351978
rect 597636 351922 597704 351978
rect 597760 351922 597828 351978
rect 597884 351922 597980 351978
rect 597360 334350 597980 351922
rect 597360 334294 597456 334350
rect 597512 334294 597580 334350
rect 597636 334294 597704 334350
rect 597760 334294 597828 334350
rect 597884 334294 597980 334350
rect 597360 334226 597980 334294
rect 597360 334170 597456 334226
rect 597512 334170 597580 334226
rect 597636 334170 597704 334226
rect 597760 334170 597828 334226
rect 597884 334170 597980 334226
rect 597360 334102 597980 334170
rect 597360 334046 597456 334102
rect 597512 334046 597580 334102
rect 597636 334046 597704 334102
rect 597760 334046 597828 334102
rect 597884 334046 597980 334102
rect 597360 333978 597980 334046
rect 597360 333922 597456 333978
rect 597512 333922 597580 333978
rect 597636 333922 597704 333978
rect 597760 333922 597828 333978
rect 597884 333922 597980 333978
rect 597360 316350 597980 333922
rect 597360 316294 597456 316350
rect 597512 316294 597580 316350
rect 597636 316294 597704 316350
rect 597760 316294 597828 316350
rect 597884 316294 597980 316350
rect 597360 316226 597980 316294
rect 597360 316170 597456 316226
rect 597512 316170 597580 316226
rect 597636 316170 597704 316226
rect 597760 316170 597828 316226
rect 597884 316170 597980 316226
rect 597360 316102 597980 316170
rect 597360 316046 597456 316102
rect 597512 316046 597580 316102
rect 597636 316046 597704 316102
rect 597760 316046 597828 316102
rect 597884 316046 597980 316102
rect 597360 315978 597980 316046
rect 597360 315922 597456 315978
rect 597512 315922 597580 315978
rect 597636 315922 597704 315978
rect 597760 315922 597828 315978
rect 597884 315922 597980 315978
rect 597360 298350 597980 315922
rect 597360 298294 597456 298350
rect 597512 298294 597580 298350
rect 597636 298294 597704 298350
rect 597760 298294 597828 298350
rect 597884 298294 597980 298350
rect 597360 298226 597980 298294
rect 597360 298170 597456 298226
rect 597512 298170 597580 298226
rect 597636 298170 597704 298226
rect 597760 298170 597828 298226
rect 597884 298170 597980 298226
rect 597360 298102 597980 298170
rect 597360 298046 597456 298102
rect 597512 298046 597580 298102
rect 597636 298046 597704 298102
rect 597760 298046 597828 298102
rect 597884 298046 597980 298102
rect 597360 297978 597980 298046
rect 597360 297922 597456 297978
rect 597512 297922 597580 297978
rect 597636 297922 597704 297978
rect 597760 297922 597828 297978
rect 597884 297922 597980 297978
rect 597360 280350 597980 297922
rect 597360 280294 597456 280350
rect 597512 280294 597580 280350
rect 597636 280294 597704 280350
rect 597760 280294 597828 280350
rect 597884 280294 597980 280350
rect 597360 280226 597980 280294
rect 597360 280170 597456 280226
rect 597512 280170 597580 280226
rect 597636 280170 597704 280226
rect 597760 280170 597828 280226
rect 597884 280170 597980 280226
rect 597360 280102 597980 280170
rect 597360 280046 597456 280102
rect 597512 280046 597580 280102
rect 597636 280046 597704 280102
rect 597760 280046 597828 280102
rect 597884 280046 597980 280102
rect 597360 279978 597980 280046
rect 597360 279922 597456 279978
rect 597512 279922 597580 279978
rect 597636 279922 597704 279978
rect 597760 279922 597828 279978
rect 597884 279922 597980 279978
rect 597360 262350 597980 279922
rect 597360 262294 597456 262350
rect 597512 262294 597580 262350
rect 597636 262294 597704 262350
rect 597760 262294 597828 262350
rect 597884 262294 597980 262350
rect 597360 262226 597980 262294
rect 597360 262170 597456 262226
rect 597512 262170 597580 262226
rect 597636 262170 597704 262226
rect 597760 262170 597828 262226
rect 597884 262170 597980 262226
rect 597360 262102 597980 262170
rect 597360 262046 597456 262102
rect 597512 262046 597580 262102
rect 597636 262046 597704 262102
rect 597760 262046 597828 262102
rect 597884 262046 597980 262102
rect 597360 261978 597980 262046
rect 597360 261922 597456 261978
rect 597512 261922 597580 261978
rect 597636 261922 597704 261978
rect 597760 261922 597828 261978
rect 597884 261922 597980 261978
rect 597360 244350 597980 261922
rect 597360 244294 597456 244350
rect 597512 244294 597580 244350
rect 597636 244294 597704 244350
rect 597760 244294 597828 244350
rect 597884 244294 597980 244350
rect 597360 244226 597980 244294
rect 597360 244170 597456 244226
rect 597512 244170 597580 244226
rect 597636 244170 597704 244226
rect 597760 244170 597828 244226
rect 597884 244170 597980 244226
rect 597360 244102 597980 244170
rect 597360 244046 597456 244102
rect 597512 244046 597580 244102
rect 597636 244046 597704 244102
rect 597760 244046 597828 244102
rect 597884 244046 597980 244102
rect 597360 243978 597980 244046
rect 597360 243922 597456 243978
rect 597512 243922 597580 243978
rect 597636 243922 597704 243978
rect 597760 243922 597828 243978
rect 597884 243922 597980 243978
rect 597360 226350 597980 243922
rect 597360 226294 597456 226350
rect 597512 226294 597580 226350
rect 597636 226294 597704 226350
rect 597760 226294 597828 226350
rect 597884 226294 597980 226350
rect 597360 226226 597980 226294
rect 597360 226170 597456 226226
rect 597512 226170 597580 226226
rect 597636 226170 597704 226226
rect 597760 226170 597828 226226
rect 597884 226170 597980 226226
rect 597360 226102 597980 226170
rect 597360 226046 597456 226102
rect 597512 226046 597580 226102
rect 597636 226046 597704 226102
rect 597760 226046 597828 226102
rect 597884 226046 597980 226102
rect 597360 225978 597980 226046
rect 597360 225922 597456 225978
rect 597512 225922 597580 225978
rect 597636 225922 597704 225978
rect 597760 225922 597828 225978
rect 597884 225922 597980 225978
rect 597360 208350 597980 225922
rect 597360 208294 597456 208350
rect 597512 208294 597580 208350
rect 597636 208294 597704 208350
rect 597760 208294 597828 208350
rect 597884 208294 597980 208350
rect 597360 208226 597980 208294
rect 597360 208170 597456 208226
rect 597512 208170 597580 208226
rect 597636 208170 597704 208226
rect 597760 208170 597828 208226
rect 597884 208170 597980 208226
rect 597360 208102 597980 208170
rect 597360 208046 597456 208102
rect 597512 208046 597580 208102
rect 597636 208046 597704 208102
rect 597760 208046 597828 208102
rect 597884 208046 597980 208102
rect 597360 207978 597980 208046
rect 597360 207922 597456 207978
rect 597512 207922 597580 207978
rect 597636 207922 597704 207978
rect 597760 207922 597828 207978
rect 597884 207922 597980 207978
rect 597360 190350 597980 207922
rect 597360 190294 597456 190350
rect 597512 190294 597580 190350
rect 597636 190294 597704 190350
rect 597760 190294 597828 190350
rect 597884 190294 597980 190350
rect 597360 190226 597980 190294
rect 597360 190170 597456 190226
rect 597512 190170 597580 190226
rect 597636 190170 597704 190226
rect 597760 190170 597828 190226
rect 597884 190170 597980 190226
rect 597360 190102 597980 190170
rect 597360 190046 597456 190102
rect 597512 190046 597580 190102
rect 597636 190046 597704 190102
rect 597760 190046 597828 190102
rect 597884 190046 597980 190102
rect 597360 189978 597980 190046
rect 597360 189922 597456 189978
rect 597512 189922 597580 189978
rect 597636 189922 597704 189978
rect 597760 189922 597828 189978
rect 597884 189922 597980 189978
rect 597360 172350 597980 189922
rect 597360 172294 597456 172350
rect 597512 172294 597580 172350
rect 597636 172294 597704 172350
rect 597760 172294 597828 172350
rect 597884 172294 597980 172350
rect 597360 172226 597980 172294
rect 597360 172170 597456 172226
rect 597512 172170 597580 172226
rect 597636 172170 597704 172226
rect 597760 172170 597828 172226
rect 597884 172170 597980 172226
rect 597360 172102 597980 172170
rect 597360 172046 597456 172102
rect 597512 172046 597580 172102
rect 597636 172046 597704 172102
rect 597760 172046 597828 172102
rect 597884 172046 597980 172102
rect 597360 171978 597980 172046
rect 597360 171922 597456 171978
rect 597512 171922 597580 171978
rect 597636 171922 597704 171978
rect 597760 171922 597828 171978
rect 597884 171922 597980 171978
rect 597360 154350 597980 171922
rect 597360 154294 597456 154350
rect 597512 154294 597580 154350
rect 597636 154294 597704 154350
rect 597760 154294 597828 154350
rect 597884 154294 597980 154350
rect 597360 154226 597980 154294
rect 597360 154170 597456 154226
rect 597512 154170 597580 154226
rect 597636 154170 597704 154226
rect 597760 154170 597828 154226
rect 597884 154170 597980 154226
rect 597360 154102 597980 154170
rect 597360 154046 597456 154102
rect 597512 154046 597580 154102
rect 597636 154046 597704 154102
rect 597760 154046 597828 154102
rect 597884 154046 597980 154102
rect 597360 153978 597980 154046
rect 597360 153922 597456 153978
rect 597512 153922 597580 153978
rect 597636 153922 597704 153978
rect 597760 153922 597828 153978
rect 597884 153922 597980 153978
rect 597360 136350 597980 153922
rect 597360 136294 597456 136350
rect 597512 136294 597580 136350
rect 597636 136294 597704 136350
rect 597760 136294 597828 136350
rect 597884 136294 597980 136350
rect 597360 136226 597980 136294
rect 597360 136170 597456 136226
rect 597512 136170 597580 136226
rect 597636 136170 597704 136226
rect 597760 136170 597828 136226
rect 597884 136170 597980 136226
rect 597360 136102 597980 136170
rect 597360 136046 597456 136102
rect 597512 136046 597580 136102
rect 597636 136046 597704 136102
rect 597760 136046 597828 136102
rect 597884 136046 597980 136102
rect 597360 135978 597980 136046
rect 597360 135922 597456 135978
rect 597512 135922 597580 135978
rect 597636 135922 597704 135978
rect 597760 135922 597828 135978
rect 597884 135922 597980 135978
rect 597360 118350 597980 135922
rect 597360 118294 597456 118350
rect 597512 118294 597580 118350
rect 597636 118294 597704 118350
rect 597760 118294 597828 118350
rect 597884 118294 597980 118350
rect 597360 118226 597980 118294
rect 597360 118170 597456 118226
rect 597512 118170 597580 118226
rect 597636 118170 597704 118226
rect 597760 118170 597828 118226
rect 597884 118170 597980 118226
rect 597360 118102 597980 118170
rect 597360 118046 597456 118102
rect 597512 118046 597580 118102
rect 597636 118046 597704 118102
rect 597760 118046 597828 118102
rect 597884 118046 597980 118102
rect 597360 117978 597980 118046
rect 597360 117922 597456 117978
rect 597512 117922 597580 117978
rect 597636 117922 597704 117978
rect 597760 117922 597828 117978
rect 597884 117922 597980 117978
rect 597360 100350 597980 117922
rect 597360 100294 597456 100350
rect 597512 100294 597580 100350
rect 597636 100294 597704 100350
rect 597760 100294 597828 100350
rect 597884 100294 597980 100350
rect 597360 100226 597980 100294
rect 597360 100170 597456 100226
rect 597512 100170 597580 100226
rect 597636 100170 597704 100226
rect 597760 100170 597828 100226
rect 597884 100170 597980 100226
rect 597360 100102 597980 100170
rect 597360 100046 597456 100102
rect 597512 100046 597580 100102
rect 597636 100046 597704 100102
rect 597760 100046 597828 100102
rect 597884 100046 597980 100102
rect 597360 99978 597980 100046
rect 597360 99922 597456 99978
rect 597512 99922 597580 99978
rect 597636 99922 597704 99978
rect 597760 99922 597828 99978
rect 597884 99922 597980 99978
rect 597360 82350 597980 99922
rect 597360 82294 597456 82350
rect 597512 82294 597580 82350
rect 597636 82294 597704 82350
rect 597760 82294 597828 82350
rect 597884 82294 597980 82350
rect 597360 82226 597980 82294
rect 597360 82170 597456 82226
rect 597512 82170 597580 82226
rect 597636 82170 597704 82226
rect 597760 82170 597828 82226
rect 597884 82170 597980 82226
rect 597360 82102 597980 82170
rect 597360 82046 597456 82102
rect 597512 82046 597580 82102
rect 597636 82046 597704 82102
rect 597760 82046 597828 82102
rect 597884 82046 597980 82102
rect 597360 81978 597980 82046
rect 597360 81922 597456 81978
rect 597512 81922 597580 81978
rect 597636 81922 597704 81978
rect 597760 81922 597828 81978
rect 597884 81922 597980 81978
rect 597360 64350 597980 81922
rect 597360 64294 597456 64350
rect 597512 64294 597580 64350
rect 597636 64294 597704 64350
rect 597760 64294 597828 64350
rect 597884 64294 597980 64350
rect 597360 64226 597980 64294
rect 597360 64170 597456 64226
rect 597512 64170 597580 64226
rect 597636 64170 597704 64226
rect 597760 64170 597828 64226
rect 597884 64170 597980 64226
rect 597360 64102 597980 64170
rect 597360 64046 597456 64102
rect 597512 64046 597580 64102
rect 597636 64046 597704 64102
rect 597760 64046 597828 64102
rect 597884 64046 597980 64102
rect 597360 63978 597980 64046
rect 597360 63922 597456 63978
rect 597512 63922 597580 63978
rect 597636 63922 597704 63978
rect 597760 63922 597828 63978
rect 597884 63922 597980 63978
rect 597360 46350 597980 63922
rect 597360 46294 597456 46350
rect 597512 46294 597580 46350
rect 597636 46294 597704 46350
rect 597760 46294 597828 46350
rect 597884 46294 597980 46350
rect 597360 46226 597980 46294
rect 597360 46170 597456 46226
rect 597512 46170 597580 46226
rect 597636 46170 597704 46226
rect 597760 46170 597828 46226
rect 597884 46170 597980 46226
rect 597360 46102 597980 46170
rect 597360 46046 597456 46102
rect 597512 46046 597580 46102
rect 597636 46046 597704 46102
rect 597760 46046 597828 46102
rect 597884 46046 597980 46102
rect 597360 45978 597980 46046
rect 597360 45922 597456 45978
rect 597512 45922 597580 45978
rect 597636 45922 597704 45978
rect 597760 45922 597828 45978
rect 597884 45922 597980 45978
rect 597360 28350 597980 45922
rect 597360 28294 597456 28350
rect 597512 28294 597580 28350
rect 597636 28294 597704 28350
rect 597760 28294 597828 28350
rect 597884 28294 597980 28350
rect 597360 28226 597980 28294
rect 597360 28170 597456 28226
rect 597512 28170 597580 28226
rect 597636 28170 597704 28226
rect 597760 28170 597828 28226
rect 597884 28170 597980 28226
rect 597360 28102 597980 28170
rect 597360 28046 597456 28102
rect 597512 28046 597580 28102
rect 597636 28046 597704 28102
rect 597760 28046 597828 28102
rect 597884 28046 597980 28102
rect 597360 27978 597980 28046
rect 597360 27922 597456 27978
rect 597512 27922 597580 27978
rect 597636 27922 597704 27978
rect 597760 27922 597828 27978
rect 597884 27922 597980 27978
rect 597360 10350 597980 27922
rect 597360 10294 597456 10350
rect 597512 10294 597580 10350
rect 597636 10294 597704 10350
rect 597760 10294 597828 10350
rect 597884 10294 597980 10350
rect 597360 10226 597980 10294
rect 597360 10170 597456 10226
rect 597512 10170 597580 10226
rect 597636 10170 597704 10226
rect 597760 10170 597828 10226
rect 597884 10170 597980 10226
rect 597360 10102 597980 10170
rect 597360 10046 597456 10102
rect 597512 10046 597580 10102
rect 597636 10046 597704 10102
rect 597760 10046 597828 10102
rect 597884 10046 597980 10102
rect 597360 9978 597980 10046
rect 597360 9922 597456 9978
rect 597512 9922 597580 9978
rect 597636 9922 597704 9978
rect 597760 9922 597828 9978
rect 597884 9922 597980 9978
rect 592818 -1176 592914 -1120
rect 592970 -1176 593038 -1120
rect 593094 -1176 593162 -1120
rect 593218 -1176 593286 -1120
rect 593342 -1176 593438 -1120
rect 592818 -1244 593438 -1176
rect 592818 -1300 592914 -1244
rect 592970 -1300 593038 -1244
rect 593094 -1300 593162 -1244
rect 593218 -1300 593286 -1244
rect 593342 -1300 593438 -1244
rect 592818 -1368 593438 -1300
rect 592818 -1424 592914 -1368
rect 592970 -1424 593038 -1368
rect 593094 -1424 593162 -1368
rect 593218 -1424 593286 -1368
rect 593342 -1424 593438 -1368
rect 592818 -1492 593438 -1424
rect 592818 -1548 592914 -1492
rect 592970 -1548 593038 -1492
rect 593094 -1548 593162 -1492
rect 593218 -1548 593286 -1492
rect 593342 -1548 593438 -1492
rect 592818 -1644 593438 -1548
rect 597360 -1120 597980 9922
rect 597360 -1176 597456 -1120
rect 597512 -1176 597580 -1120
rect 597636 -1176 597704 -1120
rect 597760 -1176 597828 -1120
rect 597884 -1176 597980 -1120
rect 597360 -1244 597980 -1176
rect 597360 -1300 597456 -1244
rect 597512 -1300 597580 -1244
rect 597636 -1300 597704 -1244
rect 597760 -1300 597828 -1244
rect 597884 -1300 597980 -1244
rect 597360 -1368 597980 -1300
rect 597360 -1424 597456 -1368
rect 597512 -1424 597580 -1368
rect 597636 -1424 597704 -1368
rect 597760 -1424 597828 -1368
rect 597884 -1424 597980 -1368
rect 597360 -1492 597980 -1424
rect 597360 -1548 597456 -1492
rect 597512 -1548 597580 -1492
rect 597636 -1548 597704 -1492
rect 597760 -1548 597828 -1492
rect 597884 -1548 597980 -1492
rect 597360 -1644 597980 -1548
<< via4 >>
rect -1820 598116 -1764 598172
rect -1696 598116 -1640 598172
rect -1572 598116 -1516 598172
rect -1448 598116 -1392 598172
rect -1820 597992 -1764 598048
rect -1696 597992 -1640 598048
rect -1572 597992 -1516 598048
rect -1448 597992 -1392 598048
rect -1820 597868 -1764 597924
rect -1696 597868 -1640 597924
rect -1572 597868 -1516 597924
rect -1448 597868 -1392 597924
rect -1820 597744 -1764 597800
rect -1696 597744 -1640 597800
rect -1572 597744 -1516 597800
rect -1448 597744 -1392 597800
rect -1820 586294 -1764 586350
rect -1696 586294 -1640 586350
rect -1572 586294 -1516 586350
rect -1448 586294 -1392 586350
rect -1820 586170 -1764 586226
rect -1696 586170 -1640 586226
rect -1572 586170 -1516 586226
rect -1448 586170 -1392 586226
rect -1820 586046 -1764 586102
rect -1696 586046 -1640 586102
rect -1572 586046 -1516 586102
rect -1448 586046 -1392 586102
rect -1820 585922 -1764 585978
rect -1696 585922 -1640 585978
rect -1572 585922 -1516 585978
rect -1448 585922 -1392 585978
rect -1820 568294 -1764 568350
rect -1696 568294 -1640 568350
rect -1572 568294 -1516 568350
rect -1448 568294 -1392 568350
rect -1820 568170 -1764 568226
rect -1696 568170 -1640 568226
rect -1572 568170 -1516 568226
rect -1448 568170 -1392 568226
rect -1820 568046 -1764 568102
rect -1696 568046 -1640 568102
rect -1572 568046 -1516 568102
rect -1448 568046 -1392 568102
rect -1820 567922 -1764 567978
rect -1696 567922 -1640 567978
rect -1572 567922 -1516 567978
rect -1448 567922 -1392 567978
rect -1820 550294 -1764 550350
rect -1696 550294 -1640 550350
rect -1572 550294 -1516 550350
rect -1448 550294 -1392 550350
rect -1820 550170 -1764 550226
rect -1696 550170 -1640 550226
rect -1572 550170 -1516 550226
rect -1448 550170 -1392 550226
rect -1820 550046 -1764 550102
rect -1696 550046 -1640 550102
rect -1572 550046 -1516 550102
rect -1448 550046 -1392 550102
rect -1820 549922 -1764 549978
rect -1696 549922 -1640 549978
rect -1572 549922 -1516 549978
rect -1448 549922 -1392 549978
rect -1820 532294 -1764 532350
rect -1696 532294 -1640 532350
rect -1572 532294 -1516 532350
rect -1448 532294 -1392 532350
rect -1820 532170 -1764 532226
rect -1696 532170 -1640 532226
rect -1572 532170 -1516 532226
rect -1448 532170 -1392 532226
rect -1820 532046 -1764 532102
rect -1696 532046 -1640 532102
rect -1572 532046 -1516 532102
rect -1448 532046 -1392 532102
rect -1820 531922 -1764 531978
rect -1696 531922 -1640 531978
rect -1572 531922 -1516 531978
rect -1448 531922 -1392 531978
rect -1820 514294 -1764 514350
rect -1696 514294 -1640 514350
rect -1572 514294 -1516 514350
rect -1448 514294 -1392 514350
rect -1820 514170 -1764 514226
rect -1696 514170 -1640 514226
rect -1572 514170 -1516 514226
rect -1448 514170 -1392 514226
rect -1820 514046 -1764 514102
rect -1696 514046 -1640 514102
rect -1572 514046 -1516 514102
rect -1448 514046 -1392 514102
rect -1820 513922 -1764 513978
rect -1696 513922 -1640 513978
rect -1572 513922 -1516 513978
rect -1448 513922 -1392 513978
rect -1820 496294 -1764 496350
rect -1696 496294 -1640 496350
rect -1572 496294 -1516 496350
rect -1448 496294 -1392 496350
rect -1820 496170 -1764 496226
rect -1696 496170 -1640 496226
rect -1572 496170 -1516 496226
rect -1448 496170 -1392 496226
rect -1820 496046 -1764 496102
rect -1696 496046 -1640 496102
rect -1572 496046 -1516 496102
rect -1448 496046 -1392 496102
rect -1820 495922 -1764 495978
rect -1696 495922 -1640 495978
rect -1572 495922 -1516 495978
rect -1448 495922 -1392 495978
rect -1820 478294 -1764 478350
rect -1696 478294 -1640 478350
rect -1572 478294 -1516 478350
rect -1448 478294 -1392 478350
rect -1820 478170 -1764 478226
rect -1696 478170 -1640 478226
rect -1572 478170 -1516 478226
rect -1448 478170 -1392 478226
rect -1820 478046 -1764 478102
rect -1696 478046 -1640 478102
rect -1572 478046 -1516 478102
rect -1448 478046 -1392 478102
rect -1820 477922 -1764 477978
rect -1696 477922 -1640 477978
rect -1572 477922 -1516 477978
rect -1448 477922 -1392 477978
rect -1820 460294 -1764 460350
rect -1696 460294 -1640 460350
rect -1572 460294 -1516 460350
rect -1448 460294 -1392 460350
rect -1820 460170 -1764 460226
rect -1696 460170 -1640 460226
rect -1572 460170 -1516 460226
rect -1448 460170 -1392 460226
rect -1820 460046 -1764 460102
rect -1696 460046 -1640 460102
rect -1572 460046 -1516 460102
rect -1448 460046 -1392 460102
rect -1820 459922 -1764 459978
rect -1696 459922 -1640 459978
rect -1572 459922 -1516 459978
rect -1448 459922 -1392 459978
rect -1820 442294 -1764 442350
rect -1696 442294 -1640 442350
rect -1572 442294 -1516 442350
rect -1448 442294 -1392 442350
rect -1820 442170 -1764 442226
rect -1696 442170 -1640 442226
rect -1572 442170 -1516 442226
rect -1448 442170 -1392 442226
rect -1820 442046 -1764 442102
rect -1696 442046 -1640 442102
rect -1572 442046 -1516 442102
rect -1448 442046 -1392 442102
rect -1820 441922 -1764 441978
rect -1696 441922 -1640 441978
rect -1572 441922 -1516 441978
rect -1448 441922 -1392 441978
rect -1820 424294 -1764 424350
rect -1696 424294 -1640 424350
rect -1572 424294 -1516 424350
rect -1448 424294 -1392 424350
rect -1820 424170 -1764 424226
rect -1696 424170 -1640 424226
rect -1572 424170 -1516 424226
rect -1448 424170 -1392 424226
rect -1820 424046 -1764 424102
rect -1696 424046 -1640 424102
rect -1572 424046 -1516 424102
rect -1448 424046 -1392 424102
rect -1820 423922 -1764 423978
rect -1696 423922 -1640 423978
rect -1572 423922 -1516 423978
rect -1448 423922 -1392 423978
rect -1820 406294 -1764 406350
rect -1696 406294 -1640 406350
rect -1572 406294 -1516 406350
rect -1448 406294 -1392 406350
rect -1820 406170 -1764 406226
rect -1696 406170 -1640 406226
rect -1572 406170 -1516 406226
rect -1448 406170 -1392 406226
rect -1820 406046 -1764 406102
rect -1696 406046 -1640 406102
rect -1572 406046 -1516 406102
rect -1448 406046 -1392 406102
rect -1820 405922 -1764 405978
rect -1696 405922 -1640 405978
rect -1572 405922 -1516 405978
rect -1448 405922 -1392 405978
rect -1820 388294 -1764 388350
rect -1696 388294 -1640 388350
rect -1572 388294 -1516 388350
rect -1448 388294 -1392 388350
rect -1820 388170 -1764 388226
rect -1696 388170 -1640 388226
rect -1572 388170 -1516 388226
rect -1448 388170 -1392 388226
rect -1820 388046 -1764 388102
rect -1696 388046 -1640 388102
rect -1572 388046 -1516 388102
rect -1448 388046 -1392 388102
rect -1820 387922 -1764 387978
rect -1696 387922 -1640 387978
rect -1572 387922 -1516 387978
rect -1448 387922 -1392 387978
rect -1820 370294 -1764 370350
rect -1696 370294 -1640 370350
rect -1572 370294 -1516 370350
rect -1448 370294 -1392 370350
rect -1820 370170 -1764 370226
rect -1696 370170 -1640 370226
rect -1572 370170 -1516 370226
rect -1448 370170 -1392 370226
rect -1820 370046 -1764 370102
rect -1696 370046 -1640 370102
rect -1572 370046 -1516 370102
rect -1448 370046 -1392 370102
rect -1820 369922 -1764 369978
rect -1696 369922 -1640 369978
rect -1572 369922 -1516 369978
rect -1448 369922 -1392 369978
rect -1820 352294 -1764 352350
rect -1696 352294 -1640 352350
rect -1572 352294 -1516 352350
rect -1448 352294 -1392 352350
rect -1820 352170 -1764 352226
rect -1696 352170 -1640 352226
rect -1572 352170 -1516 352226
rect -1448 352170 -1392 352226
rect -1820 352046 -1764 352102
rect -1696 352046 -1640 352102
rect -1572 352046 -1516 352102
rect -1448 352046 -1392 352102
rect -1820 351922 -1764 351978
rect -1696 351922 -1640 351978
rect -1572 351922 -1516 351978
rect -1448 351922 -1392 351978
rect -1820 334294 -1764 334350
rect -1696 334294 -1640 334350
rect -1572 334294 -1516 334350
rect -1448 334294 -1392 334350
rect -1820 334170 -1764 334226
rect -1696 334170 -1640 334226
rect -1572 334170 -1516 334226
rect -1448 334170 -1392 334226
rect -1820 334046 -1764 334102
rect -1696 334046 -1640 334102
rect -1572 334046 -1516 334102
rect -1448 334046 -1392 334102
rect -1820 333922 -1764 333978
rect -1696 333922 -1640 333978
rect -1572 333922 -1516 333978
rect -1448 333922 -1392 333978
rect -1820 316294 -1764 316350
rect -1696 316294 -1640 316350
rect -1572 316294 -1516 316350
rect -1448 316294 -1392 316350
rect -1820 316170 -1764 316226
rect -1696 316170 -1640 316226
rect -1572 316170 -1516 316226
rect -1448 316170 -1392 316226
rect -1820 316046 -1764 316102
rect -1696 316046 -1640 316102
rect -1572 316046 -1516 316102
rect -1448 316046 -1392 316102
rect -1820 315922 -1764 315978
rect -1696 315922 -1640 315978
rect -1572 315922 -1516 315978
rect -1448 315922 -1392 315978
rect -1820 298294 -1764 298350
rect -1696 298294 -1640 298350
rect -1572 298294 -1516 298350
rect -1448 298294 -1392 298350
rect -1820 298170 -1764 298226
rect -1696 298170 -1640 298226
rect -1572 298170 -1516 298226
rect -1448 298170 -1392 298226
rect -1820 298046 -1764 298102
rect -1696 298046 -1640 298102
rect -1572 298046 -1516 298102
rect -1448 298046 -1392 298102
rect -1820 297922 -1764 297978
rect -1696 297922 -1640 297978
rect -1572 297922 -1516 297978
rect -1448 297922 -1392 297978
rect -1820 280294 -1764 280350
rect -1696 280294 -1640 280350
rect -1572 280294 -1516 280350
rect -1448 280294 -1392 280350
rect -1820 280170 -1764 280226
rect -1696 280170 -1640 280226
rect -1572 280170 -1516 280226
rect -1448 280170 -1392 280226
rect -1820 280046 -1764 280102
rect -1696 280046 -1640 280102
rect -1572 280046 -1516 280102
rect -1448 280046 -1392 280102
rect -1820 279922 -1764 279978
rect -1696 279922 -1640 279978
rect -1572 279922 -1516 279978
rect -1448 279922 -1392 279978
rect -1820 262294 -1764 262350
rect -1696 262294 -1640 262350
rect -1572 262294 -1516 262350
rect -1448 262294 -1392 262350
rect -1820 262170 -1764 262226
rect -1696 262170 -1640 262226
rect -1572 262170 -1516 262226
rect -1448 262170 -1392 262226
rect -1820 262046 -1764 262102
rect -1696 262046 -1640 262102
rect -1572 262046 -1516 262102
rect -1448 262046 -1392 262102
rect -1820 261922 -1764 261978
rect -1696 261922 -1640 261978
rect -1572 261922 -1516 261978
rect -1448 261922 -1392 261978
rect -1820 244294 -1764 244350
rect -1696 244294 -1640 244350
rect -1572 244294 -1516 244350
rect -1448 244294 -1392 244350
rect -1820 244170 -1764 244226
rect -1696 244170 -1640 244226
rect -1572 244170 -1516 244226
rect -1448 244170 -1392 244226
rect -1820 244046 -1764 244102
rect -1696 244046 -1640 244102
rect -1572 244046 -1516 244102
rect -1448 244046 -1392 244102
rect -1820 243922 -1764 243978
rect -1696 243922 -1640 243978
rect -1572 243922 -1516 243978
rect -1448 243922 -1392 243978
rect -1820 226294 -1764 226350
rect -1696 226294 -1640 226350
rect -1572 226294 -1516 226350
rect -1448 226294 -1392 226350
rect -1820 226170 -1764 226226
rect -1696 226170 -1640 226226
rect -1572 226170 -1516 226226
rect -1448 226170 -1392 226226
rect -1820 226046 -1764 226102
rect -1696 226046 -1640 226102
rect -1572 226046 -1516 226102
rect -1448 226046 -1392 226102
rect -1820 225922 -1764 225978
rect -1696 225922 -1640 225978
rect -1572 225922 -1516 225978
rect -1448 225922 -1392 225978
rect -1820 208294 -1764 208350
rect -1696 208294 -1640 208350
rect -1572 208294 -1516 208350
rect -1448 208294 -1392 208350
rect -1820 208170 -1764 208226
rect -1696 208170 -1640 208226
rect -1572 208170 -1516 208226
rect -1448 208170 -1392 208226
rect -1820 208046 -1764 208102
rect -1696 208046 -1640 208102
rect -1572 208046 -1516 208102
rect -1448 208046 -1392 208102
rect -1820 207922 -1764 207978
rect -1696 207922 -1640 207978
rect -1572 207922 -1516 207978
rect -1448 207922 -1392 207978
rect -1820 190294 -1764 190350
rect -1696 190294 -1640 190350
rect -1572 190294 -1516 190350
rect -1448 190294 -1392 190350
rect -1820 190170 -1764 190226
rect -1696 190170 -1640 190226
rect -1572 190170 -1516 190226
rect -1448 190170 -1392 190226
rect -1820 190046 -1764 190102
rect -1696 190046 -1640 190102
rect -1572 190046 -1516 190102
rect -1448 190046 -1392 190102
rect -1820 189922 -1764 189978
rect -1696 189922 -1640 189978
rect -1572 189922 -1516 189978
rect -1448 189922 -1392 189978
rect -1820 172294 -1764 172350
rect -1696 172294 -1640 172350
rect -1572 172294 -1516 172350
rect -1448 172294 -1392 172350
rect -1820 172170 -1764 172226
rect -1696 172170 -1640 172226
rect -1572 172170 -1516 172226
rect -1448 172170 -1392 172226
rect -1820 172046 -1764 172102
rect -1696 172046 -1640 172102
rect -1572 172046 -1516 172102
rect -1448 172046 -1392 172102
rect -1820 171922 -1764 171978
rect -1696 171922 -1640 171978
rect -1572 171922 -1516 171978
rect -1448 171922 -1392 171978
rect -1820 154294 -1764 154350
rect -1696 154294 -1640 154350
rect -1572 154294 -1516 154350
rect -1448 154294 -1392 154350
rect -1820 154170 -1764 154226
rect -1696 154170 -1640 154226
rect -1572 154170 -1516 154226
rect -1448 154170 -1392 154226
rect -1820 154046 -1764 154102
rect -1696 154046 -1640 154102
rect -1572 154046 -1516 154102
rect -1448 154046 -1392 154102
rect -1820 153922 -1764 153978
rect -1696 153922 -1640 153978
rect -1572 153922 -1516 153978
rect -1448 153922 -1392 153978
rect -1820 136294 -1764 136350
rect -1696 136294 -1640 136350
rect -1572 136294 -1516 136350
rect -1448 136294 -1392 136350
rect -1820 136170 -1764 136226
rect -1696 136170 -1640 136226
rect -1572 136170 -1516 136226
rect -1448 136170 -1392 136226
rect -1820 136046 -1764 136102
rect -1696 136046 -1640 136102
rect -1572 136046 -1516 136102
rect -1448 136046 -1392 136102
rect -1820 135922 -1764 135978
rect -1696 135922 -1640 135978
rect -1572 135922 -1516 135978
rect -1448 135922 -1392 135978
rect -1820 118294 -1764 118350
rect -1696 118294 -1640 118350
rect -1572 118294 -1516 118350
rect -1448 118294 -1392 118350
rect -1820 118170 -1764 118226
rect -1696 118170 -1640 118226
rect -1572 118170 -1516 118226
rect -1448 118170 -1392 118226
rect -1820 118046 -1764 118102
rect -1696 118046 -1640 118102
rect -1572 118046 -1516 118102
rect -1448 118046 -1392 118102
rect -1820 117922 -1764 117978
rect -1696 117922 -1640 117978
rect -1572 117922 -1516 117978
rect -1448 117922 -1392 117978
rect -1820 100294 -1764 100350
rect -1696 100294 -1640 100350
rect -1572 100294 -1516 100350
rect -1448 100294 -1392 100350
rect -1820 100170 -1764 100226
rect -1696 100170 -1640 100226
rect -1572 100170 -1516 100226
rect -1448 100170 -1392 100226
rect -1820 100046 -1764 100102
rect -1696 100046 -1640 100102
rect -1572 100046 -1516 100102
rect -1448 100046 -1392 100102
rect -1820 99922 -1764 99978
rect -1696 99922 -1640 99978
rect -1572 99922 -1516 99978
rect -1448 99922 -1392 99978
rect -1820 82294 -1764 82350
rect -1696 82294 -1640 82350
rect -1572 82294 -1516 82350
rect -1448 82294 -1392 82350
rect -1820 82170 -1764 82226
rect -1696 82170 -1640 82226
rect -1572 82170 -1516 82226
rect -1448 82170 -1392 82226
rect -1820 82046 -1764 82102
rect -1696 82046 -1640 82102
rect -1572 82046 -1516 82102
rect -1448 82046 -1392 82102
rect -1820 81922 -1764 81978
rect -1696 81922 -1640 81978
rect -1572 81922 -1516 81978
rect -1448 81922 -1392 81978
rect -1820 64294 -1764 64350
rect -1696 64294 -1640 64350
rect -1572 64294 -1516 64350
rect -1448 64294 -1392 64350
rect -1820 64170 -1764 64226
rect -1696 64170 -1640 64226
rect -1572 64170 -1516 64226
rect -1448 64170 -1392 64226
rect -1820 64046 -1764 64102
rect -1696 64046 -1640 64102
rect -1572 64046 -1516 64102
rect -1448 64046 -1392 64102
rect -1820 63922 -1764 63978
rect -1696 63922 -1640 63978
rect -1572 63922 -1516 63978
rect -1448 63922 -1392 63978
rect -1820 46294 -1764 46350
rect -1696 46294 -1640 46350
rect -1572 46294 -1516 46350
rect -1448 46294 -1392 46350
rect -1820 46170 -1764 46226
rect -1696 46170 -1640 46226
rect -1572 46170 -1516 46226
rect -1448 46170 -1392 46226
rect -1820 46046 -1764 46102
rect -1696 46046 -1640 46102
rect -1572 46046 -1516 46102
rect -1448 46046 -1392 46102
rect -1820 45922 -1764 45978
rect -1696 45922 -1640 45978
rect -1572 45922 -1516 45978
rect -1448 45922 -1392 45978
rect -1820 28294 -1764 28350
rect -1696 28294 -1640 28350
rect -1572 28294 -1516 28350
rect -1448 28294 -1392 28350
rect -1820 28170 -1764 28226
rect -1696 28170 -1640 28226
rect -1572 28170 -1516 28226
rect -1448 28170 -1392 28226
rect -1820 28046 -1764 28102
rect -1696 28046 -1640 28102
rect -1572 28046 -1516 28102
rect -1448 28046 -1392 28102
rect -1820 27922 -1764 27978
rect -1696 27922 -1640 27978
rect -1572 27922 -1516 27978
rect -1448 27922 -1392 27978
rect -1820 10294 -1764 10350
rect -1696 10294 -1640 10350
rect -1572 10294 -1516 10350
rect -1448 10294 -1392 10350
rect -1820 10170 -1764 10226
rect -1696 10170 -1640 10226
rect -1572 10170 -1516 10226
rect -1448 10170 -1392 10226
rect -1820 10046 -1764 10102
rect -1696 10046 -1640 10102
rect -1572 10046 -1516 10102
rect -1448 10046 -1392 10102
rect -1820 9922 -1764 9978
rect -1696 9922 -1640 9978
rect -1572 9922 -1516 9978
rect -1448 9922 -1392 9978
rect -860 597156 -804 597212
rect -736 597156 -680 597212
rect -612 597156 -556 597212
rect -488 597156 -432 597212
rect -860 597032 -804 597088
rect -736 597032 -680 597088
rect -612 597032 -556 597088
rect -488 597032 -432 597088
rect -860 596908 -804 596964
rect -736 596908 -680 596964
rect -612 596908 -556 596964
rect -488 596908 -432 596964
rect -860 596784 -804 596840
rect -736 596784 -680 596840
rect -612 596784 -556 596840
rect -488 596784 -432 596840
rect -860 580294 -804 580350
rect -736 580294 -680 580350
rect -612 580294 -556 580350
rect -488 580294 -432 580350
rect -860 580170 -804 580226
rect -736 580170 -680 580226
rect -612 580170 -556 580226
rect -488 580170 -432 580226
rect -860 580046 -804 580102
rect -736 580046 -680 580102
rect -612 580046 -556 580102
rect -488 580046 -432 580102
rect -860 579922 -804 579978
rect -736 579922 -680 579978
rect -612 579922 -556 579978
rect -488 579922 -432 579978
rect -860 562294 -804 562350
rect -736 562294 -680 562350
rect -612 562294 -556 562350
rect -488 562294 -432 562350
rect -860 562170 -804 562226
rect -736 562170 -680 562226
rect -612 562170 -556 562226
rect -488 562170 -432 562226
rect -860 562046 -804 562102
rect -736 562046 -680 562102
rect -612 562046 -556 562102
rect -488 562046 -432 562102
rect -860 561922 -804 561978
rect -736 561922 -680 561978
rect -612 561922 -556 561978
rect -488 561922 -432 561978
rect -860 544294 -804 544350
rect -736 544294 -680 544350
rect -612 544294 -556 544350
rect -488 544294 -432 544350
rect -860 544170 -804 544226
rect -736 544170 -680 544226
rect -612 544170 -556 544226
rect -488 544170 -432 544226
rect -860 544046 -804 544102
rect -736 544046 -680 544102
rect -612 544046 -556 544102
rect -488 544046 -432 544102
rect -860 543922 -804 543978
rect -736 543922 -680 543978
rect -612 543922 -556 543978
rect -488 543922 -432 543978
rect -860 526294 -804 526350
rect -736 526294 -680 526350
rect -612 526294 -556 526350
rect -488 526294 -432 526350
rect -860 526170 -804 526226
rect -736 526170 -680 526226
rect -612 526170 -556 526226
rect -488 526170 -432 526226
rect -860 526046 -804 526102
rect -736 526046 -680 526102
rect -612 526046 -556 526102
rect -488 526046 -432 526102
rect -860 525922 -804 525978
rect -736 525922 -680 525978
rect -612 525922 -556 525978
rect -488 525922 -432 525978
rect -860 508294 -804 508350
rect -736 508294 -680 508350
rect -612 508294 -556 508350
rect -488 508294 -432 508350
rect -860 508170 -804 508226
rect -736 508170 -680 508226
rect -612 508170 -556 508226
rect -488 508170 -432 508226
rect -860 508046 -804 508102
rect -736 508046 -680 508102
rect -612 508046 -556 508102
rect -488 508046 -432 508102
rect -860 507922 -804 507978
rect -736 507922 -680 507978
rect -612 507922 -556 507978
rect -488 507922 -432 507978
rect -860 490294 -804 490350
rect -736 490294 -680 490350
rect -612 490294 -556 490350
rect -488 490294 -432 490350
rect -860 490170 -804 490226
rect -736 490170 -680 490226
rect -612 490170 -556 490226
rect -488 490170 -432 490226
rect -860 490046 -804 490102
rect -736 490046 -680 490102
rect -612 490046 -556 490102
rect -488 490046 -432 490102
rect -860 489922 -804 489978
rect -736 489922 -680 489978
rect -612 489922 -556 489978
rect -488 489922 -432 489978
rect -860 472294 -804 472350
rect -736 472294 -680 472350
rect -612 472294 -556 472350
rect -488 472294 -432 472350
rect -860 472170 -804 472226
rect -736 472170 -680 472226
rect -612 472170 -556 472226
rect -488 472170 -432 472226
rect -860 472046 -804 472102
rect -736 472046 -680 472102
rect -612 472046 -556 472102
rect -488 472046 -432 472102
rect -860 471922 -804 471978
rect -736 471922 -680 471978
rect -612 471922 -556 471978
rect -488 471922 -432 471978
rect -860 454294 -804 454350
rect -736 454294 -680 454350
rect -612 454294 -556 454350
rect -488 454294 -432 454350
rect -860 454170 -804 454226
rect -736 454170 -680 454226
rect -612 454170 -556 454226
rect -488 454170 -432 454226
rect -860 454046 -804 454102
rect -736 454046 -680 454102
rect -612 454046 -556 454102
rect -488 454046 -432 454102
rect -860 453922 -804 453978
rect -736 453922 -680 453978
rect -612 453922 -556 453978
rect -488 453922 -432 453978
rect -860 436294 -804 436350
rect -736 436294 -680 436350
rect -612 436294 -556 436350
rect -488 436294 -432 436350
rect -860 436170 -804 436226
rect -736 436170 -680 436226
rect -612 436170 -556 436226
rect -488 436170 -432 436226
rect -860 436046 -804 436102
rect -736 436046 -680 436102
rect -612 436046 -556 436102
rect -488 436046 -432 436102
rect -860 435922 -804 435978
rect -736 435922 -680 435978
rect -612 435922 -556 435978
rect -488 435922 -432 435978
rect -860 418294 -804 418350
rect -736 418294 -680 418350
rect -612 418294 -556 418350
rect -488 418294 -432 418350
rect -860 418170 -804 418226
rect -736 418170 -680 418226
rect -612 418170 -556 418226
rect -488 418170 -432 418226
rect -860 418046 -804 418102
rect -736 418046 -680 418102
rect -612 418046 -556 418102
rect -488 418046 -432 418102
rect -860 417922 -804 417978
rect -736 417922 -680 417978
rect -612 417922 -556 417978
rect -488 417922 -432 417978
rect -860 400294 -804 400350
rect -736 400294 -680 400350
rect -612 400294 -556 400350
rect -488 400294 -432 400350
rect -860 400170 -804 400226
rect -736 400170 -680 400226
rect -612 400170 -556 400226
rect -488 400170 -432 400226
rect -860 400046 -804 400102
rect -736 400046 -680 400102
rect -612 400046 -556 400102
rect -488 400046 -432 400102
rect -860 399922 -804 399978
rect -736 399922 -680 399978
rect -612 399922 -556 399978
rect -488 399922 -432 399978
rect -860 382294 -804 382350
rect -736 382294 -680 382350
rect -612 382294 -556 382350
rect -488 382294 -432 382350
rect -860 382170 -804 382226
rect -736 382170 -680 382226
rect -612 382170 -556 382226
rect -488 382170 -432 382226
rect -860 382046 -804 382102
rect -736 382046 -680 382102
rect -612 382046 -556 382102
rect -488 382046 -432 382102
rect -860 381922 -804 381978
rect -736 381922 -680 381978
rect -612 381922 -556 381978
rect -488 381922 -432 381978
rect -860 364294 -804 364350
rect -736 364294 -680 364350
rect -612 364294 -556 364350
rect -488 364294 -432 364350
rect -860 364170 -804 364226
rect -736 364170 -680 364226
rect -612 364170 -556 364226
rect -488 364170 -432 364226
rect -860 364046 -804 364102
rect -736 364046 -680 364102
rect -612 364046 -556 364102
rect -488 364046 -432 364102
rect -860 363922 -804 363978
rect -736 363922 -680 363978
rect -612 363922 -556 363978
rect -488 363922 -432 363978
rect -860 346294 -804 346350
rect -736 346294 -680 346350
rect -612 346294 -556 346350
rect -488 346294 -432 346350
rect -860 346170 -804 346226
rect -736 346170 -680 346226
rect -612 346170 -556 346226
rect -488 346170 -432 346226
rect -860 346046 -804 346102
rect -736 346046 -680 346102
rect -612 346046 -556 346102
rect -488 346046 -432 346102
rect -860 345922 -804 345978
rect -736 345922 -680 345978
rect -612 345922 -556 345978
rect -488 345922 -432 345978
rect -860 328294 -804 328350
rect -736 328294 -680 328350
rect -612 328294 -556 328350
rect -488 328294 -432 328350
rect -860 328170 -804 328226
rect -736 328170 -680 328226
rect -612 328170 -556 328226
rect -488 328170 -432 328226
rect -860 328046 -804 328102
rect -736 328046 -680 328102
rect -612 328046 -556 328102
rect -488 328046 -432 328102
rect -860 327922 -804 327978
rect -736 327922 -680 327978
rect -612 327922 -556 327978
rect -488 327922 -432 327978
rect -860 310294 -804 310350
rect -736 310294 -680 310350
rect -612 310294 -556 310350
rect -488 310294 -432 310350
rect -860 310170 -804 310226
rect -736 310170 -680 310226
rect -612 310170 -556 310226
rect -488 310170 -432 310226
rect -860 310046 -804 310102
rect -736 310046 -680 310102
rect -612 310046 -556 310102
rect -488 310046 -432 310102
rect -860 309922 -804 309978
rect -736 309922 -680 309978
rect -612 309922 -556 309978
rect -488 309922 -432 309978
rect -860 292294 -804 292350
rect -736 292294 -680 292350
rect -612 292294 -556 292350
rect -488 292294 -432 292350
rect -860 292170 -804 292226
rect -736 292170 -680 292226
rect -612 292170 -556 292226
rect -488 292170 -432 292226
rect -860 292046 -804 292102
rect -736 292046 -680 292102
rect -612 292046 -556 292102
rect -488 292046 -432 292102
rect -860 291922 -804 291978
rect -736 291922 -680 291978
rect -612 291922 -556 291978
rect -488 291922 -432 291978
rect -860 274294 -804 274350
rect -736 274294 -680 274350
rect -612 274294 -556 274350
rect -488 274294 -432 274350
rect -860 274170 -804 274226
rect -736 274170 -680 274226
rect -612 274170 -556 274226
rect -488 274170 -432 274226
rect -860 274046 -804 274102
rect -736 274046 -680 274102
rect -612 274046 -556 274102
rect -488 274046 -432 274102
rect -860 273922 -804 273978
rect -736 273922 -680 273978
rect -612 273922 -556 273978
rect -488 273922 -432 273978
rect -860 256294 -804 256350
rect -736 256294 -680 256350
rect -612 256294 -556 256350
rect -488 256294 -432 256350
rect -860 256170 -804 256226
rect -736 256170 -680 256226
rect -612 256170 -556 256226
rect -488 256170 -432 256226
rect -860 256046 -804 256102
rect -736 256046 -680 256102
rect -612 256046 -556 256102
rect -488 256046 -432 256102
rect -860 255922 -804 255978
rect -736 255922 -680 255978
rect -612 255922 -556 255978
rect -488 255922 -432 255978
rect -860 238294 -804 238350
rect -736 238294 -680 238350
rect -612 238294 -556 238350
rect -488 238294 -432 238350
rect -860 238170 -804 238226
rect -736 238170 -680 238226
rect -612 238170 -556 238226
rect -488 238170 -432 238226
rect -860 238046 -804 238102
rect -736 238046 -680 238102
rect -612 238046 -556 238102
rect -488 238046 -432 238102
rect -860 237922 -804 237978
rect -736 237922 -680 237978
rect -612 237922 -556 237978
rect -488 237922 -432 237978
rect -860 220294 -804 220350
rect -736 220294 -680 220350
rect -612 220294 -556 220350
rect -488 220294 -432 220350
rect -860 220170 -804 220226
rect -736 220170 -680 220226
rect -612 220170 -556 220226
rect -488 220170 -432 220226
rect -860 220046 -804 220102
rect -736 220046 -680 220102
rect -612 220046 -556 220102
rect -488 220046 -432 220102
rect -860 219922 -804 219978
rect -736 219922 -680 219978
rect -612 219922 -556 219978
rect -488 219922 -432 219978
rect -860 202294 -804 202350
rect -736 202294 -680 202350
rect -612 202294 -556 202350
rect -488 202294 -432 202350
rect -860 202170 -804 202226
rect -736 202170 -680 202226
rect -612 202170 -556 202226
rect -488 202170 -432 202226
rect -860 202046 -804 202102
rect -736 202046 -680 202102
rect -612 202046 -556 202102
rect -488 202046 -432 202102
rect -860 201922 -804 201978
rect -736 201922 -680 201978
rect -612 201922 -556 201978
rect -488 201922 -432 201978
rect -860 184294 -804 184350
rect -736 184294 -680 184350
rect -612 184294 -556 184350
rect -488 184294 -432 184350
rect -860 184170 -804 184226
rect -736 184170 -680 184226
rect -612 184170 -556 184226
rect -488 184170 -432 184226
rect -860 184046 -804 184102
rect -736 184046 -680 184102
rect -612 184046 -556 184102
rect -488 184046 -432 184102
rect -860 183922 -804 183978
rect -736 183922 -680 183978
rect -612 183922 -556 183978
rect -488 183922 -432 183978
rect -860 166294 -804 166350
rect -736 166294 -680 166350
rect -612 166294 -556 166350
rect -488 166294 -432 166350
rect -860 166170 -804 166226
rect -736 166170 -680 166226
rect -612 166170 -556 166226
rect -488 166170 -432 166226
rect -860 166046 -804 166102
rect -736 166046 -680 166102
rect -612 166046 -556 166102
rect -488 166046 -432 166102
rect -860 165922 -804 165978
rect -736 165922 -680 165978
rect -612 165922 -556 165978
rect -488 165922 -432 165978
rect -860 148294 -804 148350
rect -736 148294 -680 148350
rect -612 148294 -556 148350
rect -488 148294 -432 148350
rect -860 148170 -804 148226
rect -736 148170 -680 148226
rect -612 148170 -556 148226
rect -488 148170 -432 148226
rect -860 148046 -804 148102
rect -736 148046 -680 148102
rect -612 148046 -556 148102
rect -488 148046 -432 148102
rect -860 147922 -804 147978
rect -736 147922 -680 147978
rect -612 147922 -556 147978
rect -488 147922 -432 147978
rect -860 130294 -804 130350
rect -736 130294 -680 130350
rect -612 130294 -556 130350
rect -488 130294 -432 130350
rect -860 130170 -804 130226
rect -736 130170 -680 130226
rect -612 130170 -556 130226
rect -488 130170 -432 130226
rect -860 130046 -804 130102
rect -736 130046 -680 130102
rect -612 130046 -556 130102
rect -488 130046 -432 130102
rect -860 129922 -804 129978
rect -736 129922 -680 129978
rect -612 129922 -556 129978
rect -488 129922 -432 129978
rect -860 112294 -804 112350
rect -736 112294 -680 112350
rect -612 112294 -556 112350
rect -488 112294 -432 112350
rect -860 112170 -804 112226
rect -736 112170 -680 112226
rect -612 112170 -556 112226
rect -488 112170 -432 112226
rect -860 112046 -804 112102
rect -736 112046 -680 112102
rect -612 112046 -556 112102
rect -488 112046 -432 112102
rect -860 111922 -804 111978
rect -736 111922 -680 111978
rect -612 111922 -556 111978
rect -488 111922 -432 111978
rect -860 94294 -804 94350
rect -736 94294 -680 94350
rect -612 94294 -556 94350
rect -488 94294 -432 94350
rect -860 94170 -804 94226
rect -736 94170 -680 94226
rect -612 94170 -556 94226
rect -488 94170 -432 94226
rect -860 94046 -804 94102
rect -736 94046 -680 94102
rect -612 94046 -556 94102
rect -488 94046 -432 94102
rect -860 93922 -804 93978
rect -736 93922 -680 93978
rect -612 93922 -556 93978
rect -488 93922 -432 93978
rect -860 76294 -804 76350
rect -736 76294 -680 76350
rect -612 76294 -556 76350
rect -488 76294 -432 76350
rect -860 76170 -804 76226
rect -736 76170 -680 76226
rect -612 76170 -556 76226
rect -488 76170 -432 76226
rect -860 76046 -804 76102
rect -736 76046 -680 76102
rect -612 76046 -556 76102
rect -488 76046 -432 76102
rect -860 75922 -804 75978
rect -736 75922 -680 75978
rect -612 75922 -556 75978
rect -488 75922 -432 75978
rect -860 58294 -804 58350
rect -736 58294 -680 58350
rect -612 58294 -556 58350
rect -488 58294 -432 58350
rect -860 58170 -804 58226
rect -736 58170 -680 58226
rect -612 58170 -556 58226
rect -488 58170 -432 58226
rect -860 58046 -804 58102
rect -736 58046 -680 58102
rect -612 58046 -556 58102
rect -488 58046 -432 58102
rect -860 57922 -804 57978
rect -736 57922 -680 57978
rect -612 57922 -556 57978
rect -488 57922 -432 57978
rect -860 40294 -804 40350
rect -736 40294 -680 40350
rect -612 40294 -556 40350
rect -488 40294 -432 40350
rect -860 40170 -804 40226
rect -736 40170 -680 40226
rect -612 40170 -556 40226
rect -488 40170 -432 40226
rect -860 40046 -804 40102
rect -736 40046 -680 40102
rect -612 40046 -556 40102
rect -488 40046 -432 40102
rect -860 39922 -804 39978
rect -736 39922 -680 39978
rect -612 39922 -556 39978
rect -488 39922 -432 39978
rect -860 22294 -804 22350
rect -736 22294 -680 22350
rect -612 22294 -556 22350
rect -488 22294 -432 22350
rect -860 22170 -804 22226
rect -736 22170 -680 22226
rect -612 22170 -556 22226
rect -488 22170 -432 22226
rect -860 22046 -804 22102
rect -736 22046 -680 22102
rect -612 22046 -556 22102
rect -488 22046 -432 22102
rect -860 21922 -804 21978
rect -736 21922 -680 21978
rect -612 21922 -556 21978
rect -488 21922 -432 21978
rect -860 4294 -804 4350
rect -736 4294 -680 4350
rect -612 4294 -556 4350
rect -488 4294 -432 4350
rect -860 4170 -804 4226
rect -736 4170 -680 4226
rect -612 4170 -556 4226
rect -488 4170 -432 4226
rect -860 4046 -804 4102
rect -736 4046 -680 4102
rect -612 4046 -556 4102
rect -488 4046 -432 4102
rect -860 3922 -804 3978
rect -736 3922 -680 3978
rect -612 3922 -556 3978
rect -488 3922 -432 3978
rect -860 -216 -804 -160
rect -736 -216 -680 -160
rect -612 -216 -556 -160
rect -488 -216 -432 -160
rect -860 -340 -804 -284
rect -736 -340 -680 -284
rect -612 -340 -556 -284
rect -488 -340 -432 -284
rect -860 -464 -804 -408
rect -736 -464 -680 -408
rect -612 -464 -556 -408
rect -488 -464 -432 -408
rect -860 -588 -804 -532
rect -736 -588 -680 -532
rect -612 -588 -556 -532
rect -488 -588 -432 -532
rect 5514 597156 5570 597212
rect 5638 597156 5694 597212
rect 5762 597156 5818 597212
rect 5886 597156 5942 597212
rect 5514 597032 5570 597088
rect 5638 597032 5694 597088
rect 5762 597032 5818 597088
rect 5886 597032 5942 597088
rect 5514 596908 5570 596964
rect 5638 596908 5694 596964
rect 5762 596908 5818 596964
rect 5886 596908 5942 596964
rect 5514 596784 5570 596840
rect 5638 596784 5694 596840
rect 5762 596784 5818 596840
rect 5886 596784 5942 596840
rect 5514 580294 5570 580350
rect 5638 580294 5694 580350
rect 5762 580294 5818 580350
rect 5886 580294 5942 580350
rect 5514 580170 5570 580226
rect 5638 580170 5694 580226
rect 5762 580170 5818 580226
rect 5886 580170 5942 580226
rect 5514 580046 5570 580102
rect 5638 580046 5694 580102
rect 5762 580046 5818 580102
rect 5886 580046 5942 580102
rect 5514 579922 5570 579978
rect 5638 579922 5694 579978
rect 5762 579922 5818 579978
rect 5886 579922 5942 579978
rect 5514 562294 5570 562350
rect 5638 562294 5694 562350
rect 5762 562294 5818 562350
rect 5886 562294 5942 562350
rect 5514 562170 5570 562226
rect 5638 562170 5694 562226
rect 5762 562170 5818 562226
rect 5886 562170 5942 562226
rect 5514 562046 5570 562102
rect 5638 562046 5694 562102
rect 5762 562046 5818 562102
rect 5886 562046 5942 562102
rect 5514 561922 5570 561978
rect 5638 561922 5694 561978
rect 5762 561922 5818 561978
rect 5886 561922 5942 561978
rect 5514 544294 5570 544350
rect 5638 544294 5694 544350
rect 5762 544294 5818 544350
rect 5886 544294 5942 544350
rect 5514 544170 5570 544226
rect 5638 544170 5694 544226
rect 5762 544170 5818 544226
rect 5886 544170 5942 544226
rect 5514 544046 5570 544102
rect 5638 544046 5694 544102
rect 5762 544046 5818 544102
rect 5886 544046 5942 544102
rect 5514 543922 5570 543978
rect 5638 543922 5694 543978
rect 5762 543922 5818 543978
rect 5886 543922 5942 543978
rect 5514 526294 5570 526350
rect 5638 526294 5694 526350
rect 5762 526294 5818 526350
rect 5886 526294 5942 526350
rect 5514 526170 5570 526226
rect 5638 526170 5694 526226
rect 5762 526170 5818 526226
rect 5886 526170 5942 526226
rect 5514 526046 5570 526102
rect 5638 526046 5694 526102
rect 5762 526046 5818 526102
rect 5886 526046 5942 526102
rect 5514 525922 5570 525978
rect 5638 525922 5694 525978
rect 5762 525922 5818 525978
rect 5886 525922 5942 525978
rect 5514 508294 5570 508350
rect 5638 508294 5694 508350
rect 5762 508294 5818 508350
rect 5886 508294 5942 508350
rect 5514 508170 5570 508226
rect 5638 508170 5694 508226
rect 5762 508170 5818 508226
rect 5886 508170 5942 508226
rect 5514 508046 5570 508102
rect 5638 508046 5694 508102
rect 5762 508046 5818 508102
rect 5886 508046 5942 508102
rect 5514 507922 5570 507978
rect 5638 507922 5694 507978
rect 5762 507922 5818 507978
rect 5886 507922 5942 507978
rect 5514 490294 5570 490350
rect 5638 490294 5694 490350
rect 5762 490294 5818 490350
rect 5886 490294 5942 490350
rect 5514 490170 5570 490226
rect 5638 490170 5694 490226
rect 5762 490170 5818 490226
rect 5886 490170 5942 490226
rect 5514 490046 5570 490102
rect 5638 490046 5694 490102
rect 5762 490046 5818 490102
rect 5886 490046 5942 490102
rect 5514 489922 5570 489978
rect 5638 489922 5694 489978
rect 5762 489922 5818 489978
rect 5886 489922 5942 489978
rect 5514 472294 5570 472350
rect 5638 472294 5694 472350
rect 5762 472294 5818 472350
rect 5886 472294 5942 472350
rect 5514 472170 5570 472226
rect 5638 472170 5694 472226
rect 5762 472170 5818 472226
rect 5886 472170 5942 472226
rect 5514 472046 5570 472102
rect 5638 472046 5694 472102
rect 5762 472046 5818 472102
rect 5886 472046 5942 472102
rect 5514 471922 5570 471978
rect 5638 471922 5694 471978
rect 5762 471922 5818 471978
rect 5886 471922 5942 471978
rect 5514 454294 5570 454350
rect 5638 454294 5694 454350
rect 5762 454294 5818 454350
rect 5886 454294 5942 454350
rect 5514 454170 5570 454226
rect 5638 454170 5694 454226
rect 5762 454170 5818 454226
rect 5886 454170 5942 454226
rect 5514 454046 5570 454102
rect 5638 454046 5694 454102
rect 5762 454046 5818 454102
rect 5886 454046 5942 454102
rect 5514 453922 5570 453978
rect 5638 453922 5694 453978
rect 5762 453922 5818 453978
rect 5886 453922 5942 453978
rect 5514 436294 5570 436350
rect 5638 436294 5694 436350
rect 5762 436294 5818 436350
rect 5886 436294 5942 436350
rect 5514 436170 5570 436226
rect 5638 436170 5694 436226
rect 5762 436170 5818 436226
rect 5886 436170 5942 436226
rect 5514 436046 5570 436102
rect 5638 436046 5694 436102
rect 5762 436046 5818 436102
rect 5886 436046 5942 436102
rect 5514 435922 5570 435978
rect 5638 435922 5694 435978
rect 5762 435922 5818 435978
rect 5886 435922 5942 435978
rect 5514 418294 5570 418350
rect 5638 418294 5694 418350
rect 5762 418294 5818 418350
rect 5886 418294 5942 418350
rect 5514 418170 5570 418226
rect 5638 418170 5694 418226
rect 5762 418170 5818 418226
rect 5886 418170 5942 418226
rect 5514 418046 5570 418102
rect 5638 418046 5694 418102
rect 5762 418046 5818 418102
rect 5886 418046 5942 418102
rect 5514 417922 5570 417978
rect 5638 417922 5694 417978
rect 5762 417922 5818 417978
rect 5886 417922 5942 417978
rect 5514 400294 5570 400350
rect 5638 400294 5694 400350
rect 5762 400294 5818 400350
rect 5886 400294 5942 400350
rect 5514 400170 5570 400226
rect 5638 400170 5694 400226
rect 5762 400170 5818 400226
rect 5886 400170 5942 400226
rect 5514 400046 5570 400102
rect 5638 400046 5694 400102
rect 5762 400046 5818 400102
rect 5886 400046 5942 400102
rect 5514 399922 5570 399978
rect 5638 399922 5694 399978
rect 5762 399922 5818 399978
rect 5886 399922 5942 399978
rect 5514 382294 5570 382350
rect 5638 382294 5694 382350
rect 5762 382294 5818 382350
rect 5886 382294 5942 382350
rect 5514 382170 5570 382226
rect 5638 382170 5694 382226
rect 5762 382170 5818 382226
rect 5886 382170 5942 382226
rect 5514 382046 5570 382102
rect 5638 382046 5694 382102
rect 5762 382046 5818 382102
rect 5886 382046 5942 382102
rect 5514 381922 5570 381978
rect 5638 381922 5694 381978
rect 5762 381922 5818 381978
rect 5886 381922 5942 381978
rect 5514 364294 5570 364350
rect 5638 364294 5694 364350
rect 5762 364294 5818 364350
rect 5886 364294 5942 364350
rect 5514 364170 5570 364226
rect 5638 364170 5694 364226
rect 5762 364170 5818 364226
rect 5886 364170 5942 364226
rect 5514 364046 5570 364102
rect 5638 364046 5694 364102
rect 5762 364046 5818 364102
rect 5886 364046 5942 364102
rect 5514 363922 5570 363978
rect 5638 363922 5694 363978
rect 5762 363922 5818 363978
rect 5886 363922 5942 363978
rect 5514 346294 5570 346350
rect 5638 346294 5694 346350
rect 5762 346294 5818 346350
rect 5886 346294 5942 346350
rect 5514 346170 5570 346226
rect 5638 346170 5694 346226
rect 5762 346170 5818 346226
rect 5886 346170 5942 346226
rect 5514 346046 5570 346102
rect 5638 346046 5694 346102
rect 5762 346046 5818 346102
rect 5886 346046 5942 346102
rect 5514 345922 5570 345978
rect 5638 345922 5694 345978
rect 5762 345922 5818 345978
rect 5886 345922 5942 345978
rect 5514 328294 5570 328350
rect 5638 328294 5694 328350
rect 5762 328294 5818 328350
rect 5886 328294 5942 328350
rect 5514 328170 5570 328226
rect 5638 328170 5694 328226
rect 5762 328170 5818 328226
rect 5886 328170 5942 328226
rect 5514 328046 5570 328102
rect 5638 328046 5694 328102
rect 5762 328046 5818 328102
rect 5886 328046 5942 328102
rect 5514 327922 5570 327978
rect 5638 327922 5694 327978
rect 5762 327922 5818 327978
rect 5886 327922 5942 327978
rect 5514 310294 5570 310350
rect 5638 310294 5694 310350
rect 5762 310294 5818 310350
rect 5886 310294 5942 310350
rect 5514 310170 5570 310226
rect 5638 310170 5694 310226
rect 5762 310170 5818 310226
rect 5886 310170 5942 310226
rect 5514 310046 5570 310102
rect 5638 310046 5694 310102
rect 5762 310046 5818 310102
rect 5886 310046 5942 310102
rect 5514 309922 5570 309978
rect 5638 309922 5694 309978
rect 5762 309922 5818 309978
rect 5886 309922 5942 309978
rect 5514 292294 5570 292350
rect 5638 292294 5694 292350
rect 5762 292294 5818 292350
rect 5886 292294 5942 292350
rect 5514 292170 5570 292226
rect 5638 292170 5694 292226
rect 5762 292170 5818 292226
rect 5886 292170 5942 292226
rect 5514 292046 5570 292102
rect 5638 292046 5694 292102
rect 5762 292046 5818 292102
rect 5886 292046 5942 292102
rect 5514 291922 5570 291978
rect 5638 291922 5694 291978
rect 5762 291922 5818 291978
rect 5886 291922 5942 291978
rect 5514 274294 5570 274350
rect 5638 274294 5694 274350
rect 5762 274294 5818 274350
rect 5886 274294 5942 274350
rect 5514 274170 5570 274226
rect 5638 274170 5694 274226
rect 5762 274170 5818 274226
rect 5886 274170 5942 274226
rect 5514 274046 5570 274102
rect 5638 274046 5694 274102
rect 5762 274046 5818 274102
rect 5886 274046 5942 274102
rect 5514 273922 5570 273978
rect 5638 273922 5694 273978
rect 5762 273922 5818 273978
rect 5886 273922 5942 273978
rect 5514 256294 5570 256350
rect 5638 256294 5694 256350
rect 5762 256294 5818 256350
rect 5886 256294 5942 256350
rect 5514 256170 5570 256226
rect 5638 256170 5694 256226
rect 5762 256170 5818 256226
rect 5886 256170 5942 256226
rect 5514 256046 5570 256102
rect 5638 256046 5694 256102
rect 5762 256046 5818 256102
rect 5886 256046 5942 256102
rect 5514 255922 5570 255978
rect 5638 255922 5694 255978
rect 5762 255922 5818 255978
rect 5886 255922 5942 255978
rect 5514 238294 5570 238350
rect 5638 238294 5694 238350
rect 5762 238294 5818 238350
rect 5886 238294 5942 238350
rect 5514 238170 5570 238226
rect 5638 238170 5694 238226
rect 5762 238170 5818 238226
rect 5886 238170 5942 238226
rect 5514 238046 5570 238102
rect 5638 238046 5694 238102
rect 5762 238046 5818 238102
rect 5886 238046 5942 238102
rect 5514 237922 5570 237978
rect 5638 237922 5694 237978
rect 5762 237922 5818 237978
rect 5886 237922 5942 237978
rect 5514 220294 5570 220350
rect 5638 220294 5694 220350
rect 5762 220294 5818 220350
rect 5886 220294 5942 220350
rect 5514 220170 5570 220226
rect 5638 220170 5694 220226
rect 5762 220170 5818 220226
rect 5886 220170 5942 220226
rect 5514 220046 5570 220102
rect 5638 220046 5694 220102
rect 5762 220046 5818 220102
rect 5886 220046 5942 220102
rect 5514 219922 5570 219978
rect 5638 219922 5694 219978
rect 5762 219922 5818 219978
rect 5886 219922 5942 219978
rect 5514 202294 5570 202350
rect 5638 202294 5694 202350
rect 5762 202294 5818 202350
rect 5886 202294 5942 202350
rect 5514 202170 5570 202226
rect 5638 202170 5694 202226
rect 5762 202170 5818 202226
rect 5886 202170 5942 202226
rect 5514 202046 5570 202102
rect 5638 202046 5694 202102
rect 5762 202046 5818 202102
rect 5886 202046 5942 202102
rect 5514 201922 5570 201978
rect 5638 201922 5694 201978
rect 5762 201922 5818 201978
rect 5886 201922 5942 201978
rect 5514 184294 5570 184350
rect 5638 184294 5694 184350
rect 5762 184294 5818 184350
rect 5886 184294 5942 184350
rect 5514 184170 5570 184226
rect 5638 184170 5694 184226
rect 5762 184170 5818 184226
rect 5886 184170 5942 184226
rect 5514 184046 5570 184102
rect 5638 184046 5694 184102
rect 5762 184046 5818 184102
rect 5886 184046 5942 184102
rect 5514 183922 5570 183978
rect 5638 183922 5694 183978
rect 5762 183922 5818 183978
rect 5886 183922 5942 183978
rect 5514 166294 5570 166350
rect 5638 166294 5694 166350
rect 5762 166294 5818 166350
rect 5886 166294 5942 166350
rect 5514 166170 5570 166226
rect 5638 166170 5694 166226
rect 5762 166170 5818 166226
rect 5886 166170 5942 166226
rect 5514 166046 5570 166102
rect 5638 166046 5694 166102
rect 5762 166046 5818 166102
rect 5886 166046 5942 166102
rect 5514 165922 5570 165978
rect 5638 165922 5694 165978
rect 5762 165922 5818 165978
rect 5886 165922 5942 165978
rect 5514 148294 5570 148350
rect 5638 148294 5694 148350
rect 5762 148294 5818 148350
rect 5886 148294 5942 148350
rect 5514 148170 5570 148226
rect 5638 148170 5694 148226
rect 5762 148170 5818 148226
rect 5886 148170 5942 148226
rect 5514 148046 5570 148102
rect 5638 148046 5694 148102
rect 5762 148046 5818 148102
rect 5886 148046 5942 148102
rect 5514 147922 5570 147978
rect 5638 147922 5694 147978
rect 5762 147922 5818 147978
rect 5886 147922 5942 147978
rect 5514 130294 5570 130350
rect 5638 130294 5694 130350
rect 5762 130294 5818 130350
rect 5886 130294 5942 130350
rect 5514 130170 5570 130226
rect 5638 130170 5694 130226
rect 5762 130170 5818 130226
rect 5886 130170 5942 130226
rect 5514 130046 5570 130102
rect 5638 130046 5694 130102
rect 5762 130046 5818 130102
rect 5886 130046 5942 130102
rect 5514 129922 5570 129978
rect 5638 129922 5694 129978
rect 5762 129922 5818 129978
rect 5886 129922 5942 129978
rect 5514 112294 5570 112350
rect 5638 112294 5694 112350
rect 5762 112294 5818 112350
rect 5886 112294 5942 112350
rect 5514 112170 5570 112226
rect 5638 112170 5694 112226
rect 5762 112170 5818 112226
rect 5886 112170 5942 112226
rect 5514 112046 5570 112102
rect 5638 112046 5694 112102
rect 5762 112046 5818 112102
rect 5886 112046 5942 112102
rect 5514 111922 5570 111978
rect 5638 111922 5694 111978
rect 5762 111922 5818 111978
rect 5886 111922 5942 111978
rect 5514 94294 5570 94350
rect 5638 94294 5694 94350
rect 5762 94294 5818 94350
rect 5886 94294 5942 94350
rect 5514 94170 5570 94226
rect 5638 94170 5694 94226
rect 5762 94170 5818 94226
rect 5886 94170 5942 94226
rect 5514 94046 5570 94102
rect 5638 94046 5694 94102
rect 5762 94046 5818 94102
rect 5886 94046 5942 94102
rect 5514 93922 5570 93978
rect 5638 93922 5694 93978
rect 5762 93922 5818 93978
rect 5886 93922 5942 93978
rect 5514 76294 5570 76350
rect 5638 76294 5694 76350
rect 5762 76294 5818 76350
rect 5886 76294 5942 76350
rect 5514 76170 5570 76226
rect 5638 76170 5694 76226
rect 5762 76170 5818 76226
rect 5886 76170 5942 76226
rect 5514 76046 5570 76102
rect 5638 76046 5694 76102
rect 5762 76046 5818 76102
rect 5886 76046 5942 76102
rect 5514 75922 5570 75978
rect 5638 75922 5694 75978
rect 5762 75922 5818 75978
rect 5886 75922 5942 75978
rect 5514 58294 5570 58350
rect 5638 58294 5694 58350
rect 5762 58294 5818 58350
rect 5886 58294 5942 58350
rect 5514 58170 5570 58226
rect 5638 58170 5694 58226
rect 5762 58170 5818 58226
rect 5886 58170 5942 58226
rect 5514 58046 5570 58102
rect 5638 58046 5694 58102
rect 5762 58046 5818 58102
rect 5886 58046 5942 58102
rect 5514 57922 5570 57978
rect 5638 57922 5694 57978
rect 5762 57922 5818 57978
rect 5886 57922 5942 57978
rect 5514 40294 5570 40350
rect 5638 40294 5694 40350
rect 5762 40294 5818 40350
rect 5886 40294 5942 40350
rect 5514 40170 5570 40226
rect 5638 40170 5694 40226
rect 5762 40170 5818 40226
rect 5886 40170 5942 40226
rect 5514 40046 5570 40102
rect 5638 40046 5694 40102
rect 5762 40046 5818 40102
rect 5886 40046 5942 40102
rect 5514 39922 5570 39978
rect 5638 39922 5694 39978
rect 5762 39922 5818 39978
rect 5886 39922 5942 39978
rect 5514 22294 5570 22350
rect 5638 22294 5694 22350
rect 5762 22294 5818 22350
rect 5886 22294 5942 22350
rect 5514 22170 5570 22226
rect 5638 22170 5694 22226
rect 5762 22170 5818 22226
rect 5886 22170 5942 22226
rect 5514 22046 5570 22102
rect 5638 22046 5694 22102
rect 5762 22046 5818 22102
rect 5886 22046 5942 22102
rect 5514 21922 5570 21978
rect 5638 21922 5694 21978
rect 5762 21922 5818 21978
rect 5886 21922 5942 21978
rect 5514 4294 5570 4350
rect 5638 4294 5694 4350
rect 5762 4294 5818 4350
rect 5886 4294 5942 4350
rect 5514 4170 5570 4226
rect 5638 4170 5694 4226
rect 5762 4170 5818 4226
rect 5886 4170 5942 4226
rect 5514 4046 5570 4102
rect 5638 4046 5694 4102
rect 5762 4046 5818 4102
rect 5886 4046 5942 4102
rect 5514 3922 5570 3978
rect 5638 3922 5694 3978
rect 5762 3922 5818 3978
rect 5886 3922 5942 3978
rect 5514 -216 5570 -160
rect 5638 -216 5694 -160
rect 5762 -216 5818 -160
rect 5886 -216 5942 -160
rect 5514 -340 5570 -284
rect 5638 -340 5694 -284
rect 5762 -340 5818 -284
rect 5886 -340 5942 -284
rect 5514 -464 5570 -408
rect 5638 -464 5694 -408
rect 5762 -464 5818 -408
rect 5886 -464 5942 -408
rect 5514 -588 5570 -532
rect 5638 -588 5694 -532
rect 5762 -588 5818 -532
rect 5886 -588 5942 -532
rect -1820 -1176 -1764 -1120
rect -1696 -1176 -1640 -1120
rect -1572 -1176 -1516 -1120
rect -1448 -1176 -1392 -1120
rect -1820 -1300 -1764 -1244
rect -1696 -1300 -1640 -1244
rect -1572 -1300 -1516 -1244
rect -1448 -1300 -1392 -1244
rect -1820 -1424 -1764 -1368
rect -1696 -1424 -1640 -1368
rect -1572 -1424 -1516 -1368
rect -1448 -1424 -1392 -1368
rect -1820 -1548 -1764 -1492
rect -1696 -1548 -1640 -1492
rect -1572 -1548 -1516 -1492
rect -1448 -1548 -1392 -1492
rect 9234 598116 9290 598172
rect 9358 598116 9414 598172
rect 9482 598116 9538 598172
rect 9606 598116 9662 598172
rect 9234 597992 9290 598048
rect 9358 597992 9414 598048
rect 9482 597992 9538 598048
rect 9606 597992 9662 598048
rect 9234 597868 9290 597924
rect 9358 597868 9414 597924
rect 9482 597868 9538 597924
rect 9606 597868 9662 597924
rect 9234 597744 9290 597800
rect 9358 597744 9414 597800
rect 9482 597744 9538 597800
rect 9606 597744 9662 597800
rect 9234 586294 9290 586350
rect 9358 586294 9414 586350
rect 9482 586294 9538 586350
rect 9606 586294 9662 586350
rect 9234 586170 9290 586226
rect 9358 586170 9414 586226
rect 9482 586170 9538 586226
rect 9606 586170 9662 586226
rect 9234 586046 9290 586102
rect 9358 586046 9414 586102
rect 9482 586046 9538 586102
rect 9606 586046 9662 586102
rect 9234 585922 9290 585978
rect 9358 585922 9414 585978
rect 9482 585922 9538 585978
rect 9606 585922 9662 585978
rect 9234 568294 9290 568350
rect 9358 568294 9414 568350
rect 9482 568294 9538 568350
rect 9606 568294 9662 568350
rect 9234 568170 9290 568226
rect 9358 568170 9414 568226
rect 9482 568170 9538 568226
rect 9606 568170 9662 568226
rect 9234 568046 9290 568102
rect 9358 568046 9414 568102
rect 9482 568046 9538 568102
rect 9606 568046 9662 568102
rect 9234 567922 9290 567978
rect 9358 567922 9414 567978
rect 9482 567922 9538 567978
rect 9606 567922 9662 567978
rect 36234 597156 36290 597212
rect 36358 597156 36414 597212
rect 36482 597156 36538 597212
rect 36606 597156 36662 597212
rect 36234 597032 36290 597088
rect 36358 597032 36414 597088
rect 36482 597032 36538 597088
rect 36606 597032 36662 597088
rect 36234 596908 36290 596964
rect 36358 596908 36414 596964
rect 36482 596908 36538 596964
rect 36606 596908 36662 596964
rect 36234 596784 36290 596840
rect 36358 596784 36414 596840
rect 36482 596784 36538 596840
rect 36606 596784 36662 596840
rect 36234 580294 36290 580350
rect 36358 580294 36414 580350
rect 36482 580294 36538 580350
rect 36606 580294 36662 580350
rect 36234 580170 36290 580226
rect 36358 580170 36414 580226
rect 36482 580170 36538 580226
rect 36606 580170 36662 580226
rect 36234 580046 36290 580102
rect 36358 580046 36414 580102
rect 36482 580046 36538 580102
rect 36606 580046 36662 580102
rect 36234 579922 36290 579978
rect 36358 579922 36414 579978
rect 36482 579922 36538 579978
rect 36606 579922 36662 579978
rect 24518 562294 24574 562350
rect 24642 562294 24698 562350
rect 24518 562170 24574 562226
rect 24642 562170 24698 562226
rect 24518 562046 24574 562102
rect 24642 562046 24698 562102
rect 24518 561922 24574 561978
rect 24642 561922 24698 561978
rect 39954 598116 40010 598172
rect 40078 598116 40134 598172
rect 40202 598116 40258 598172
rect 40326 598116 40382 598172
rect 39954 597992 40010 598048
rect 40078 597992 40134 598048
rect 40202 597992 40258 598048
rect 40326 597992 40382 598048
rect 39954 597868 40010 597924
rect 40078 597868 40134 597924
rect 40202 597868 40258 597924
rect 40326 597868 40382 597924
rect 39954 597744 40010 597800
rect 40078 597744 40134 597800
rect 40202 597744 40258 597800
rect 40326 597744 40382 597800
rect 39954 586294 40010 586350
rect 40078 586294 40134 586350
rect 40202 586294 40258 586350
rect 40326 586294 40382 586350
rect 39954 586170 40010 586226
rect 40078 586170 40134 586226
rect 40202 586170 40258 586226
rect 40326 586170 40382 586226
rect 39954 586046 40010 586102
rect 40078 586046 40134 586102
rect 40202 586046 40258 586102
rect 40326 586046 40382 586102
rect 39954 585922 40010 585978
rect 40078 585922 40134 585978
rect 40202 585922 40258 585978
rect 40326 585922 40382 585978
rect 39954 568351 40010 568407
rect 40078 568351 40134 568407
rect 40202 568351 40258 568407
rect 40326 568351 40382 568407
rect 39954 568227 40010 568283
rect 40078 568227 40134 568283
rect 40202 568227 40258 568283
rect 40326 568227 40382 568283
rect 66954 597156 67010 597212
rect 67078 597156 67134 597212
rect 67202 597156 67258 597212
rect 67326 597156 67382 597212
rect 66954 597032 67010 597088
rect 67078 597032 67134 597088
rect 67202 597032 67258 597088
rect 67326 597032 67382 597088
rect 66954 596908 67010 596964
rect 67078 596908 67134 596964
rect 67202 596908 67258 596964
rect 67326 596908 67382 596964
rect 66954 596784 67010 596840
rect 67078 596784 67134 596840
rect 67202 596784 67258 596840
rect 67326 596784 67382 596840
rect 66954 580294 67010 580350
rect 67078 580294 67134 580350
rect 67202 580294 67258 580350
rect 67326 580294 67382 580350
rect 66954 580170 67010 580226
rect 67078 580170 67134 580226
rect 67202 580170 67258 580226
rect 67326 580170 67382 580226
rect 66954 580046 67010 580102
rect 67078 580046 67134 580102
rect 67202 580046 67258 580102
rect 67326 580046 67382 580102
rect 66954 579922 67010 579978
rect 67078 579922 67134 579978
rect 67202 579922 67258 579978
rect 67326 579922 67382 579978
rect 36234 562294 36290 562350
rect 36358 562294 36414 562350
rect 36482 562294 36538 562350
rect 36606 562294 36662 562350
rect 36234 562170 36290 562226
rect 36358 562170 36414 562226
rect 36482 562170 36538 562226
rect 36606 562170 36662 562226
rect 36234 562046 36290 562102
rect 36358 562046 36414 562102
rect 36482 562046 36538 562102
rect 36606 562046 36662 562102
rect 36234 561922 36290 561978
rect 36358 561922 36414 561978
rect 36482 561922 36538 561978
rect 36606 561922 36662 561978
rect 18396 554484 18452 554518
rect 18396 554462 18452 554484
rect 9234 550294 9290 550350
rect 9358 550294 9414 550350
rect 9482 550294 9538 550350
rect 9606 550294 9662 550350
rect 9234 550170 9290 550226
rect 9358 550170 9414 550226
rect 9482 550170 9538 550226
rect 9606 550170 9662 550226
rect 9234 550046 9290 550102
rect 9358 550046 9414 550102
rect 9482 550046 9538 550102
rect 9606 550046 9662 550102
rect 9234 549922 9290 549978
rect 9358 549922 9414 549978
rect 9482 549922 9538 549978
rect 9606 549922 9662 549978
rect 9234 532294 9290 532350
rect 9358 532294 9414 532350
rect 9482 532294 9538 532350
rect 9606 532294 9662 532350
rect 9234 532170 9290 532226
rect 9358 532170 9414 532226
rect 9482 532170 9538 532226
rect 9606 532170 9662 532226
rect 9234 532046 9290 532102
rect 9358 532046 9414 532102
rect 9482 532046 9538 532102
rect 9606 532046 9662 532102
rect 9234 531922 9290 531978
rect 9358 531922 9414 531978
rect 9482 531922 9538 531978
rect 9606 531922 9662 531978
rect 9234 514294 9290 514350
rect 9358 514294 9414 514350
rect 9482 514294 9538 514350
rect 9606 514294 9662 514350
rect 9234 514170 9290 514226
rect 9358 514170 9414 514226
rect 9482 514170 9538 514226
rect 9606 514170 9662 514226
rect 9234 514046 9290 514102
rect 9358 514046 9414 514102
rect 9482 514046 9538 514102
rect 9606 514046 9662 514102
rect 9234 513922 9290 513978
rect 9358 513922 9414 513978
rect 9482 513922 9538 513978
rect 9606 513922 9662 513978
rect 24518 544294 24574 544350
rect 24642 544294 24698 544350
rect 24518 544170 24574 544226
rect 24642 544170 24698 544226
rect 24518 544046 24574 544102
rect 24642 544046 24698 544102
rect 24518 543922 24574 543978
rect 24642 543922 24698 543978
rect 55238 562294 55294 562350
rect 55362 562294 55418 562350
rect 55238 562170 55294 562226
rect 55362 562170 55418 562226
rect 55238 562046 55294 562102
rect 55362 562046 55418 562102
rect 55238 561922 55294 561978
rect 55362 561922 55418 561978
rect 66954 562294 67010 562350
rect 67078 562294 67134 562350
rect 67202 562294 67258 562350
rect 67326 562294 67382 562350
rect 66954 562170 67010 562226
rect 67078 562170 67134 562226
rect 67202 562170 67258 562226
rect 67326 562170 67382 562226
rect 66954 562046 67010 562102
rect 67078 562046 67134 562102
rect 67202 562046 67258 562102
rect 67326 562046 67382 562102
rect 66954 561922 67010 561978
rect 67078 561922 67134 561978
rect 67202 561922 67258 561978
rect 67326 561922 67382 561978
rect 39878 550294 39934 550350
rect 40002 550294 40058 550350
rect 39878 550170 39934 550226
rect 40002 550170 40058 550226
rect 39878 550046 39934 550102
rect 40002 550046 40058 550102
rect 39878 549922 39934 549978
rect 40002 549922 40058 549978
rect 36234 544294 36290 544350
rect 36358 544294 36414 544350
rect 36482 544294 36538 544350
rect 36606 544294 36662 544350
rect 36234 544170 36290 544226
rect 36358 544170 36414 544226
rect 36482 544170 36538 544226
rect 36606 544170 36662 544226
rect 36234 544046 36290 544102
rect 36358 544046 36414 544102
rect 36482 544046 36538 544102
rect 36606 544046 36662 544102
rect 36234 543922 36290 543978
rect 36358 543922 36414 543978
rect 36482 543922 36538 543978
rect 36606 543922 36662 543978
rect 55238 544294 55294 544350
rect 55362 544294 55418 544350
rect 55238 544170 55294 544226
rect 55362 544170 55418 544226
rect 55238 544046 55294 544102
rect 55362 544046 55418 544102
rect 55238 543922 55294 543978
rect 55362 543922 55418 543978
rect 39878 532294 39934 532350
rect 40002 532294 40058 532350
rect 39878 532170 39934 532226
rect 40002 532170 40058 532226
rect 39878 532046 39934 532102
rect 40002 532046 40058 532102
rect 39878 531922 39934 531978
rect 40002 531922 40058 531978
rect 36234 526294 36290 526350
rect 36358 526294 36414 526350
rect 36482 526294 36538 526350
rect 36606 526294 36662 526350
rect 36234 526170 36290 526226
rect 36358 526170 36414 526226
rect 36482 526170 36538 526226
rect 36606 526170 36662 526226
rect 36234 526046 36290 526102
rect 36358 526046 36414 526102
rect 36482 526046 36538 526102
rect 36606 526046 36662 526102
rect 36234 525922 36290 525978
rect 36358 525922 36414 525978
rect 36482 525922 36538 525978
rect 36606 525922 36662 525978
rect 36234 508294 36290 508350
rect 36358 508294 36414 508350
rect 36482 508294 36538 508350
rect 36606 508294 36662 508350
rect 36234 508170 36290 508226
rect 36358 508170 36414 508226
rect 36482 508170 36538 508226
rect 36606 508170 36662 508226
rect 36234 508046 36290 508102
rect 36358 508046 36414 508102
rect 36482 508046 36538 508102
rect 36606 508046 36662 508102
rect 36234 507922 36290 507978
rect 36358 507922 36414 507978
rect 36482 507922 36538 507978
rect 36606 507922 36662 507978
rect 9234 496294 9290 496350
rect 9358 496294 9414 496350
rect 9482 496294 9538 496350
rect 9606 496294 9662 496350
rect 9234 496170 9290 496226
rect 9358 496170 9414 496226
rect 9482 496170 9538 496226
rect 9606 496170 9662 496226
rect 9234 496046 9290 496102
rect 9358 496046 9414 496102
rect 9482 496046 9538 496102
rect 9606 496046 9662 496102
rect 9234 495922 9290 495978
rect 9358 495922 9414 495978
rect 9482 495922 9538 495978
rect 9606 495922 9662 495978
rect 24518 490294 24574 490350
rect 24642 490294 24698 490350
rect 24518 490170 24574 490226
rect 24642 490170 24698 490226
rect 24518 490046 24574 490102
rect 24642 490046 24698 490102
rect 24518 489922 24574 489978
rect 24642 489922 24698 489978
rect 66954 544294 67010 544350
rect 67078 544294 67134 544350
rect 67202 544294 67258 544350
rect 67326 544294 67382 544350
rect 66954 544170 67010 544226
rect 67078 544170 67134 544226
rect 67202 544170 67258 544226
rect 67326 544170 67382 544226
rect 66954 544046 67010 544102
rect 67078 544046 67134 544102
rect 67202 544046 67258 544102
rect 67326 544046 67382 544102
rect 66954 543922 67010 543978
rect 67078 543922 67134 543978
rect 67202 543922 67258 543978
rect 67326 543922 67382 543978
rect 66954 526294 67010 526350
rect 67078 526294 67134 526350
rect 67202 526294 67258 526350
rect 67326 526294 67382 526350
rect 66954 526170 67010 526226
rect 67078 526170 67134 526226
rect 67202 526170 67258 526226
rect 67326 526170 67382 526226
rect 66954 526046 67010 526102
rect 67078 526046 67134 526102
rect 67202 526046 67258 526102
rect 67326 526046 67382 526102
rect 66954 525922 67010 525978
rect 67078 525922 67134 525978
rect 67202 525922 67258 525978
rect 67326 525922 67382 525978
rect 66954 508294 67010 508350
rect 67078 508294 67134 508350
rect 67202 508294 67258 508350
rect 67326 508294 67382 508350
rect 66954 508170 67010 508226
rect 67078 508170 67134 508226
rect 67202 508170 67258 508226
rect 67326 508170 67382 508226
rect 66954 508046 67010 508102
rect 67078 508046 67134 508102
rect 67202 508046 67258 508102
rect 67326 508046 67382 508102
rect 66954 507922 67010 507978
rect 67078 507922 67134 507978
rect 67202 507922 67258 507978
rect 67326 507922 67382 507978
rect 36234 490294 36290 490350
rect 36358 490294 36414 490350
rect 36482 490294 36538 490350
rect 36606 490294 36662 490350
rect 36234 490170 36290 490226
rect 36358 490170 36414 490226
rect 36482 490170 36538 490226
rect 36606 490170 36662 490226
rect 36234 490046 36290 490102
rect 36358 490046 36414 490102
rect 36482 490046 36538 490102
rect 36606 490046 36662 490102
rect 36234 489922 36290 489978
rect 36358 489922 36414 489978
rect 36482 489922 36538 489978
rect 36606 489922 36662 489978
rect 9234 478294 9290 478350
rect 9358 478294 9414 478350
rect 9482 478294 9538 478350
rect 9606 478294 9662 478350
rect 9234 478170 9290 478226
rect 9358 478170 9414 478226
rect 9482 478170 9538 478226
rect 9606 478170 9662 478226
rect 9234 478046 9290 478102
rect 9358 478046 9414 478102
rect 9482 478046 9538 478102
rect 9606 478046 9662 478102
rect 9234 477922 9290 477978
rect 9358 477922 9414 477978
rect 9482 477922 9538 477978
rect 9606 477922 9662 477978
rect 9234 460294 9290 460350
rect 9358 460294 9414 460350
rect 9482 460294 9538 460350
rect 9606 460294 9662 460350
rect 9234 460170 9290 460226
rect 9358 460170 9414 460226
rect 9482 460170 9538 460226
rect 9606 460170 9662 460226
rect 9234 460046 9290 460102
rect 9358 460046 9414 460102
rect 9482 460046 9538 460102
rect 9606 460046 9662 460102
rect 9234 459922 9290 459978
rect 9358 459922 9414 459978
rect 9482 459922 9538 459978
rect 9606 459922 9662 459978
rect 9234 442294 9290 442350
rect 9358 442294 9414 442350
rect 9482 442294 9538 442350
rect 9606 442294 9662 442350
rect 9234 442170 9290 442226
rect 9358 442170 9414 442226
rect 9482 442170 9538 442226
rect 9606 442170 9662 442226
rect 9234 442046 9290 442102
rect 9358 442046 9414 442102
rect 9482 442046 9538 442102
rect 9606 442046 9662 442102
rect 9234 441922 9290 441978
rect 9358 441922 9414 441978
rect 9482 441922 9538 441978
rect 9606 441922 9662 441978
rect 9234 424294 9290 424350
rect 9358 424294 9414 424350
rect 9482 424294 9538 424350
rect 9606 424294 9662 424350
rect 9234 424170 9290 424226
rect 9358 424170 9414 424226
rect 9482 424170 9538 424226
rect 9606 424170 9662 424226
rect 9234 424046 9290 424102
rect 9358 424046 9414 424102
rect 9482 424046 9538 424102
rect 9606 424046 9662 424102
rect 9234 423922 9290 423978
rect 9358 423922 9414 423978
rect 9482 423922 9538 423978
rect 9606 423922 9662 423978
rect 20076 482822 20132 482878
rect 24518 472294 24574 472350
rect 24642 472294 24698 472350
rect 24518 472170 24574 472226
rect 24642 472170 24698 472226
rect 24518 472046 24574 472102
rect 24642 472046 24698 472102
rect 24518 471922 24574 471978
rect 24642 471922 24698 471978
rect 55238 490294 55294 490350
rect 55362 490294 55418 490350
rect 55238 490170 55294 490226
rect 55362 490170 55418 490226
rect 55238 490046 55294 490102
rect 55362 490046 55418 490102
rect 55238 489922 55294 489978
rect 55362 489922 55418 489978
rect 70674 598116 70730 598172
rect 70798 598116 70854 598172
rect 70922 598116 70978 598172
rect 71046 598116 71102 598172
rect 70674 597992 70730 598048
rect 70798 597992 70854 598048
rect 70922 597992 70978 598048
rect 71046 597992 71102 598048
rect 70674 597868 70730 597924
rect 70798 597868 70854 597924
rect 70922 597868 70978 597924
rect 71046 597868 71102 597924
rect 70674 597744 70730 597800
rect 70798 597744 70854 597800
rect 70922 597744 70978 597800
rect 71046 597744 71102 597800
rect 70674 586294 70730 586350
rect 70798 586294 70854 586350
rect 70922 586294 70978 586350
rect 71046 586294 71102 586350
rect 70674 586170 70730 586226
rect 70798 586170 70854 586226
rect 70922 586170 70978 586226
rect 71046 586170 71102 586226
rect 70674 586046 70730 586102
rect 70798 586046 70854 586102
rect 70922 586046 70978 586102
rect 71046 586046 71102 586102
rect 70674 585922 70730 585978
rect 70798 585922 70854 585978
rect 70922 585922 70978 585978
rect 71046 585922 71102 585978
rect 70674 568294 70730 568350
rect 70798 568294 70854 568350
rect 70922 568294 70978 568350
rect 71046 568294 71102 568350
rect 70674 568170 70730 568226
rect 70798 568170 70854 568226
rect 70922 568170 70978 568226
rect 71046 568170 71102 568226
rect 70674 568046 70730 568102
rect 70798 568046 70854 568102
rect 70922 568046 70978 568102
rect 71046 568046 71102 568102
rect 70674 567922 70730 567978
rect 70798 567922 70854 567978
rect 70922 567922 70978 567978
rect 71046 567922 71102 567978
rect 97674 597156 97730 597212
rect 97798 597156 97854 597212
rect 97922 597156 97978 597212
rect 98046 597156 98102 597212
rect 97674 597032 97730 597088
rect 97798 597032 97854 597088
rect 97922 597032 97978 597088
rect 98046 597032 98102 597088
rect 97674 596908 97730 596964
rect 97798 596908 97854 596964
rect 97922 596908 97978 596964
rect 98046 596908 98102 596964
rect 97674 596784 97730 596840
rect 97798 596784 97854 596840
rect 97922 596784 97978 596840
rect 98046 596784 98102 596840
rect 97674 580294 97730 580350
rect 97798 580294 97854 580350
rect 97922 580294 97978 580350
rect 98046 580294 98102 580350
rect 97674 580170 97730 580226
rect 97798 580170 97854 580226
rect 97922 580170 97978 580226
rect 98046 580170 98102 580226
rect 97674 580046 97730 580102
rect 97798 580046 97854 580102
rect 97922 580046 97978 580102
rect 98046 580046 98102 580102
rect 97674 579922 97730 579978
rect 97798 579922 97854 579978
rect 97922 579922 97978 579978
rect 98046 579922 98102 579978
rect 86518 562294 86574 562350
rect 86642 562294 86698 562350
rect 86518 562170 86574 562226
rect 86642 562170 86698 562226
rect 86518 562046 86574 562102
rect 86642 562046 86698 562102
rect 86518 561922 86574 561978
rect 86642 561922 86698 561978
rect 101394 598116 101450 598172
rect 101518 598116 101574 598172
rect 101642 598116 101698 598172
rect 101766 598116 101822 598172
rect 101394 597992 101450 598048
rect 101518 597992 101574 598048
rect 101642 597992 101698 598048
rect 101766 597992 101822 598048
rect 101394 597868 101450 597924
rect 101518 597868 101574 597924
rect 101642 597868 101698 597924
rect 101766 597868 101822 597924
rect 101394 597744 101450 597800
rect 101518 597744 101574 597800
rect 101642 597744 101698 597800
rect 101766 597744 101822 597800
rect 101394 586294 101450 586350
rect 101518 586294 101574 586350
rect 101642 586294 101698 586350
rect 101766 586294 101822 586350
rect 101394 586170 101450 586226
rect 101518 586170 101574 586226
rect 101642 586170 101698 586226
rect 101766 586170 101822 586226
rect 101394 586046 101450 586102
rect 101518 586046 101574 586102
rect 101642 586046 101698 586102
rect 101766 586046 101822 586102
rect 101394 585922 101450 585978
rect 101518 585922 101574 585978
rect 101642 585922 101698 585978
rect 101766 585922 101822 585978
rect 101394 568351 101450 568407
rect 101518 568351 101574 568407
rect 101642 568351 101698 568407
rect 101766 568351 101822 568407
rect 101394 568227 101450 568283
rect 101518 568227 101574 568283
rect 101642 568227 101698 568283
rect 101766 568227 101822 568283
rect 128394 597156 128450 597212
rect 128518 597156 128574 597212
rect 128642 597156 128698 597212
rect 128766 597156 128822 597212
rect 128394 597032 128450 597088
rect 128518 597032 128574 597088
rect 128642 597032 128698 597088
rect 128766 597032 128822 597088
rect 128394 596908 128450 596964
rect 128518 596908 128574 596964
rect 128642 596908 128698 596964
rect 128766 596908 128822 596964
rect 128394 596784 128450 596840
rect 128518 596784 128574 596840
rect 128642 596784 128698 596840
rect 128766 596784 128822 596840
rect 128394 580294 128450 580350
rect 128518 580294 128574 580350
rect 128642 580294 128698 580350
rect 128766 580294 128822 580350
rect 128394 580170 128450 580226
rect 128518 580170 128574 580226
rect 128642 580170 128698 580226
rect 128766 580170 128822 580226
rect 128394 580046 128450 580102
rect 128518 580046 128574 580102
rect 128642 580046 128698 580102
rect 128766 580046 128822 580102
rect 128394 579922 128450 579978
rect 128518 579922 128574 579978
rect 128642 579922 128698 579978
rect 128766 579922 128822 579978
rect 97674 562294 97730 562350
rect 97798 562294 97854 562350
rect 97922 562294 97978 562350
rect 98046 562294 98102 562350
rect 97674 562170 97730 562226
rect 97798 562170 97854 562226
rect 97922 562170 97978 562226
rect 98046 562170 98102 562226
rect 97674 562046 97730 562102
rect 97798 562046 97854 562102
rect 97922 562046 97978 562102
rect 98046 562046 98102 562102
rect 97674 561922 97730 561978
rect 97798 561922 97854 561978
rect 97922 561922 97978 561978
rect 98046 561922 98102 561978
rect 70674 550294 70730 550350
rect 70798 550294 70854 550350
rect 70922 550294 70978 550350
rect 71046 550294 71102 550350
rect 70674 550170 70730 550226
rect 70798 550170 70854 550226
rect 70922 550170 70978 550226
rect 71046 550170 71102 550226
rect 70674 550046 70730 550102
rect 70798 550046 70854 550102
rect 70922 550046 70978 550102
rect 71046 550046 71102 550102
rect 70674 549922 70730 549978
rect 70798 549922 70854 549978
rect 70922 549922 70978 549978
rect 71046 549922 71102 549978
rect 70674 532294 70730 532350
rect 70798 532294 70854 532350
rect 70922 532294 70978 532350
rect 71046 532294 71102 532350
rect 70674 532170 70730 532226
rect 70798 532170 70854 532226
rect 70922 532170 70978 532226
rect 71046 532170 71102 532226
rect 70674 532046 70730 532102
rect 70798 532046 70854 532102
rect 70922 532046 70978 532102
rect 71046 532046 71102 532102
rect 70674 531922 70730 531978
rect 70798 531922 70854 531978
rect 70922 531922 70978 531978
rect 71046 531922 71102 531978
rect 70674 514294 70730 514350
rect 70798 514294 70854 514350
rect 70922 514294 70978 514350
rect 71046 514294 71102 514350
rect 70674 514170 70730 514226
rect 70798 514170 70854 514226
rect 70922 514170 70978 514226
rect 71046 514170 71102 514226
rect 70674 514046 70730 514102
rect 70798 514046 70854 514102
rect 70922 514046 70978 514102
rect 71046 514046 71102 514102
rect 70674 513922 70730 513978
rect 70798 513922 70854 513978
rect 70922 513922 70978 513978
rect 71046 513922 71102 513978
rect 82684 554462 82740 554518
rect 86518 544294 86574 544350
rect 86642 544294 86698 544350
rect 86518 544170 86574 544226
rect 86642 544170 86698 544226
rect 86518 544046 86574 544102
rect 86642 544046 86698 544102
rect 86518 543922 86574 543978
rect 86642 543922 86698 543978
rect 117238 562294 117294 562350
rect 117362 562294 117418 562350
rect 117238 562170 117294 562226
rect 117362 562170 117418 562226
rect 117238 562046 117294 562102
rect 117362 562046 117418 562102
rect 117238 561922 117294 561978
rect 117362 561922 117418 561978
rect 128394 562294 128450 562350
rect 128518 562294 128574 562350
rect 128642 562294 128698 562350
rect 128766 562294 128822 562350
rect 128394 562170 128450 562226
rect 128518 562170 128574 562226
rect 128642 562170 128698 562226
rect 128766 562170 128822 562226
rect 128394 562046 128450 562102
rect 128518 562046 128574 562102
rect 128642 562046 128698 562102
rect 128766 562046 128822 562102
rect 128394 561922 128450 561978
rect 128518 561922 128574 561978
rect 128642 561922 128698 561978
rect 128766 561922 128822 561978
rect 101878 550294 101934 550350
rect 102002 550294 102058 550350
rect 101878 550170 101934 550226
rect 102002 550170 102058 550226
rect 101878 550046 101934 550102
rect 102002 550046 102058 550102
rect 101878 549922 101934 549978
rect 102002 549922 102058 549978
rect 97674 544294 97730 544350
rect 97798 544294 97854 544350
rect 97922 544294 97978 544350
rect 98046 544294 98102 544350
rect 97674 544170 97730 544226
rect 97798 544170 97854 544226
rect 97922 544170 97978 544226
rect 98046 544170 98102 544226
rect 97674 544046 97730 544102
rect 97798 544046 97854 544102
rect 97922 544046 97978 544102
rect 98046 544046 98102 544102
rect 97674 543922 97730 543978
rect 97798 543922 97854 543978
rect 97922 543922 97978 543978
rect 98046 543922 98102 543978
rect 117238 544294 117294 544350
rect 117362 544294 117418 544350
rect 117238 544170 117294 544226
rect 117362 544170 117418 544226
rect 117238 544046 117294 544102
rect 117362 544046 117418 544102
rect 117238 543922 117294 543978
rect 117362 543922 117418 543978
rect 101878 532294 101934 532350
rect 102002 532294 102058 532350
rect 101878 532170 101934 532226
rect 102002 532170 102058 532226
rect 101878 532046 101934 532102
rect 102002 532046 102058 532102
rect 101878 531922 101934 531978
rect 102002 531922 102058 531978
rect 97674 526294 97730 526350
rect 97798 526294 97854 526350
rect 97922 526294 97978 526350
rect 98046 526294 98102 526350
rect 97674 526170 97730 526226
rect 97798 526170 97854 526226
rect 97922 526170 97978 526226
rect 98046 526170 98102 526226
rect 97674 526046 97730 526102
rect 97798 526046 97854 526102
rect 97922 526046 97978 526102
rect 98046 526046 98102 526102
rect 97674 525922 97730 525978
rect 97798 525922 97854 525978
rect 97922 525922 97978 525978
rect 98046 525922 98102 525978
rect 128394 544294 128450 544350
rect 128518 544294 128574 544350
rect 128642 544294 128698 544350
rect 128766 544294 128822 544350
rect 128394 544170 128450 544226
rect 128518 544170 128574 544226
rect 128642 544170 128698 544226
rect 128766 544170 128822 544226
rect 128394 544046 128450 544102
rect 128518 544046 128574 544102
rect 128642 544046 128698 544102
rect 128766 544046 128822 544102
rect 128394 543922 128450 543978
rect 128518 543922 128574 543978
rect 128642 543922 128698 543978
rect 128766 543922 128822 543978
rect 128394 526294 128450 526350
rect 128518 526294 128574 526350
rect 128642 526294 128698 526350
rect 128766 526294 128822 526350
rect 128394 526170 128450 526226
rect 128518 526170 128574 526226
rect 128642 526170 128698 526226
rect 128766 526170 128822 526226
rect 128394 526046 128450 526102
rect 128518 526046 128574 526102
rect 128642 526046 128698 526102
rect 128766 526046 128822 526102
rect 128394 525922 128450 525978
rect 128518 525922 128574 525978
rect 128642 525922 128698 525978
rect 128766 525922 128822 525978
rect 97674 508294 97730 508350
rect 97798 508294 97854 508350
rect 97922 508294 97978 508350
rect 98046 508294 98102 508350
rect 97674 508170 97730 508226
rect 97798 508170 97854 508226
rect 97922 508170 97978 508226
rect 98046 508170 98102 508226
rect 97674 508046 97730 508102
rect 97798 508046 97854 508102
rect 97922 508046 97978 508102
rect 98046 508046 98102 508102
rect 97674 507922 97730 507978
rect 97798 507922 97854 507978
rect 97922 507922 97978 507978
rect 98046 507922 98102 507978
rect 70674 496294 70730 496350
rect 70798 496294 70854 496350
rect 70922 496294 70978 496350
rect 71046 496294 71102 496350
rect 70674 496170 70730 496226
rect 70798 496170 70854 496226
rect 70922 496170 70978 496226
rect 71046 496170 71102 496226
rect 70674 496046 70730 496102
rect 70798 496046 70854 496102
rect 70922 496046 70978 496102
rect 71046 496046 71102 496102
rect 70674 495922 70730 495978
rect 70798 495922 70854 495978
rect 70922 495922 70978 495978
rect 71046 495922 71102 495978
rect 66954 490294 67010 490350
rect 67078 490294 67134 490350
rect 67202 490294 67258 490350
rect 67326 490294 67382 490350
rect 66954 490170 67010 490226
rect 67078 490170 67134 490226
rect 67202 490170 67258 490226
rect 67326 490170 67382 490226
rect 66954 490046 67010 490102
rect 67078 490046 67134 490102
rect 67202 490046 67258 490102
rect 67326 490046 67382 490102
rect 66954 489922 67010 489978
rect 67078 489922 67134 489978
rect 67202 489922 67258 489978
rect 67326 489922 67382 489978
rect 39878 478294 39934 478350
rect 40002 478294 40058 478350
rect 39878 478170 39934 478226
rect 40002 478170 40058 478226
rect 39878 478046 39934 478102
rect 40002 478046 40058 478102
rect 39878 477922 39934 477978
rect 40002 477922 40058 477978
rect 36234 472294 36290 472350
rect 36358 472294 36414 472350
rect 36482 472294 36538 472350
rect 36606 472294 36662 472350
rect 36234 472170 36290 472226
rect 36358 472170 36414 472226
rect 36482 472170 36538 472226
rect 36606 472170 36662 472226
rect 36234 472046 36290 472102
rect 36358 472046 36414 472102
rect 36482 472046 36538 472102
rect 36606 472046 36662 472102
rect 36234 471922 36290 471978
rect 36358 471922 36414 471978
rect 36482 471922 36538 471978
rect 36606 471922 36662 471978
rect 55238 472294 55294 472350
rect 55362 472294 55418 472350
rect 55238 472170 55294 472226
rect 55362 472170 55418 472226
rect 55238 472046 55294 472102
rect 55362 472046 55418 472102
rect 55238 471922 55294 471978
rect 55362 471922 55418 471978
rect 39878 460294 39934 460350
rect 40002 460294 40058 460350
rect 39878 460170 39934 460226
rect 40002 460170 40058 460226
rect 39878 460046 39934 460102
rect 40002 460046 40058 460102
rect 39878 459922 39934 459978
rect 40002 459922 40058 459978
rect 36234 454294 36290 454350
rect 36358 454294 36414 454350
rect 36482 454294 36538 454350
rect 36606 454294 36662 454350
rect 36234 454170 36290 454226
rect 36358 454170 36414 454226
rect 36482 454170 36538 454226
rect 36606 454170 36662 454226
rect 36234 454046 36290 454102
rect 36358 454046 36414 454102
rect 36482 454046 36538 454102
rect 36606 454046 36662 454102
rect 36234 453922 36290 453978
rect 36358 453922 36414 453978
rect 36482 453922 36538 453978
rect 36606 453922 36662 453978
rect 66954 472294 67010 472350
rect 67078 472294 67134 472350
rect 67202 472294 67258 472350
rect 67326 472294 67382 472350
rect 66954 472170 67010 472226
rect 67078 472170 67134 472226
rect 67202 472170 67258 472226
rect 67326 472170 67382 472226
rect 66954 472046 67010 472102
rect 67078 472046 67134 472102
rect 67202 472046 67258 472102
rect 67326 472046 67382 472102
rect 66954 471922 67010 471978
rect 67078 471922 67134 471978
rect 67202 471922 67258 471978
rect 67326 471922 67382 471978
rect 86518 490294 86574 490350
rect 86642 490294 86698 490350
rect 86518 490170 86574 490226
rect 86642 490170 86698 490226
rect 86518 490046 86574 490102
rect 86642 490046 86698 490102
rect 86518 489922 86574 489978
rect 86642 489922 86698 489978
rect 128394 508294 128450 508350
rect 128518 508294 128574 508350
rect 128642 508294 128698 508350
rect 128766 508294 128822 508350
rect 128394 508170 128450 508226
rect 128518 508170 128574 508226
rect 128642 508170 128698 508226
rect 128766 508170 128822 508226
rect 128394 508046 128450 508102
rect 128518 508046 128574 508102
rect 128642 508046 128698 508102
rect 128766 508046 128822 508102
rect 128394 507922 128450 507978
rect 128518 507922 128574 507978
rect 128642 507922 128698 507978
rect 128766 507922 128822 507978
rect 97674 490294 97730 490350
rect 97798 490294 97854 490350
rect 97922 490294 97978 490350
rect 98046 490294 98102 490350
rect 97674 490170 97730 490226
rect 97798 490170 97854 490226
rect 97922 490170 97978 490226
rect 98046 490170 98102 490226
rect 97674 490046 97730 490102
rect 97798 490046 97854 490102
rect 97922 490046 97978 490102
rect 98046 490046 98102 490102
rect 97674 489922 97730 489978
rect 97798 489922 97854 489978
rect 97922 489922 97978 489978
rect 98046 489922 98102 489978
rect 82684 483002 82740 483058
rect 70674 478294 70730 478350
rect 70798 478294 70854 478350
rect 70922 478294 70978 478350
rect 71046 478294 71102 478350
rect 70674 478170 70730 478226
rect 70798 478170 70854 478226
rect 70922 478170 70978 478226
rect 71046 478170 71102 478226
rect 70674 478046 70730 478102
rect 70798 478046 70854 478102
rect 70922 478046 70978 478102
rect 71046 478046 71102 478102
rect 70674 477922 70730 477978
rect 70798 477922 70854 477978
rect 70922 477922 70978 477978
rect 71046 477922 71102 477978
rect 66954 454294 67010 454350
rect 67078 454294 67134 454350
rect 67202 454294 67258 454350
rect 67326 454294 67382 454350
rect 66954 454170 67010 454226
rect 67078 454170 67134 454226
rect 67202 454170 67258 454226
rect 67326 454170 67382 454226
rect 66954 454046 67010 454102
rect 67078 454046 67134 454102
rect 67202 454046 67258 454102
rect 67326 454046 67382 454102
rect 66954 453922 67010 453978
rect 67078 453922 67134 453978
rect 67202 453922 67258 453978
rect 67326 453922 67382 453978
rect 36234 436294 36290 436350
rect 36358 436294 36414 436350
rect 36482 436294 36538 436350
rect 36606 436294 36662 436350
rect 36234 436170 36290 436226
rect 36358 436170 36414 436226
rect 36482 436170 36538 436226
rect 36606 436170 36662 436226
rect 36234 436046 36290 436102
rect 36358 436046 36414 436102
rect 36482 436046 36538 436102
rect 36606 436046 36662 436102
rect 36234 435922 36290 435978
rect 36358 435922 36414 435978
rect 36482 435922 36538 435978
rect 36606 435922 36662 435978
rect 24518 418294 24574 418350
rect 24642 418294 24698 418350
rect 24518 418170 24574 418226
rect 24642 418170 24698 418226
rect 24518 418046 24574 418102
rect 24642 418046 24698 418102
rect 24518 417922 24574 417978
rect 24642 417922 24698 417978
rect 70674 460294 70730 460350
rect 70798 460294 70854 460350
rect 70922 460294 70978 460350
rect 71046 460294 71102 460350
rect 70674 460170 70730 460226
rect 70798 460170 70854 460226
rect 70922 460170 70978 460226
rect 71046 460170 71102 460226
rect 70674 460046 70730 460102
rect 70798 460046 70854 460102
rect 70922 460046 70978 460102
rect 71046 460046 71102 460102
rect 70674 459922 70730 459978
rect 70798 459922 70854 459978
rect 70922 459922 70978 459978
rect 71046 459922 71102 459978
rect 70674 442294 70730 442350
rect 70798 442294 70854 442350
rect 70922 442294 70978 442350
rect 71046 442294 71102 442350
rect 70674 442170 70730 442226
rect 70798 442170 70854 442226
rect 70922 442170 70978 442226
rect 71046 442170 71102 442226
rect 70674 442046 70730 442102
rect 70798 442046 70854 442102
rect 70922 442046 70978 442102
rect 71046 442046 71102 442102
rect 70674 441922 70730 441978
rect 70798 441922 70854 441978
rect 70922 441922 70978 441978
rect 71046 441922 71102 441978
rect 66954 436294 67010 436350
rect 67078 436294 67134 436350
rect 67202 436294 67258 436350
rect 67326 436294 67382 436350
rect 66954 436170 67010 436226
rect 67078 436170 67134 436226
rect 67202 436170 67258 436226
rect 67326 436170 67382 436226
rect 66954 436046 67010 436102
rect 67078 436046 67134 436102
rect 67202 436046 67258 436102
rect 67326 436046 67382 436102
rect 66954 435922 67010 435978
rect 67078 435922 67134 435978
rect 67202 435922 67258 435978
rect 67326 435922 67382 435978
rect 36234 418294 36290 418350
rect 36358 418294 36414 418350
rect 36482 418294 36538 418350
rect 36606 418294 36662 418350
rect 36234 418170 36290 418226
rect 36358 418170 36414 418226
rect 36482 418170 36538 418226
rect 36606 418170 36662 418226
rect 36234 418046 36290 418102
rect 36358 418046 36414 418102
rect 36482 418046 36538 418102
rect 36606 418046 36662 418102
rect 36234 417922 36290 417978
rect 36358 417922 36414 417978
rect 36482 417922 36538 417978
rect 36606 417922 36662 417978
rect 18396 413162 18452 413218
rect 9234 406294 9290 406350
rect 9358 406294 9414 406350
rect 9482 406294 9538 406350
rect 9606 406294 9662 406350
rect 9234 406170 9290 406226
rect 9358 406170 9414 406226
rect 9482 406170 9538 406226
rect 9606 406170 9662 406226
rect 9234 406046 9290 406102
rect 9358 406046 9414 406102
rect 9482 406046 9538 406102
rect 9606 406046 9662 406102
rect 9234 405922 9290 405978
rect 9358 405922 9414 405978
rect 9482 405922 9538 405978
rect 9606 405922 9662 405978
rect 9234 388294 9290 388350
rect 9358 388294 9414 388350
rect 9482 388294 9538 388350
rect 9606 388294 9662 388350
rect 9234 388170 9290 388226
rect 9358 388170 9414 388226
rect 9482 388170 9538 388226
rect 9606 388170 9662 388226
rect 9234 388046 9290 388102
rect 9358 388046 9414 388102
rect 9482 388046 9538 388102
rect 9606 388046 9662 388102
rect 9234 387922 9290 387978
rect 9358 387922 9414 387978
rect 9482 387922 9538 387978
rect 9606 387922 9662 387978
rect 9234 370294 9290 370350
rect 9358 370294 9414 370350
rect 9482 370294 9538 370350
rect 9606 370294 9662 370350
rect 9234 370170 9290 370226
rect 9358 370170 9414 370226
rect 9482 370170 9538 370226
rect 9606 370170 9662 370226
rect 9234 370046 9290 370102
rect 9358 370046 9414 370102
rect 9482 370046 9538 370102
rect 9606 370046 9662 370102
rect 9234 369922 9290 369978
rect 9358 369922 9414 369978
rect 9482 369922 9538 369978
rect 9606 369922 9662 369978
rect 20636 406700 20692 406738
rect 20636 406682 20692 406700
rect 24518 400294 24574 400350
rect 24642 400294 24698 400350
rect 24518 400170 24574 400226
rect 24642 400170 24698 400226
rect 24518 400046 24574 400102
rect 24642 400046 24698 400102
rect 24518 399922 24574 399978
rect 24642 399922 24698 399978
rect 55238 418294 55294 418350
rect 55362 418294 55418 418350
rect 55238 418170 55294 418226
rect 55362 418170 55418 418226
rect 55238 418046 55294 418102
rect 55362 418046 55418 418102
rect 55238 417922 55294 417978
rect 55362 417922 55418 417978
rect 66954 418294 67010 418350
rect 67078 418294 67134 418350
rect 67202 418294 67258 418350
rect 67326 418294 67382 418350
rect 66954 418170 67010 418226
rect 67078 418170 67134 418226
rect 67202 418170 67258 418226
rect 67326 418170 67382 418226
rect 66954 418046 67010 418102
rect 67078 418046 67134 418102
rect 67202 418046 67258 418102
rect 67326 418046 67382 418102
rect 66954 417922 67010 417978
rect 67078 417922 67134 417978
rect 67202 417922 67258 417978
rect 67326 417922 67382 417978
rect 62972 406682 63028 406738
rect 39878 406294 39934 406350
rect 40002 406294 40058 406350
rect 39878 406170 39934 406226
rect 40002 406170 40058 406226
rect 39878 406046 39934 406102
rect 40002 406046 40058 406102
rect 39878 405922 39934 405978
rect 40002 405922 40058 405978
rect 36234 400294 36290 400350
rect 36358 400294 36414 400350
rect 36482 400294 36538 400350
rect 36606 400294 36662 400350
rect 36234 400170 36290 400226
rect 36358 400170 36414 400226
rect 36482 400170 36538 400226
rect 36606 400170 36662 400226
rect 36234 400046 36290 400102
rect 36358 400046 36414 400102
rect 36482 400046 36538 400102
rect 36606 400046 36662 400102
rect 36234 399922 36290 399978
rect 36358 399922 36414 399978
rect 36482 399922 36538 399978
rect 36606 399922 36662 399978
rect 55238 400294 55294 400350
rect 55362 400294 55418 400350
rect 55238 400170 55294 400226
rect 55362 400170 55418 400226
rect 55238 400046 55294 400102
rect 55362 400046 55418 400102
rect 55238 399922 55294 399978
rect 55362 399922 55418 399978
rect 62972 391382 63028 391438
rect 39836 388333 39892 388389
rect 39940 388333 39996 388389
rect 40044 388333 40100 388389
rect 36234 382294 36290 382350
rect 36358 382294 36414 382350
rect 36482 382294 36538 382350
rect 36606 382294 36662 382350
rect 36234 382170 36290 382226
rect 36358 382170 36414 382226
rect 36482 382170 36538 382226
rect 36606 382170 36662 382226
rect 36234 382046 36290 382102
rect 36358 382046 36414 382102
rect 36482 382046 36538 382102
rect 36606 382046 36662 382102
rect 36234 381922 36290 381978
rect 36358 381922 36414 381978
rect 36482 381922 36538 381978
rect 36606 381922 36662 381978
rect 36234 364294 36290 364350
rect 36358 364294 36414 364350
rect 36482 364294 36538 364350
rect 36606 364294 36662 364350
rect 36234 364170 36290 364226
rect 36358 364170 36414 364226
rect 36482 364170 36538 364226
rect 36606 364170 36662 364226
rect 36234 364046 36290 364102
rect 36358 364046 36414 364102
rect 36482 364046 36538 364102
rect 36606 364046 36662 364102
rect 36234 363922 36290 363978
rect 36358 363922 36414 363978
rect 36482 363922 36538 363978
rect 36606 363922 36662 363978
rect 9234 352294 9290 352350
rect 9358 352294 9414 352350
rect 9482 352294 9538 352350
rect 9606 352294 9662 352350
rect 9234 352170 9290 352226
rect 9358 352170 9414 352226
rect 9482 352170 9538 352226
rect 9606 352170 9662 352226
rect 9234 352046 9290 352102
rect 9358 352046 9414 352102
rect 9482 352046 9538 352102
rect 9606 352046 9662 352102
rect 9234 351922 9290 351978
rect 9358 351922 9414 351978
rect 9482 351922 9538 351978
rect 9606 351922 9662 351978
rect 24518 346294 24574 346350
rect 24642 346294 24698 346350
rect 24518 346170 24574 346226
rect 24642 346170 24698 346226
rect 24518 346046 24574 346102
rect 24642 346046 24698 346102
rect 24518 345922 24574 345978
rect 24642 345922 24698 345978
rect 117238 490294 117294 490350
rect 117362 490294 117418 490350
rect 117238 490170 117294 490226
rect 117362 490170 117418 490226
rect 117238 490046 117294 490102
rect 117362 490046 117418 490102
rect 117238 489922 117294 489978
rect 117362 489922 117418 489978
rect 128394 490294 128450 490350
rect 128518 490294 128574 490350
rect 128642 490294 128698 490350
rect 128766 490294 128822 490350
rect 128394 490170 128450 490226
rect 128518 490170 128574 490226
rect 128642 490170 128698 490226
rect 128766 490170 128822 490226
rect 128394 490046 128450 490102
rect 128518 490046 128574 490102
rect 128642 490046 128698 490102
rect 128766 490046 128822 490102
rect 128394 489922 128450 489978
rect 128518 489922 128574 489978
rect 128642 489922 128698 489978
rect 128766 489922 128822 489978
rect 101878 478294 101934 478350
rect 102002 478294 102058 478350
rect 101878 478170 101934 478226
rect 102002 478170 102058 478226
rect 101878 478046 101934 478102
rect 102002 478046 102058 478102
rect 101878 477922 101934 477978
rect 102002 477922 102058 477978
rect 86518 472294 86574 472350
rect 86642 472294 86698 472350
rect 86518 472170 86574 472226
rect 86642 472170 86698 472226
rect 86518 472046 86574 472102
rect 86642 472046 86698 472102
rect 86518 471922 86574 471978
rect 86642 471922 86698 471978
rect 97674 472294 97730 472350
rect 97798 472294 97854 472350
rect 97922 472294 97978 472350
rect 98046 472294 98102 472350
rect 97674 472170 97730 472226
rect 97798 472170 97854 472226
rect 97922 472170 97978 472226
rect 98046 472170 98102 472226
rect 97674 472046 97730 472102
rect 97798 472046 97854 472102
rect 97922 472046 97978 472102
rect 98046 472046 98102 472102
rect 97674 471922 97730 471978
rect 97798 471922 97854 471978
rect 97922 471922 97978 471978
rect 98046 471922 98102 471978
rect 117238 472294 117294 472350
rect 117362 472294 117418 472350
rect 117238 472170 117294 472226
rect 117362 472170 117418 472226
rect 117238 472046 117294 472102
rect 117362 472046 117418 472102
rect 117238 471922 117294 471978
rect 117362 471922 117418 471978
rect 101878 460294 101934 460350
rect 102002 460294 102058 460350
rect 101878 460170 101934 460226
rect 102002 460170 102058 460226
rect 101878 460046 101934 460102
rect 102002 460046 102058 460102
rect 101878 459922 101934 459978
rect 102002 459922 102058 459978
rect 97674 454294 97730 454350
rect 97798 454294 97854 454350
rect 97922 454294 97978 454350
rect 98046 454294 98102 454350
rect 97674 454170 97730 454226
rect 97798 454170 97854 454226
rect 97922 454170 97978 454226
rect 98046 454170 98102 454226
rect 97674 454046 97730 454102
rect 97798 454046 97854 454102
rect 97922 454046 97978 454102
rect 98046 454046 98102 454102
rect 97674 453922 97730 453978
rect 97798 453922 97854 453978
rect 97922 453922 97978 453978
rect 98046 453922 98102 453978
rect 132114 598116 132170 598172
rect 132238 598116 132294 598172
rect 132362 598116 132418 598172
rect 132486 598116 132542 598172
rect 132114 597992 132170 598048
rect 132238 597992 132294 598048
rect 132362 597992 132418 598048
rect 132486 597992 132542 598048
rect 132114 597868 132170 597924
rect 132238 597868 132294 597924
rect 132362 597868 132418 597924
rect 132486 597868 132542 597924
rect 132114 597744 132170 597800
rect 132238 597744 132294 597800
rect 132362 597744 132418 597800
rect 132486 597744 132542 597800
rect 132114 586294 132170 586350
rect 132238 586294 132294 586350
rect 132362 586294 132418 586350
rect 132486 586294 132542 586350
rect 132114 586170 132170 586226
rect 132238 586170 132294 586226
rect 132362 586170 132418 586226
rect 132486 586170 132542 586226
rect 132114 586046 132170 586102
rect 132238 586046 132294 586102
rect 132362 586046 132418 586102
rect 132486 586046 132542 586102
rect 132114 585922 132170 585978
rect 132238 585922 132294 585978
rect 132362 585922 132418 585978
rect 132486 585922 132542 585978
rect 132114 568294 132170 568350
rect 132238 568294 132294 568350
rect 132362 568294 132418 568350
rect 132486 568294 132542 568350
rect 132114 568170 132170 568226
rect 132238 568170 132294 568226
rect 132362 568170 132418 568226
rect 132486 568170 132542 568226
rect 132114 568046 132170 568102
rect 132238 568046 132294 568102
rect 132362 568046 132418 568102
rect 132486 568046 132542 568102
rect 132114 567922 132170 567978
rect 132238 567922 132294 567978
rect 132362 567922 132418 567978
rect 132486 567922 132542 567978
rect 159114 597156 159170 597212
rect 159238 597156 159294 597212
rect 159362 597156 159418 597212
rect 159486 597156 159542 597212
rect 159114 597032 159170 597088
rect 159238 597032 159294 597088
rect 159362 597032 159418 597088
rect 159486 597032 159542 597088
rect 159114 596908 159170 596964
rect 159238 596908 159294 596964
rect 159362 596908 159418 596964
rect 159486 596908 159542 596964
rect 159114 596784 159170 596840
rect 159238 596784 159294 596840
rect 159362 596784 159418 596840
rect 159486 596784 159542 596840
rect 159114 580294 159170 580350
rect 159238 580294 159294 580350
rect 159362 580294 159418 580350
rect 159486 580294 159542 580350
rect 159114 580170 159170 580226
rect 159238 580170 159294 580226
rect 159362 580170 159418 580226
rect 159486 580170 159542 580226
rect 159114 580046 159170 580102
rect 159238 580046 159294 580102
rect 159362 580046 159418 580102
rect 159486 580046 159542 580102
rect 159114 579922 159170 579978
rect 159238 579922 159294 579978
rect 159362 579922 159418 579978
rect 159486 579922 159542 579978
rect 148518 562294 148574 562350
rect 148642 562294 148698 562350
rect 148518 562170 148574 562226
rect 148642 562170 148698 562226
rect 148518 562046 148574 562102
rect 148642 562046 148698 562102
rect 148518 561922 148574 561978
rect 148642 561922 148698 561978
rect 159114 562294 159170 562350
rect 159238 562294 159294 562350
rect 159362 562294 159418 562350
rect 159486 562294 159542 562350
rect 159114 562170 159170 562226
rect 159238 562170 159294 562226
rect 159362 562170 159418 562226
rect 159486 562170 159542 562226
rect 159114 562046 159170 562102
rect 159238 562046 159294 562102
rect 159362 562046 159418 562102
rect 159486 562046 159542 562102
rect 159114 561922 159170 561978
rect 159238 561922 159294 561978
rect 159362 561922 159418 561978
rect 159486 561922 159542 561978
rect 141036 554462 141092 554518
rect 132114 550294 132170 550350
rect 132238 550294 132294 550350
rect 132362 550294 132418 550350
rect 132486 550294 132542 550350
rect 132114 550170 132170 550226
rect 132238 550170 132294 550226
rect 132362 550170 132418 550226
rect 132486 550170 132542 550226
rect 132114 550046 132170 550102
rect 132238 550046 132294 550102
rect 132362 550046 132418 550102
rect 132486 550046 132542 550102
rect 132114 549922 132170 549978
rect 132238 549922 132294 549978
rect 132362 549922 132418 549978
rect 132486 549922 132542 549978
rect 132114 532294 132170 532350
rect 132238 532294 132294 532350
rect 132362 532294 132418 532350
rect 132486 532294 132542 532350
rect 132114 532170 132170 532226
rect 132238 532170 132294 532226
rect 132362 532170 132418 532226
rect 132486 532170 132542 532226
rect 132114 532046 132170 532102
rect 132238 532046 132294 532102
rect 132362 532046 132418 532102
rect 132486 532046 132542 532102
rect 132114 531922 132170 531978
rect 132238 531922 132294 531978
rect 132362 531922 132418 531978
rect 132486 531922 132542 531978
rect 132114 514294 132170 514350
rect 132238 514294 132294 514350
rect 132362 514294 132418 514350
rect 132486 514294 132542 514350
rect 132114 514170 132170 514226
rect 132238 514170 132294 514226
rect 132362 514170 132418 514226
rect 132486 514170 132542 514226
rect 132114 514046 132170 514102
rect 132238 514046 132294 514102
rect 132362 514046 132418 514102
rect 132486 514046 132542 514102
rect 132114 513922 132170 513978
rect 132238 513922 132294 513978
rect 132362 513922 132418 513978
rect 132486 513922 132542 513978
rect 144060 555212 144116 555238
rect 144060 555182 144116 555212
rect 148518 544294 148574 544350
rect 148642 544294 148698 544350
rect 148518 544170 148574 544226
rect 148642 544170 148698 544226
rect 148518 544046 148574 544102
rect 148642 544046 148698 544102
rect 148518 543922 148574 543978
rect 148642 543922 148698 543978
rect 162834 598116 162890 598172
rect 162958 598116 163014 598172
rect 163082 598116 163138 598172
rect 163206 598116 163262 598172
rect 162834 597992 162890 598048
rect 162958 597992 163014 598048
rect 163082 597992 163138 598048
rect 163206 597992 163262 598048
rect 162834 597868 162890 597924
rect 162958 597868 163014 597924
rect 163082 597868 163138 597924
rect 163206 597868 163262 597924
rect 162834 597744 162890 597800
rect 162958 597744 163014 597800
rect 163082 597744 163138 597800
rect 163206 597744 163262 597800
rect 162834 586294 162890 586350
rect 162958 586294 163014 586350
rect 163082 586294 163138 586350
rect 163206 586294 163262 586350
rect 162834 586170 162890 586226
rect 162958 586170 163014 586226
rect 163082 586170 163138 586226
rect 163206 586170 163262 586226
rect 162834 586046 162890 586102
rect 162958 586046 163014 586102
rect 163082 586046 163138 586102
rect 163206 586046 163262 586102
rect 162834 585922 162890 585978
rect 162958 585922 163014 585978
rect 163082 585922 163138 585978
rect 163206 585922 163262 585978
rect 162834 568294 162890 568350
rect 162958 568294 163014 568350
rect 163082 568294 163138 568350
rect 163206 568294 163262 568350
rect 162834 568170 162890 568226
rect 162958 568170 163014 568226
rect 163082 568170 163138 568226
rect 163206 568170 163262 568226
rect 162834 568046 162890 568102
rect 162958 568046 163014 568102
rect 163082 568046 163138 568102
rect 163206 568046 163262 568102
rect 162834 567922 162890 567978
rect 162958 567922 163014 567978
rect 163082 567922 163138 567978
rect 163206 567922 163262 567978
rect 189834 597156 189890 597212
rect 189958 597156 190014 597212
rect 190082 597156 190138 597212
rect 190206 597156 190262 597212
rect 189834 597032 189890 597088
rect 189958 597032 190014 597088
rect 190082 597032 190138 597088
rect 190206 597032 190262 597088
rect 189834 596908 189890 596964
rect 189958 596908 190014 596964
rect 190082 596908 190138 596964
rect 190206 596908 190262 596964
rect 189834 596784 189890 596840
rect 189958 596784 190014 596840
rect 190082 596784 190138 596840
rect 190206 596784 190262 596840
rect 189834 580294 189890 580350
rect 189958 580294 190014 580350
rect 190082 580294 190138 580350
rect 190206 580294 190262 580350
rect 189834 580170 189890 580226
rect 189958 580170 190014 580226
rect 190082 580170 190138 580226
rect 190206 580170 190262 580226
rect 189834 580046 189890 580102
rect 189958 580046 190014 580102
rect 190082 580046 190138 580102
rect 190206 580046 190262 580102
rect 189834 579922 189890 579978
rect 189958 579922 190014 579978
rect 190082 579922 190138 579978
rect 190206 579922 190262 579978
rect 179238 562294 179294 562350
rect 179362 562294 179418 562350
rect 179238 562170 179294 562226
rect 179362 562170 179418 562226
rect 179238 562046 179294 562102
rect 179362 562046 179418 562102
rect 179238 561922 179294 561978
rect 179362 561922 179418 561978
rect 189834 562294 189890 562350
rect 189958 562294 190014 562350
rect 190082 562294 190138 562350
rect 190206 562294 190262 562350
rect 189834 562170 189890 562226
rect 189958 562170 190014 562226
rect 190082 562170 190138 562226
rect 190206 562170 190262 562226
rect 189834 562046 189890 562102
rect 189958 562046 190014 562102
rect 190082 562046 190138 562102
rect 190206 562046 190262 562102
rect 189834 561922 189890 561978
rect 189958 561922 190014 561978
rect 190082 561922 190138 561978
rect 190206 561922 190262 561978
rect 163878 550294 163934 550350
rect 164002 550294 164058 550350
rect 163878 550170 163934 550226
rect 164002 550170 164058 550226
rect 163878 550046 163934 550102
rect 164002 550046 164058 550102
rect 163878 549922 163934 549978
rect 164002 549922 164058 549978
rect 159114 544294 159170 544350
rect 159238 544294 159294 544350
rect 159362 544294 159418 544350
rect 159486 544294 159542 544350
rect 159114 544170 159170 544226
rect 159238 544170 159294 544226
rect 159362 544170 159418 544226
rect 159486 544170 159542 544226
rect 159114 544046 159170 544102
rect 159238 544046 159294 544102
rect 159362 544046 159418 544102
rect 159486 544046 159542 544102
rect 159114 543922 159170 543978
rect 159238 543922 159294 543978
rect 159362 543922 159418 543978
rect 159486 543922 159542 543978
rect 179238 544294 179294 544350
rect 179362 544294 179418 544350
rect 179238 544170 179294 544226
rect 179362 544170 179418 544226
rect 179238 544046 179294 544102
rect 179362 544046 179418 544102
rect 179238 543922 179294 543978
rect 179362 543922 179418 543978
rect 159114 526294 159170 526350
rect 159238 526294 159294 526350
rect 159362 526294 159418 526350
rect 159486 526294 159542 526350
rect 159114 526170 159170 526226
rect 159238 526170 159294 526226
rect 159362 526170 159418 526226
rect 159486 526170 159542 526226
rect 159114 526046 159170 526102
rect 159238 526046 159294 526102
rect 159362 526046 159418 526102
rect 159486 526046 159542 526102
rect 159114 525922 159170 525978
rect 159238 525922 159294 525978
rect 159362 525922 159418 525978
rect 159486 525922 159542 525978
rect 132114 496294 132170 496350
rect 132238 496294 132294 496350
rect 132362 496294 132418 496350
rect 132486 496294 132542 496350
rect 132114 496170 132170 496226
rect 132238 496170 132294 496226
rect 132362 496170 132418 496226
rect 132486 496170 132542 496226
rect 132114 496046 132170 496102
rect 132238 496046 132294 496102
rect 132362 496046 132418 496102
rect 132486 496046 132542 496102
rect 132114 495922 132170 495978
rect 132238 495922 132294 495978
rect 132362 495922 132418 495978
rect 132486 495922 132542 495978
rect 128394 472294 128450 472350
rect 128518 472294 128574 472350
rect 128642 472294 128698 472350
rect 128766 472294 128822 472350
rect 128394 472170 128450 472226
rect 128518 472170 128574 472226
rect 128642 472170 128698 472226
rect 128766 472170 128822 472226
rect 128394 472046 128450 472102
rect 128518 472046 128574 472102
rect 128642 472046 128698 472102
rect 128766 472046 128822 472102
rect 128394 471922 128450 471978
rect 128518 471922 128574 471978
rect 128642 471922 128698 471978
rect 128766 471922 128822 471978
rect 159114 508294 159170 508350
rect 159238 508294 159294 508350
rect 159362 508294 159418 508350
rect 159486 508294 159542 508350
rect 159114 508170 159170 508226
rect 159238 508170 159294 508226
rect 159362 508170 159418 508226
rect 159486 508170 159542 508226
rect 159114 508046 159170 508102
rect 159238 508046 159294 508102
rect 159362 508046 159418 508102
rect 159486 508046 159542 508102
rect 159114 507922 159170 507978
rect 159238 507922 159294 507978
rect 159362 507922 159418 507978
rect 159486 507922 159542 507978
rect 132114 478294 132170 478350
rect 132238 478294 132294 478350
rect 132362 478294 132418 478350
rect 132486 478294 132542 478350
rect 132114 478170 132170 478226
rect 132238 478170 132294 478226
rect 132362 478170 132418 478226
rect 132486 478170 132542 478226
rect 132114 478046 132170 478102
rect 132238 478046 132294 478102
rect 132362 478046 132418 478102
rect 132486 478046 132542 478102
rect 132114 477922 132170 477978
rect 132238 477922 132294 477978
rect 132362 477922 132418 477978
rect 132486 477922 132542 477978
rect 132114 460294 132170 460350
rect 132238 460294 132294 460350
rect 132362 460294 132418 460350
rect 132486 460294 132542 460350
rect 132114 460170 132170 460226
rect 132238 460170 132294 460226
rect 132362 460170 132418 460226
rect 132486 460170 132542 460226
rect 132114 460046 132170 460102
rect 132238 460046 132294 460102
rect 132362 460046 132418 460102
rect 132486 460046 132542 460102
rect 132114 459922 132170 459978
rect 132238 459922 132294 459978
rect 132362 459922 132418 459978
rect 132486 459922 132542 459978
rect 128394 454294 128450 454350
rect 128518 454294 128574 454350
rect 128642 454294 128698 454350
rect 128766 454294 128822 454350
rect 128394 454170 128450 454226
rect 128518 454170 128574 454226
rect 128642 454170 128698 454226
rect 128766 454170 128822 454226
rect 128394 454046 128450 454102
rect 128518 454046 128574 454102
rect 128642 454046 128698 454102
rect 128766 454046 128822 454102
rect 128394 453922 128450 453978
rect 128518 453922 128574 453978
rect 128642 453922 128698 453978
rect 128766 453922 128822 453978
rect 97674 436294 97730 436350
rect 97798 436294 97854 436350
rect 97922 436294 97978 436350
rect 98046 436294 98102 436350
rect 97674 436170 97730 436226
rect 97798 436170 97854 436226
rect 97922 436170 97978 436226
rect 98046 436170 98102 436226
rect 97674 436046 97730 436102
rect 97798 436046 97854 436102
rect 97922 436046 97978 436102
rect 98046 436046 98102 436102
rect 97674 435922 97730 435978
rect 97798 435922 97854 435978
rect 97922 435922 97978 435978
rect 98046 435922 98102 435978
rect 70674 424294 70730 424350
rect 70798 424294 70854 424350
rect 70922 424294 70978 424350
rect 71046 424294 71102 424350
rect 70674 424170 70730 424226
rect 70798 424170 70854 424226
rect 70922 424170 70978 424226
rect 71046 424170 71102 424226
rect 70674 424046 70730 424102
rect 70798 424046 70854 424102
rect 70922 424046 70978 424102
rect 71046 424046 71102 424102
rect 70674 423922 70730 423978
rect 70798 423922 70854 423978
rect 70922 423922 70978 423978
rect 71046 423922 71102 423978
rect 66954 400294 67010 400350
rect 67078 400294 67134 400350
rect 67202 400294 67258 400350
rect 67326 400294 67382 400350
rect 66954 400170 67010 400226
rect 67078 400170 67134 400226
rect 67202 400170 67258 400226
rect 67326 400170 67382 400226
rect 66954 400046 67010 400102
rect 67078 400046 67134 400102
rect 67202 400046 67258 400102
rect 67326 400046 67382 400102
rect 66954 399922 67010 399978
rect 67078 399922 67134 399978
rect 67202 399922 67258 399978
rect 67326 399922 67382 399978
rect 66954 382294 67010 382350
rect 67078 382294 67134 382350
rect 67202 382294 67258 382350
rect 67326 382294 67382 382350
rect 66954 382170 67010 382226
rect 67078 382170 67134 382226
rect 67202 382170 67258 382226
rect 67326 382170 67382 382226
rect 66954 382046 67010 382102
rect 67078 382046 67134 382102
rect 67202 382046 67258 382102
rect 67326 382046 67382 382102
rect 66954 381922 67010 381978
rect 67078 381922 67134 381978
rect 67202 381922 67258 381978
rect 67326 381922 67382 381978
rect 86518 418294 86574 418350
rect 86642 418294 86698 418350
rect 86518 418170 86574 418226
rect 86642 418170 86698 418226
rect 86518 418046 86574 418102
rect 86642 418046 86698 418102
rect 86518 417922 86574 417978
rect 86642 417922 86698 417978
rect 128394 436294 128450 436350
rect 128518 436294 128574 436350
rect 128642 436294 128698 436350
rect 128766 436294 128822 436350
rect 128394 436170 128450 436226
rect 128518 436170 128574 436226
rect 128642 436170 128698 436226
rect 128766 436170 128822 436226
rect 128394 436046 128450 436102
rect 128518 436046 128574 436102
rect 128642 436046 128698 436102
rect 128766 436046 128822 436102
rect 128394 435922 128450 435978
rect 128518 435922 128574 435978
rect 128642 435922 128698 435978
rect 128766 435922 128822 435978
rect 97674 418294 97730 418350
rect 97798 418294 97854 418350
rect 97922 418294 97978 418350
rect 98046 418294 98102 418350
rect 97674 418170 97730 418226
rect 97798 418170 97854 418226
rect 97922 418170 97978 418226
rect 98046 418170 98102 418226
rect 97674 418046 97730 418102
rect 97798 418046 97854 418102
rect 97922 418046 97978 418102
rect 98046 418046 98102 418102
rect 97674 417922 97730 417978
rect 97798 417922 97854 417978
rect 97922 417922 97978 417978
rect 98046 417922 98102 417978
rect 82684 412442 82740 412498
rect 70674 406294 70730 406350
rect 70798 406294 70854 406350
rect 70922 406294 70978 406350
rect 71046 406294 71102 406350
rect 70674 406170 70730 406226
rect 70798 406170 70854 406226
rect 70922 406170 70978 406226
rect 71046 406170 71102 406226
rect 70674 406046 70730 406102
rect 70798 406046 70854 406102
rect 70922 406046 70978 406102
rect 71046 406046 71102 406102
rect 70674 405922 70730 405978
rect 70798 405922 70854 405978
rect 70922 405922 70978 405978
rect 71046 405922 71102 405978
rect 70674 388294 70730 388350
rect 70798 388294 70854 388350
rect 70922 388294 70978 388350
rect 71046 388294 71102 388350
rect 70674 388170 70730 388226
rect 70798 388170 70854 388226
rect 70922 388170 70978 388226
rect 71046 388170 71102 388226
rect 70674 388046 70730 388102
rect 70798 388046 70854 388102
rect 70922 388046 70978 388102
rect 71046 388046 71102 388102
rect 70674 387922 70730 387978
rect 70798 387922 70854 387978
rect 70922 387922 70978 387978
rect 71046 387922 71102 387978
rect 66954 364294 67010 364350
rect 67078 364294 67134 364350
rect 67202 364294 67258 364350
rect 67326 364294 67382 364350
rect 66954 364170 67010 364226
rect 67078 364170 67134 364226
rect 67202 364170 67258 364226
rect 67326 364170 67382 364226
rect 66954 364046 67010 364102
rect 67078 364046 67134 364102
rect 67202 364046 67258 364102
rect 67326 364046 67382 364102
rect 66954 363922 67010 363978
rect 67078 363922 67134 363978
rect 67202 363922 67258 363978
rect 67326 363922 67382 363978
rect 39878 352294 39934 352350
rect 40002 352294 40058 352350
rect 39878 352170 39934 352226
rect 40002 352170 40058 352226
rect 39878 352046 39934 352102
rect 40002 352046 40058 352102
rect 39878 351922 39934 351978
rect 40002 351922 40058 351978
rect 36234 346294 36290 346350
rect 36358 346294 36414 346350
rect 36482 346294 36538 346350
rect 36606 346294 36662 346350
rect 36234 346170 36290 346226
rect 36358 346170 36414 346226
rect 36482 346170 36538 346226
rect 36606 346170 36662 346226
rect 36234 346046 36290 346102
rect 36358 346046 36414 346102
rect 36482 346046 36538 346102
rect 36606 346046 36662 346102
rect 36234 345922 36290 345978
rect 36358 345922 36414 345978
rect 36482 345922 36538 345978
rect 36606 345922 36662 345978
rect 20076 341702 20132 341758
rect 9234 334294 9290 334350
rect 9358 334294 9414 334350
rect 9482 334294 9538 334350
rect 9606 334294 9662 334350
rect 9234 334170 9290 334226
rect 9358 334170 9414 334226
rect 9482 334170 9538 334226
rect 9606 334170 9662 334226
rect 9234 334046 9290 334102
rect 9358 334046 9414 334102
rect 9482 334046 9538 334102
rect 9606 334046 9662 334102
rect 9234 333922 9290 333978
rect 9358 333922 9414 333978
rect 9482 333922 9538 333978
rect 9606 333922 9662 333978
rect 18060 331802 18116 331858
rect 9234 316294 9290 316350
rect 9358 316294 9414 316350
rect 9482 316294 9538 316350
rect 9606 316294 9662 316350
rect 9234 316170 9290 316226
rect 9358 316170 9414 316226
rect 9482 316170 9538 316226
rect 9606 316170 9662 316226
rect 9234 316046 9290 316102
rect 9358 316046 9414 316102
rect 9482 316046 9538 316102
rect 9606 316046 9662 316102
rect 9234 315922 9290 315978
rect 9358 315922 9414 315978
rect 9482 315922 9538 315978
rect 9606 315922 9662 315978
rect 20636 336122 20692 336178
rect 24518 328294 24574 328350
rect 24642 328294 24698 328350
rect 24518 328170 24574 328226
rect 24642 328170 24698 328226
rect 24518 328046 24574 328102
rect 24642 328046 24698 328102
rect 24518 327922 24574 327978
rect 24642 327922 24698 327978
rect 55238 346294 55294 346350
rect 55362 346294 55418 346350
rect 55238 346170 55294 346226
rect 55362 346170 55418 346226
rect 55238 346046 55294 346102
rect 55362 346046 55418 346102
rect 55238 345922 55294 345978
rect 55362 345922 55418 345978
rect 66954 346294 67010 346350
rect 67078 346294 67134 346350
rect 67202 346294 67258 346350
rect 67326 346294 67382 346350
rect 66954 346170 67010 346226
rect 67078 346170 67134 346226
rect 67202 346170 67258 346226
rect 67326 346170 67382 346226
rect 66954 346046 67010 346102
rect 67078 346046 67134 346102
rect 67202 346046 67258 346102
rect 67326 346046 67382 346102
rect 66954 345922 67010 345978
rect 67078 345922 67134 345978
rect 67202 345922 67258 345978
rect 67326 345922 67382 345978
rect 64204 337562 64260 337618
rect 39878 334294 39934 334350
rect 40002 334294 40058 334350
rect 39878 334170 39934 334226
rect 40002 334170 40058 334226
rect 39878 334046 39934 334102
rect 40002 334046 40058 334102
rect 39878 333922 39934 333978
rect 40002 333922 40058 333978
rect 64204 331442 64260 331498
rect 64204 330362 64260 330418
rect 36234 328294 36290 328350
rect 36358 328294 36414 328350
rect 36482 328294 36538 328350
rect 36606 328294 36662 328350
rect 36234 328170 36290 328226
rect 36358 328170 36414 328226
rect 36482 328170 36538 328226
rect 36606 328170 36662 328226
rect 36234 328046 36290 328102
rect 36358 328046 36414 328102
rect 36482 328046 36538 328102
rect 36606 328046 36662 328102
rect 36234 327922 36290 327978
rect 36358 327922 36414 327978
rect 36482 327922 36538 327978
rect 36606 327922 36662 327978
rect 20076 327482 20132 327538
rect 55238 328294 55294 328350
rect 55362 328294 55418 328350
rect 55238 328170 55294 328226
rect 55362 328170 55418 328226
rect 55238 328046 55294 328102
rect 55362 328046 55418 328102
rect 55238 327922 55294 327978
rect 55362 327922 55418 327978
rect 36234 310294 36290 310350
rect 36358 310294 36414 310350
rect 36482 310294 36538 310350
rect 36606 310294 36662 310350
rect 36234 310170 36290 310226
rect 36358 310170 36414 310226
rect 36482 310170 36538 310226
rect 36606 310170 36662 310226
rect 36234 310046 36290 310102
rect 36358 310046 36414 310102
rect 36482 310046 36538 310102
rect 36606 310046 36662 310102
rect 36234 309922 36290 309978
rect 36358 309922 36414 309978
rect 36482 309922 36538 309978
rect 36606 309922 36662 309978
rect 9234 298294 9290 298350
rect 9358 298294 9414 298350
rect 9482 298294 9538 298350
rect 9606 298294 9662 298350
rect 9234 298170 9290 298226
rect 9358 298170 9414 298226
rect 9482 298170 9538 298226
rect 9606 298170 9662 298226
rect 9234 298046 9290 298102
rect 9358 298046 9414 298102
rect 9482 298046 9538 298102
rect 9606 298046 9662 298102
rect 9234 297922 9290 297978
rect 9358 297922 9414 297978
rect 9482 297922 9538 297978
rect 9606 297922 9662 297978
rect 9234 280294 9290 280350
rect 9358 280294 9414 280350
rect 9482 280294 9538 280350
rect 9606 280294 9662 280350
rect 9234 280170 9290 280226
rect 9358 280170 9414 280226
rect 9482 280170 9538 280226
rect 9606 280170 9662 280226
rect 9234 280046 9290 280102
rect 9358 280046 9414 280102
rect 9482 280046 9538 280102
rect 9606 280046 9662 280102
rect 9234 279922 9290 279978
rect 9358 279922 9414 279978
rect 9482 279922 9538 279978
rect 9606 279922 9662 279978
rect 65212 330902 65268 330958
rect 82684 409022 82740 409078
rect 117238 418294 117294 418350
rect 117362 418294 117418 418350
rect 117238 418170 117294 418226
rect 117362 418170 117418 418226
rect 117238 418046 117294 418102
rect 117362 418046 117418 418102
rect 117238 417922 117294 417978
rect 117362 417922 117418 417978
rect 128394 418294 128450 418350
rect 128518 418294 128574 418350
rect 128642 418294 128698 418350
rect 128766 418294 128822 418350
rect 128394 418170 128450 418226
rect 128518 418170 128574 418226
rect 128642 418170 128698 418226
rect 128766 418170 128822 418226
rect 128394 418046 128450 418102
rect 128518 418046 128574 418102
rect 128642 418046 128698 418102
rect 128766 418046 128822 418102
rect 128394 417922 128450 417978
rect 128518 417922 128574 417978
rect 128642 417922 128698 417978
rect 128766 417922 128822 417978
rect 82348 406682 82404 406738
rect 125132 406682 125188 406738
rect 101878 406294 101934 406350
rect 102002 406294 102058 406350
rect 101878 406170 101934 406226
rect 102002 406170 102058 406226
rect 101878 406046 101934 406102
rect 102002 406046 102058 406102
rect 101878 405922 101934 405978
rect 102002 405922 102058 405978
rect 86518 400294 86574 400350
rect 86642 400294 86698 400350
rect 86518 400170 86574 400226
rect 86642 400170 86698 400226
rect 86518 400046 86574 400102
rect 86642 400046 86698 400102
rect 86518 399922 86574 399978
rect 86642 399922 86698 399978
rect 117238 400294 117294 400350
rect 117362 400294 117418 400350
rect 117238 400170 117294 400226
rect 117362 400170 117418 400226
rect 117238 400046 117294 400102
rect 117362 400046 117418 400102
rect 117238 399922 117294 399978
rect 117362 399922 117418 399978
rect 82348 398042 82404 398098
rect 126252 402362 126308 402418
rect 125132 396422 125188 396478
rect 101836 388333 101892 388389
rect 101940 388333 101996 388389
rect 102044 388333 102100 388389
rect 97674 382294 97730 382350
rect 97798 382294 97854 382350
rect 97922 382294 97978 382350
rect 98046 382294 98102 382350
rect 97674 382170 97730 382226
rect 97798 382170 97854 382226
rect 97922 382170 97978 382226
rect 98046 382170 98102 382226
rect 97674 382046 97730 382102
rect 97798 382046 97854 382102
rect 97922 382046 97978 382102
rect 98046 382046 98102 382102
rect 97674 381922 97730 381978
rect 97798 381922 97854 381978
rect 97922 381922 97978 381978
rect 98046 381922 98102 381978
rect 70674 370294 70730 370350
rect 70798 370294 70854 370350
rect 70922 370294 70978 370350
rect 71046 370294 71102 370350
rect 70674 370170 70730 370226
rect 70798 370170 70854 370226
rect 70922 370170 70978 370226
rect 71046 370170 71102 370226
rect 70674 370046 70730 370102
rect 70798 370046 70854 370102
rect 70922 370046 70978 370102
rect 71046 370046 71102 370102
rect 70674 369922 70730 369978
rect 70798 369922 70854 369978
rect 70922 369922 70978 369978
rect 71046 369922 71102 369978
rect 70674 352294 70730 352350
rect 70798 352294 70854 352350
rect 70922 352294 70978 352350
rect 71046 352294 71102 352350
rect 70674 352170 70730 352226
rect 70798 352170 70854 352226
rect 70922 352170 70978 352226
rect 71046 352170 71102 352226
rect 70674 352046 70730 352102
rect 70798 352046 70854 352102
rect 70922 352046 70978 352102
rect 71046 352046 71102 352102
rect 70674 351922 70730 351978
rect 70798 351922 70854 351978
rect 70922 351922 70978 351978
rect 71046 351922 71102 351978
rect 128394 400294 128450 400350
rect 128518 400294 128574 400350
rect 128642 400294 128698 400350
rect 128766 400294 128822 400350
rect 128394 400170 128450 400226
rect 128518 400170 128574 400226
rect 128642 400170 128698 400226
rect 128766 400170 128822 400226
rect 128394 400046 128450 400102
rect 128518 400046 128574 400102
rect 128642 400046 128698 400102
rect 128766 400046 128822 400102
rect 128394 399922 128450 399978
rect 128518 399922 128574 399978
rect 128642 399922 128698 399978
rect 128766 399922 128822 399978
rect 128394 382294 128450 382350
rect 128518 382294 128574 382350
rect 128642 382294 128698 382350
rect 128766 382294 128822 382350
rect 128394 382170 128450 382226
rect 128518 382170 128574 382226
rect 128642 382170 128698 382226
rect 128766 382170 128822 382226
rect 128394 382046 128450 382102
rect 128518 382046 128574 382102
rect 128642 382046 128698 382102
rect 128766 382046 128822 382102
rect 128394 381922 128450 381978
rect 128518 381922 128574 381978
rect 128642 381922 128698 381978
rect 128766 381922 128822 381978
rect 97674 364294 97730 364350
rect 97798 364294 97854 364350
rect 97922 364294 97978 364350
rect 98046 364294 98102 364350
rect 97674 364170 97730 364226
rect 97798 364170 97854 364226
rect 97922 364170 97978 364226
rect 98046 364170 98102 364226
rect 97674 364046 97730 364102
rect 97798 364046 97854 364102
rect 97922 364046 97978 364102
rect 98046 364046 98102 364102
rect 97674 363922 97730 363978
rect 97798 363922 97854 363978
rect 97922 363922 97978 363978
rect 98046 363922 98102 363978
rect 86518 346294 86574 346350
rect 86642 346294 86698 346350
rect 86518 346170 86574 346226
rect 86642 346170 86698 346226
rect 86518 346046 86574 346102
rect 86642 346046 86698 346102
rect 86518 345922 86574 345978
rect 86642 345922 86698 345978
rect 128394 364294 128450 364350
rect 128518 364294 128574 364350
rect 128642 364294 128698 364350
rect 128766 364294 128822 364350
rect 128394 364170 128450 364226
rect 128518 364170 128574 364226
rect 128642 364170 128698 364226
rect 128766 364170 128822 364226
rect 128394 364046 128450 364102
rect 128518 364046 128574 364102
rect 128642 364046 128698 364102
rect 128766 364046 128822 364102
rect 128394 363922 128450 363978
rect 128518 363922 128574 363978
rect 128642 363922 128698 363978
rect 128766 363922 128822 363978
rect 101878 352294 101934 352350
rect 102002 352294 102058 352350
rect 101878 352170 101934 352226
rect 102002 352170 102058 352226
rect 101878 352046 101934 352102
rect 102002 352046 102058 352102
rect 101878 351922 101934 351978
rect 102002 351922 102058 351978
rect 97674 346294 97730 346350
rect 97798 346294 97854 346350
rect 97922 346294 97978 346350
rect 98046 346294 98102 346350
rect 97674 346170 97730 346226
rect 97798 346170 97854 346226
rect 97922 346170 97978 346226
rect 98046 346170 98102 346226
rect 97674 346046 97730 346102
rect 97798 346046 97854 346102
rect 97922 346046 97978 346102
rect 98046 346046 98102 346102
rect 97674 345922 97730 345978
rect 97798 345922 97854 345978
rect 97922 345922 97978 345978
rect 98046 345922 98102 345978
rect 82684 341882 82740 341938
rect 82460 340284 82516 340318
rect 82460 340262 82516 340284
rect 82236 338462 82292 338518
rect 70674 334294 70730 334350
rect 70798 334294 70854 334350
rect 70922 334294 70978 334350
rect 71046 334294 71102 334350
rect 70674 334170 70730 334226
rect 70798 334170 70854 334226
rect 70922 334170 70978 334226
rect 71046 334170 71102 334226
rect 70674 334046 70730 334102
rect 70798 334046 70854 334102
rect 70922 334046 70978 334102
rect 71046 334046 71102 334102
rect 70674 333922 70730 333978
rect 70798 333922 70854 333978
rect 70922 333922 70978 333978
rect 71046 333922 71102 333978
rect 66954 328294 67010 328350
rect 67078 328294 67134 328350
rect 67202 328294 67258 328350
rect 67326 328294 67382 328350
rect 66954 328170 67010 328226
rect 67078 328170 67134 328226
rect 67202 328170 67258 328226
rect 67326 328170 67382 328226
rect 66954 328046 67010 328102
rect 67078 328046 67134 328102
rect 67202 328046 67258 328102
rect 67326 328046 67382 328102
rect 66954 327922 67010 327978
rect 67078 327922 67134 327978
rect 67202 327922 67258 327978
rect 67326 327922 67382 327978
rect 66954 310294 67010 310350
rect 67078 310294 67134 310350
rect 67202 310294 67258 310350
rect 67326 310294 67382 310350
rect 66954 310170 67010 310226
rect 67078 310170 67134 310226
rect 67202 310170 67258 310226
rect 67326 310170 67382 310226
rect 66954 310046 67010 310102
rect 67078 310046 67134 310102
rect 67202 310046 67258 310102
rect 67326 310046 67382 310102
rect 66954 309922 67010 309978
rect 67078 309922 67134 309978
rect 67202 309922 67258 309978
rect 67326 309922 67382 309978
rect 36234 292294 36290 292350
rect 36358 292294 36414 292350
rect 36482 292294 36538 292350
rect 36606 292294 36662 292350
rect 36234 292170 36290 292226
rect 36358 292170 36414 292226
rect 36482 292170 36538 292226
rect 36606 292170 36662 292226
rect 36234 292046 36290 292102
rect 36358 292046 36414 292102
rect 36482 292046 36538 292102
rect 36606 292046 36662 292102
rect 36234 291922 36290 291978
rect 36358 291922 36414 291978
rect 36482 291922 36538 291978
rect 36606 291922 36662 291978
rect 24518 274294 24574 274350
rect 24642 274294 24698 274350
rect 24518 274170 24574 274226
rect 24642 274170 24698 274226
rect 24518 274046 24574 274102
rect 24642 274046 24698 274102
rect 24518 273922 24574 273978
rect 24642 273922 24698 273978
rect 70674 316294 70730 316350
rect 70798 316294 70854 316350
rect 70922 316294 70978 316350
rect 71046 316294 71102 316350
rect 70674 316170 70730 316226
rect 70798 316170 70854 316226
rect 70922 316170 70978 316226
rect 71046 316170 71102 316226
rect 70674 316046 70730 316102
rect 70798 316046 70854 316102
rect 70922 316046 70978 316102
rect 71046 316046 71102 316102
rect 70674 315922 70730 315978
rect 70798 315922 70854 315978
rect 70922 315922 70978 315978
rect 71046 315922 71102 315978
rect 66954 292294 67010 292350
rect 67078 292294 67134 292350
rect 67202 292294 67258 292350
rect 67326 292294 67382 292350
rect 66954 292170 67010 292226
rect 67078 292170 67134 292226
rect 67202 292170 67258 292226
rect 67326 292170 67382 292226
rect 66954 292046 67010 292102
rect 67078 292046 67134 292102
rect 67202 292046 67258 292102
rect 67326 292046 67382 292102
rect 66954 291922 67010 291978
rect 67078 291922 67134 291978
rect 67202 291922 67258 291978
rect 67326 291922 67382 291978
rect 39878 280294 39934 280350
rect 40002 280294 40058 280350
rect 39878 280170 39934 280226
rect 40002 280170 40058 280226
rect 39878 280046 39934 280102
rect 40002 280046 40058 280102
rect 39878 279922 39934 279978
rect 40002 279922 40058 279978
rect 64204 275642 64260 275698
rect 36234 274294 36290 274350
rect 36358 274294 36414 274350
rect 36482 274294 36538 274350
rect 36606 274294 36662 274350
rect 36234 274170 36290 274226
rect 36358 274170 36414 274226
rect 36482 274170 36538 274226
rect 36606 274170 36662 274226
rect 36234 274046 36290 274102
rect 36358 274046 36414 274102
rect 36482 274046 36538 274102
rect 36606 274046 36662 274102
rect 36234 273922 36290 273978
rect 36358 273922 36414 273978
rect 36482 273922 36538 273978
rect 36606 273922 36662 273978
rect 20076 270452 20132 270478
rect 20076 270422 20132 270452
rect 9234 262294 9290 262350
rect 9358 262294 9414 262350
rect 9482 262294 9538 262350
rect 9606 262294 9662 262350
rect 9234 262170 9290 262226
rect 9358 262170 9414 262226
rect 9482 262170 9538 262226
rect 9606 262170 9662 262226
rect 9234 262046 9290 262102
rect 9358 262046 9414 262102
rect 9482 262046 9538 262102
rect 9606 262046 9662 262102
rect 9234 261922 9290 261978
rect 9358 261922 9414 261978
rect 9482 261922 9538 261978
rect 9606 261922 9662 261978
rect 55238 274294 55294 274350
rect 55362 274294 55418 274350
rect 55238 274170 55294 274226
rect 55362 274170 55418 274226
rect 55238 274046 55294 274102
rect 55362 274046 55418 274102
rect 55238 273922 55294 273978
rect 55362 273922 55418 273978
rect 66954 274294 67010 274350
rect 67078 274294 67134 274350
rect 67202 274294 67258 274350
rect 67326 274294 67382 274350
rect 66954 274170 67010 274226
rect 67078 274170 67134 274226
rect 67202 274170 67258 274226
rect 67326 274170 67382 274226
rect 66954 274046 67010 274102
rect 67078 274046 67134 274102
rect 67202 274046 67258 274102
rect 67326 274046 67382 274102
rect 66954 273922 67010 273978
rect 67078 273922 67134 273978
rect 67202 273922 67258 273978
rect 67326 273922 67382 273978
rect 64652 270782 64708 270838
rect 64204 270242 64260 270298
rect 64204 270062 64260 270118
rect 64204 268622 64260 268678
rect 9234 244294 9290 244350
rect 9358 244294 9414 244350
rect 9482 244294 9538 244350
rect 9606 244294 9662 244350
rect 9234 244170 9290 244226
rect 9358 244170 9414 244226
rect 9482 244170 9538 244226
rect 9606 244170 9662 244226
rect 9234 244046 9290 244102
rect 9358 244046 9414 244102
rect 9482 244046 9538 244102
rect 9606 244046 9662 244102
rect 9234 243922 9290 243978
rect 9358 243922 9414 243978
rect 9482 243922 9538 243978
rect 9606 243922 9662 243978
rect 64204 264482 64260 264538
rect 39878 262294 39934 262350
rect 40002 262294 40058 262350
rect 39878 262170 39934 262226
rect 40002 262170 40058 262226
rect 39878 262046 39934 262102
rect 40002 262046 40058 262102
rect 39878 261922 39934 261978
rect 40002 261922 40058 261978
rect 24518 256294 24574 256350
rect 24642 256294 24698 256350
rect 24518 256170 24574 256226
rect 24642 256170 24698 256226
rect 24518 256046 24574 256102
rect 24642 256046 24698 256102
rect 24518 255922 24574 255978
rect 24642 255922 24698 255978
rect 36234 256294 36290 256350
rect 36358 256294 36414 256350
rect 36482 256294 36538 256350
rect 36606 256294 36662 256350
rect 36234 256170 36290 256226
rect 36358 256170 36414 256226
rect 36482 256170 36538 256226
rect 36606 256170 36662 256226
rect 36234 256046 36290 256102
rect 36358 256046 36414 256102
rect 36482 256046 36538 256102
rect 36606 256046 36662 256102
rect 36234 255922 36290 255978
rect 36358 255922 36414 255978
rect 36482 255922 36538 255978
rect 36606 255922 36662 255978
rect 9234 226294 9290 226350
rect 9358 226294 9414 226350
rect 9482 226294 9538 226350
rect 9606 226294 9662 226350
rect 9234 226170 9290 226226
rect 9358 226170 9414 226226
rect 9482 226170 9538 226226
rect 9606 226170 9662 226226
rect 9234 226046 9290 226102
rect 9358 226046 9414 226102
rect 9482 226046 9538 226102
rect 9606 226046 9662 226102
rect 9234 225922 9290 225978
rect 9358 225922 9414 225978
rect 9482 225922 9538 225978
rect 9606 225922 9662 225978
rect 55238 256294 55294 256350
rect 55362 256294 55418 256350
rect 55238 256170 55294 256226
rect 55362 256170 55418 256226
rect 55238 256046 55294 256102
rect 55362 256046 55418 256102
rect 55238 255922 55294 255978
rect 55362 255922 55418 255978
rect 86518 328294 86574 328350
rect 86642 328294 86698 328350
rect 86518 328170 86574 328226
rect 86642 328170 86698 328226
rect 86518 328046 86574 328102
rect 86642 328046 86698 328102
rect 86518 327922 86574 327978
rect 86642 327922 86698 327978
rect 117238 346294 117294 346350
rect 117362 346294 117418 346350
rect 117238 346170 117294 346226
rect 117362 346170 117418 346226
rect 117238 346046 117294 346102
rect 117362 346046 117418 346102
rect 117238 345922 117294 345978
rect 117362 345922 117418 345978
rect 128394 346294 128450 346350
rect 128518 346294 128574 346350
rect 128642 346294 128698 346350
rect 128766 346294 128822 346350
rect 128394 346170 128450 346226
rect 128518 346170 128574 346226
rect 128642 346170 128698 346226
rect 128766 346170 128822 346226
rect 128394 346046 128450 346102
rect 128518 346046 128574 346102
rect 128642 346046 128698 346102
rect 128766 346046 128822 346102
rect 128394 345922 128450 345978
rect 128518 345922 128574 345978
rect 128642 345922 128698 345978
rect 128766 345922 128822 345978
rect 122668 340442 122724 340498
rect 122668 338462 122724 338518
rect 124348 336122 124404 336178
rect 101878 334294 101934 334350
rect 102002 334294 102058 334350
rect 101878 334170 101934 334226
rect 102002 334170 102058 334226
rect 101878 334046 101934 334102
rect 102002 334046 102058 334102
rect 101878 333922 101934 333978
rect 102002 333922 102058 333978
rect 97674 328294 97730 328350
rect 97798 328294 97854 328350
rect 97922 328294 97978 328350
rect 98046 328294 98102 328350
rect 97674 328170 97730 328226
rect 97798 328170 97854 328226
rect 97922 328170 97978 328226
rect 98046 328170 98102 328226
rect 97674 328046 97730 328102
rect 97798 328046 97854 328102
rect 97922 328046 97978 328102
rect 98046 328046 98102 328102
rect 97674 327922 97730 327978
rect 97798 327922 97854 327978
rect 97922 327922 97978 327978
rect 98046 327922 98102 327978
rect 117238 328294 117294 328350
rect 117362 328294 117418 328350
rect 117238 328170 117294 328226
rect 117362 328170 117418 328226
rect 117238 328046 117294 328102
rect 117362 328046 117418 328102
rect 117238 327922 117294 327978
rect 117362 327922 117418 327978
rect 127596 339182 127652 339238
rect 127596 336122 127652 336178
rect 127596 332702 127652 332758
rect 127596 330722 127652 330778
rect 124348 327302 124404 327358
rect 141036 483002 141092 483058
rect 140924 466082 140980 466138
rect 132114 442294 132170 442350
rect 132238 442294 132294 442350
rect 132362 442294 132418 442350
rect 132486 442294 132542 442350
rect 132114 442170 132170 442226
rect 132238 442170 132294 442226
rect 132362 442170 132418 442226
rect 132486 442170 132542 442226
rect 132114 442046 132170 442102
rect 132238 442046 132294 442102
rect 132362 442046 132418 442102
rect 132486 442046 132542 442102
rect 132114 441922 132170 441978
rect 132238 441922 132294 441978
rect 132362 441922 132418 441978
rect 132486 441922 132542 441978
rect 148518 490294 148574 490350
rect 148642 490294 148698 490350
rect 148518 490170 148574 490226
rect 148642 490170 148698 490226
rect 148518 490046 148574 490102
rect 148642 490046 148698 490102
rect 148518 489922 148574 489978
rect 148642 489922 148698 489978
rect 159114 490294 159170 490350
rect 159238 490294 159294 490350
rect 159362 490294 159418 490350
rect 159486 490294 159542 490350
rect 159114 490170 159170 490226
rect 159238 490170 159294 490226
rect 159362 490170 159418 490226
rect 159486 490170 159542 490226
rect 159114 490046 159170 490102
rect 159238 490046 159294 490102
rect 159362 490046 159418 490102
rect 159486 490046 159542 490102
rect 159114 489922 159170 489978
rect 159238 489922 159294 489978
rect 159362 489922 159418 489978
rect 159486 489922 159542 489978
rect 148518 472294 148574 472350
rect 148642 472294 148698 472350
rect 148518 472170 148574 472226
rect 148642 472170 148698 472226
rect 148518 472046 148574 472102
rect 148642 472046 148698 472102
rect 148518 471922 148574 471978
rect 148642 471922 148698 471978
rect 159114 472294 159170 472350
rect 159238 472294 159294 472350
rect 159362 472294 159418 472350
rect 159486 472294 159542 472350
rect 159114 472170 159170 472226
rect 159238 472170 159294 472226
rect 159362 472170 159418 472226
rect 159486 472170 159542 472226
rect 159114 472046 159170 472102
rect 159238 472046 159294 472102
rect 159362 472046 159418 472102
rect 159486 472046 159542 472102
rect 159114 471922 159170 471978
rect 159238 471922 159294 471978
rect 159362 471922 159418 471978
rect 159486 471922 159542 471978
rect 144396 469502 144452 469558
rect 162834 532294 162890 532350
rect 162958 532294 163014 532350
rect 163082 532294 163138 532350
rect 163206 532294 163262 532350
rect 162834 532170 162890 532226
rect 162958 532170 163014 532226
rect 163082 532170 163138 532226
rect 163206 532170 163262 532226
rect 162834 532046 162890 532102
rect 162958 532046 163014 532102
rect 163082 532046 163138 532102
rect 163206 532046 163262 532102
rect 162834 531922 162890 531978
rect 162958 531922 163014 531978
rect 163082 531922 163138 531978
rect 163206 531922 163262 531978
rect 163878 532294 163934 532350
rect 164002 532294 164058 532350
rect 163878 532170 163934 532226
rect 164002 532170 164058 532226
rect 163878 532046 163934 532102
rect 164002 532046 164058 532102
rect 163878 531922 163934 531978
rect 164002 531922 164058 531978
rect 162834 514294 162890 514350
rect 162958 514294 163014 514350
rect 163082 514294 163138 514350
rect 163206 514294 163262 514350
rect 162834 514170 162890 514226
rect 162958 514170 163014 514226
rect 163082 514170 163138 514226
rect 163206 514170 163262 514226
rect 162834 514046 162890 514102
rect 162958 514046 163014 514102
rect 163082 514046 163138 514102
rect 163206 514046 163262 514102
rect 162834 513922 162890 513978
rect 162958 513922 163014 513978
rect 163082 513922 163138 513978
rect 163206 513922 163262 513978
rect 189834 544294 189890 544350
rect 189958 544294 190014 544350
rect 190082 544294 190138 544350
rect 190206 544294 190262 544350
rect 189834 544170 189890 544226
rect 189958 544170 190014 544226
rect 190082 544170 190138 544226
rect 190206 544170 190262 544226
rect 189834 544046 189890 544102
rect 189958 544046 190014 544102
rect 190082 544046 190138 544102
rect 190206 544046 190262 544102
rect 189834 543922 189890 543978
rect 189958 543922 190014 543978
rect 190082 543922 190138 543978
rect 190206 543922 190262 543978
rect 189834 526294 189890 526350
rect 189958 526294 190014 526350
rect 190082 526294 190138 526350
rect 190206 526294 190262 526350
rect 189834 526170 189890 526226
rect 189958 526170 190014 526226
rect 190082 526170 190138 526226
rect 190206 526170 190262 526226
rect 189834 526046 189890 526102
rect 189958 526046 190014 526102
rect 190082 526046 190138 526102
rect 190206 526046 190262 526102
rect 189834 525922 189890 525978
rect 189958 525922 190014 525978
rect 190082 525922 190138 525978
rect 190206 525922 190262 525978
rect 189834 508294 189890 508350
rect 189958 508294 190014 508350
rect 190082 508294 190138 508350
rect 190206 508294 190262 508350
rect 189834 508170 189890 508226
rect 189958 508170 190014 508226
rect 190082 508170 190138 508226
rect 190206 508170 190262 508226
rect 189834 508046 189890 508102
rect 189958 508046 190014 508102
rect 190082 508046 190138 508102
rect 190206 508046 190262 508102
rect 189834 507922 189890 507978
rect 189958 507922 190014 507978
rect 190082 507922 190138 507978
rect 190206 507922 190262 507978
rect 162834 496294 162890 496350
rect 162958 496294 163014 496350
rect 163082 496294 163138 496350
rect 163206 496294 163262 496350
rect 162834 496170 162890 496226
rect 162958 496170 163014 496226
rect 163082 496170 163138 496226
rect 163206 496170 163262 496226
rect 162834 496046 162890 496102
rect 162958 496046 163014 496102
rect 163082 496046 163138 496102
rect 163206 496046 163262 496102
rect 162834 495922 162890 495978
rect 162958 495922 163014 495978
rect 163082 495922 163138 495978
rect 163206 495922 163262 495978
rect 179238 490294 179294 490350
rect 179362 490294 179418 490350
rect 179238 490170 179294 490226
rect 179362 490170 179418 490226
rect 179238 490046 179294 490102
rect 179362 490046 179418 490102
rect 179238 489922 179294 489978
rect 179362 489922 179418 489978
rect 189834 490294 189890 490350
rect 189958 490294 190014 490350
rect 190082 490294 190138 490350
rect 190206 490294 190262 490350
rect 189834 490170 189890 490226
rect 189958 490170 190014 490226
rect 190082 490170 190138 490226
rect 190206 490170 190262 490226
rect 189834 490046 189890 490102
rect 189958 490046 190014 490102
rect 190082 490046 190138 490102
rect 190206 490046 190262 490102
rect 189834 489922 189890 489978
rect 189958 489922 190014 489978
rect 190082 489922 190138 489978
rect 190206 489922 190262 489978
rect 162834 478294 162890 478350
rect 162958 478294 163014 478350
rect 163082 478294 163138 478350
rect 163206 478294 163262 478350
rect 162834 478170 162890 478226
rect 162958 478170 163014 478226
rect 163082 478170 163138 478226
rect 163206 478170 163262 478226
rect 162834 478046 162890 478102
rect 162958 478046 163014 478102
rect 163082 478046 163138 478102
rect 163206 478046 163262 478102
rect 162834 477922 162890 477978
rect 162958 477922 163014 477978
rect 163082 477922 163138 477978
rect 163206 477922 163262 477978
rect 163878 478294 163934 478350
rect 164002 478294 164058 478350
rect 163878 478170 163934 478226
rect 164002 478170 164058 478226
rect 163878 478046 163934 478102
rect 164002 478046 164058 478102
rect 163878 477922 163934 477978
rect 164002 477922 164058 477978
rect 179238 472294 179294 472350
rect 179362 472294 179418 472350
rect 179238 472170 179294 472226
rect 179362 472170 179418 472226
rect 179238 472046 179294 472102
rect 179362 472046 179418 472102
rect 179238 471922 179294 471978
rect 179362 471922 179418 471978
rect 189532 475442 189588 475498
rect 189532 473822 189588 473878
rect 189834 472294 189890 472350
rect 189958 472294 190014 472350
rect 190082 472294 190138 472350
rect 190206 472294 190262 472350
rect 189834 472170 189890 472226
rect 189958 472170 190014 472226
rect 190082 472170 190138 472226
rect 190206 472170 190262 472226
rect 189834 472046 189890 472102
rect 189958 472046 190014 472102
rect 190082 472046 190138 472102
rect 190206 472046 190262 472102
rect 189834 471922 189890 471978
rect 189958 471922 190014 471978
rect 190082 471922 190138 471978
rect 190206 471922 190262 471978
rect 162834 460294 162890 460350
rect 162958 460294 163014 460350
rect 163082 460294 163138 460350
rect 163206 460294 163262 460350
rect 162834 460170 162890 460226
rect 162958 460170 163014 460226
rect 163082 460170 163138 460226
rect 163206 460170 163262 460226
rect 162834 460046 162890 460102
rect 162958 460046 163014 460102
rect 163082 460046 163138 460102
rect 163206 460046 163262 460102
rect 162834 459922 162890 459978
rect 162958 459922 163014 459978
rect 163082 459922 163138 459978
rect 163206 459922 163262 459978
rect 159114 454294 159170 454350
rect 159238 454294 159294 454350
rect 159362 454294 159418 454350
rect 159486 454294 159542 454350
rect 159114 454170 159170 454226
rect 159238 454170 159294 454226
rect 159362 454170 159418 454226
rect 159486 454170 159542 454226
rect 159114 454046 159170 454102
rect 159238 454046 159294 454102
rect 159362 454046 159418 454102
rect 159486 454046 159542 454102
rect 159114 453922 159170 453978
rect 159238 453922 159294 453978
rect 159362 453922 159418 453978
rect 159486 453922 159542 453978
rect 159114 436294 159170 436350
rect 159238 436294 159294 436350
rect 159362 436294 159418 436350
rect 159486 436294 159542 436350
rect 159114 436170 159170 436226
rect 159238 436170 159294 436226
rect 159362 436170 159418 436226
rect 159486 436170 159542 436226
rect 159114 436046 159170 436102
rect 159238 436046 159294 436102
rect 159362 436046 159418 436102
rect 159486 436046 159542 436102
rect 159114 435922 159170 435978
rect 159238 435922 159294 435978
rect 159362 435922 159418 435978
rect 159486 435922 159542 435978
rect 132114 424294 132170 424350
rect 132238 424294 132294 424350
rect 132362 424294 132418 424350
rect 132486 424294 132542 424350
rect 132114 424170 132170 424226
rect 132238 424170 132294 424226
rect 132362 424170 132418 424226
rect 132486 424170 132542 424226
rect 132114 424046 132170 424102
rect 132238 424046 132294 424102
rect 132362 424046 132418 424102
rect 132486 424046 132542 424102
rect 132114 423922 132170 423978
rect 132238 423922 132294 423978
rect 132362 423922 132418 423978
rect 132486 423922 132542 423978
rect 148518 418294 148574 418350
rect 148642 418294 148698 418350
rect 148518 418170 148574 418226
rect 148642 418170 148698 418226
rect 148518 418046 148574 418102
rect 148642 418046 148698 418102
rect 148518 417922 148574 417978
rect 148642 417922 148698 417978
rect 159114 418294 159170 418350
rect 159238 418294 159294 418350
rect 159362 418294 159418 418350
rect 159486 418294 159542 418350
rect 159114 418170 159170 418226
rect 159238 418170 159294 418226
rect 159362 418170 159418 418226
rect 159486 418170 159542 418226
rect 159114 418046 159170 418102
rect 159238 418046 159294 418102
rect 159362 418046 159418 418102
rect 159486 418046 159542 418102
rect 159114 417922 159170 417978
rect 159238 417922 159294 417978
rect 159362 417922 159418 417978
rect 159486 417922 159542 417978
rect 144060 412622 144116 412678
rect 141036 412442 141092 412498
rect 132114 406294 132170 406350
rect 132238 406294 132294 406350
rect 132362 406294 132418 406350
rect 132486 406294 132542 406350
rect 132114 406170 132170 406226
rect 132238 406170 132294 406226
rect 132362 406170 132418 406226
rect 132486 406170 132542 406226
rect 132114 406046 132170 406102
rect 132238 406046 132294 406102
rect 132362 406046 132418 406102
rect 132486 406046 132542 406102
rect 132114 405922 132170 405978
rect 132238 405922 132294 405978
rect 132362 405922 132418 405978
rect 132486 405922 132542 405978
rect 132114 388294 132170 388350
rect 132238 388294 132294 388350
rect 132362 388294 132418 388350
rect 132486 388294 132542 388350
rect 132114 388170 132170 388226
rect 132238 388170 132294 388226
rect 132362 388170 132418 388226
rect 132486 388170 132542 388226
rect 132114 388046 132170 388102
rect 132238 388046 132294 388102
rect 132362 388046 132418 388102
rect 132486 388046 132542 388102
rect 132114 387922 132170 387978
rect 132238 387922 132294 387978
rect 132362 387922 132418 387978
rect 132486 387922 132542 387978
rect 136108 399662 136164 399718
rect 135212 393002 135268 393058
rect 144284 409922 144340 409978
rect 144284 408302 144340 408358
rect 144396 406682 144452 406738
rect 144284 404162 144340 404218
rect 132114 370294 132170 370350
rect 132238 370294 132294 370350
rect 132362 370294 132418 370350
rect 132486 370294 132542 370350
rect 132114 370170 132170 370226
rect 132238 370170 132294 370226
rect 132362 370170 132418 370226
rect 132486 370170 132542 370226
rect 132114 370046 132170 370102
rect 132238 370046 132294 370102
rect 132362 370046 132418 370102
rect 132486 370046 132542 370102
rect 132114 369922 132170 369978
rect 132238 369922 132294 369978
rect 132362 369922 132418 369978
rect 132486 369922 132542 369978
rect 148518 400294 148574 400350
rect 148642 400294 148698 400350
rect 148518 400170 148574 400226
rect 148642 400170 148698 400226
rect 148518 400046 148574 400102
rect 148642 400046 148698 400102
rect 148518 399922 148574 399978
rect 148642 399922 148698 399978
rect 159114 400294 159170 400350
rect 159238 400294 159294 400350
rect 159362 400294 159418 400350
rect 159486 400294 159542 400350
rect 159114 400170 159170 400226
rect 159238 400170 159294 400226
rect 159362 400170 159418 400226
rect 159486 400170 159542 400226
rect 159114 400046 159170 400102
rect 159238 400046 159294 400102
rect 159362 400046 159418 400102
rect 159486 400046 159542 400102
rect 159114 399922 159170 399978
rect 159238 399922 159294 399978
rect 159362 399922 159418 399978
rect 159486 399922 159542 399978
rect 159114 382294 159170 382350
rect 159238 382294 159294 382350
rect 159362 382294 159418 382350
rect 159486 382294 159542 382350
rect 159114 382170 159170 382226
rect 159238 382170 159294 382226
rect 159362 382170 159418 382226
rect 159486 382170 159542 382226
rect 159114 382046 159170 382102
rect 159238 382046 159294 382102
rect 159362 382046 159418 382102
rect 159486 382046 159542 382102
rect 159114 381922 159170 381978
rect 159238 381922 159294 381978
rect 159362 381922 159418 381978
rect 159486 381922 159542 381978
rect 159114 364294 159170 364350
rect 159238 364294 159294 364350
rect 159362 364294 159418 364350
rect 159486 364294 159542 364350
rect 159114 364170 159170 364226
rect 159238 364170 159294 364226
rect 159362 364170 159418 364226
rect 159486 364170 159542 364226
rect 132114 352294 132170 352350
rect 132238 352294 132294 352350
rect 132362 352294 132418 352350
rect 132486 352294 132542 352350
rect 132114 352170 132170 352226
rect 132238 352170 132294 352226
rect 132362 352170 132418 352226
rect 132486 352170 132542 352226
rect 132114 352046 132170 352102
rect 132238 352046 132294 352102
rect 132362 352046 132418 352102
rect 132486 352046 132542 352102
rect 132114 351922 132170 351978
rect 132238 351922 132294 351978
rect 132362 351922 132418 351978
rect 132486 351922 132542 351978
rect 130060 341702 130116 341758
rect 128394 328294 128450 328350
rect 128518 328294 128574 328350
rect 128642 328294 128698 328350
rect 128766 328294 128822 328350
rect 128394 328170 128450 328226
rect 128518 328170 128574 328226
rect 128642 328170 128698 328226
rect 128766 328170 128822 328226
rect 128394 328046 128450 328102
rect 128518 328046 128574 328102
rect 128642 328046 128698 328102
rect 128766 328046 128822 328102
rect 128394 327922 128450 327978
rect 128518 327922 128574 327978
rect 128642 327922 128698 327978
rect 128766 327922 128822 327978
rect 97674 310294 97730 310350
rect 97798 310294 97854 310350
rect 97922 310294 97978 310350
rect 98046 310294 98102 310350
rect 97674 310170 97730 310226
rect 97798 310170 97854 310226
rect 97922 310170 97978 310226
rect 98046 310170 98102 310226
rect 97674 310046 97730 310102
rect 97798 310046 97854 310102
rect 97922 310046 97978 310102
rect 98046 310046 98102 310102
rect 97674 309922 97730 309978
rect 97798 309922 97854 309978
rect 97922 309922 97978 309978
rect 98046 309922 98102 309978
rect 70674 298294 70730 298350
rect 70798 298294 70854 298350
rect 70922 298294 70978 298350
rect 71046 298294 71102 298350
rect 70674 298170 70730 298226
rect 70798 298170 70854 298226
rect 70922 298170 70978 298226
rect 71046 298170 71102 298226
rect 70674 298046 70730 298102
rect 70798 298046 70854 298102
rect 70922 298046 70978 298102
rect 71046 298046 71102 298102
rect 70674 297922 70730 297978
rect 70798 297922 70854 297978
rect 70922 297922 70978 297978
rect 71046 297922 71102 297978
rect 97674 292294 97730 292350
rect 97798 292294 97854 292350
rect 97922 292294 97978 292350
rect 98046 292294 98102 292350
rect 97674 292170 97730 292226
rect 97798 292170 97854 292226
rect 97922 292170 97978 292226
rect 98046 292170 98102 292226
rect 97674 292046 97730 292102
rect 97798 292046 97854 292102
rect 97922 292046 97978 292102
rect 98046 292046 98102 292102
rect 97674 291922 97730 291978
rect 97798 291922 97854 291978
rect 97922 291922 97978 291978
rect 98046 291922 98102 291978
rect 70674 280294 70730 280350
rect 70798 280294 70854 280350
rect 70922 280294 70978 280350
rect 71046 280294 71102 280350
rect 70674 280170 70730 280226
rect 70798 280170 70854 280226
rect 70922 280170 70978 280226
rect 71046 280170 71102 280226
rect 70674 280046 70730 280102
rect 70798 280046 70854 280102
rect 70922 280046 70978 280102
rect 71046 280046 71102 280102
rect 70674 279922 70730 279978
rect 70798 279922 70854 279978
rect 70922 279922 70978 279978
rect 71046 279922 71102 279978
rect 66954 256294 67010 256350
rect 67078 256294 67134 256350
rect 67202 256294 67258 256350
rect 67326 256294 67382 256350
rect 66954 256170 67010 256226
rect 67078 256170 67134 256226
rect 67202 256170 67258 256226
rect 67326 256170 67382 256226
rect 66954 256046 67010 256102
rect 67078 256046 67134 256102
rect 67202 256046 67258 256102
rect 67326 256046 67382 256102
rect 66954 255922 67010 255978
rect 67078 255922 67134 255978
rect 67202 255922 67258 255978
rect 67326 255922 67382 255978
rect 36234 238294 36290 238350
rect 36358 238294 36414 238350
rect 36482 238294 36538 238350
rect 36606 238294 36662 238350
rect 36234 238170 36290 238226
rect 36358 238170 36414 238226
rect 36482 238170 36538 238226
rect 36606 238170 36662 238226
rect 36234 238046 36290 238102
rect 36358 238046 36414 238102
rect 36482 238046 36538 238102
rect 36606 238046 36662 238102
rect 36234 237922 36290 237978
rect 36358 237922 36414 237978
rect 36482 237922 36538 237978
rect 36606 237922 36662 237978
rect 36234 220294 36290 220350
rect 36358 220294 36414 220350
rect 36482 220294 36538 220350
rect 36606 220294 36662 220350
rect 36234 220170 36290 220226
rect 36358 220170 36414 220226
rect 36482 220170 36538 220226
rect 36606 220170 36662 220226
rect 36234 220046 36290 220102
rect 36358 220046 36414 220102
rect 36482 220046 36538 220102
rect 36606 220046 36662 220102
rect 36234 219922 36290 219978
rect 36358 219922 36414 219978
rect 36482 219922 36538 219978
rect 36606 219922 36662 219978
rect 9234 208294 9290 208350
rect 9358 208294 9414 208350
rect 9482 208294 9538 208350
rect 9606 208294 9662 208350
rect 9234 208170 9290 208226
rect 9358 208170 9414 208226
rect 9482 208170 9538 208226
rect 9606 208170 9662 208226
rect 9234 208046 9290 208102
rect 9358 208046 9414 208102
rect 9482 208046 9538 208102
rect 9606 208046 9662 208102
rect 9234 207922 9290 207978
rect 9358 207922 9414 207978
rect 9482 207922 9538 207978
rect 9606 207922 9662 207978
rect 18396 198996 18452 199018
rect 18396 198962 18452 198996
rect 24518 202294 24574 202350
rect 24642 202294 24698 202350
rect 24518 202170 24574 202226
rect 24642 202170 24698 202226
rect 24518 202046 24574 202102
rect 24642 202046 24698 202102
rect 24518 201922 24574 201978
rect 24642 201922 24698 201978
rect 70674 262294 70730 262350
rect 70798 262294 70854 262350
rect 70922 262294 70978 262350
rect 71046 262294 71102 262350
rect 70674 262170 70730 262226
rect 70798 262170 70854 262226
rect 70922 262170 70978 262226
rect 71046 262170 71102 262226
rect 70674 262046 70730 262102
rect 70798 262046 70854 262102
rect 70922 262046 70978 262102
rect 71046 262046 71102 262102
rect 70674 261922 70730 261978
rect 70798 261922 70854 261978
rect 70922 261922 70978 261978
rect 71046 261922 71102 261978
rect 80444 253502 80500 253558
rect 70674 244294 70730 244350
rect 70798 244294 70854 244350
rect 70922 244294 70978 244350
rect 71046 244294 71102 244350
rect 70674 244170 70730 244226
rect 70798 244170 70854 244226
rect 70922 244170 70978 244226
rect 71046 244170 71102 244226
rect 70674 244046 70730 244102
rect 70798 244046 70854 244102
rect 70922 244046 70978 244102
rect 71046 244046 71102 244102
rect 70674 243922 70730 243978
rect 70798 243922 70854 243978
rect 70922 243922 70978 243978
rect 71046 243922 71102 243978
rect 66954 238294 67010 238350
rect 67078 238294 67134 238350
rect 67202 238294 67258 238350
rect 67326 238294 67382 238350
rect 66954 238170 67010 238226
rect 67078 238170 67134 238226
rect 67202 238170 67258 238226
rect 67326 238170 67382 238226
rect 66954 238046 67010 238102
rect 67078 238046 67134 238102
rect 67202 238046 67258 238102
rect 67326 238046 67382 238102
rect 66954 237922 67010 237978
rect 67078 237922 67134 237978
rect 67202 237922 67258 237978
rect 67326 237922 67382 237978
rect 66954 220294 67010 220350
rect 67078 220294 67134 220350
rect 67202 220294 67258 220350
rect 67326 220294 67382 220350
rect 66954 220170 67010 220226
rect 67078 220170 67134 220226
rect 67202 220170 67258 220226
rect 67326 220170 67382 220226
rect 66954 220046 67010 220102
rect 67078 220046 67134 220102
rect 67202 220046 67258 220102
rect 67326 220046 67382 220102
rect 66954 219922 67010 219978
rect 67078 219922 67134 219978
rect 67202 219922 67258 219978
rect 67326 219922 67382 219978
rect 39878 208294 39934 208350
rect 40002 208294 40058 208350
rect 39878 208170 39934 208226
rect 40002 208170 40058 208226
rect 39878 208046 39934 208102
rect 40002 208046 40058 208102
rect 39878 207922 39934 207978
rect 40002 207922 40058 207978
rect 36234 202294 36290 202350
rect 36358 202294 36414 202350
rect 36482 202294 36538 202350
rect 36606 202294 36662 202350
rect 36234 202170 36290 202226
rect 36358 202170 36414 202226
rect 36482 202170 36538 202226
rect 36606 202170 36662 202226
rect 36234 202046 36290 202102
rect 36358 202046 36414 202102
rect 36482 202046 36538 202102
rect 36606 202046 36662 202102
rect 36234 201922 36290 201978
rect 36358 201922 36414 201978
rect 36482 201922 36538 201978
rect 36606 201922 36662 201978
rect 20636 195002 20692 195058
rect 20300 194102 20356 194158
rect 9234 190294 9290 190350
rect 9358 190294 9414 190350
rect 9482 190294 9538 190350
rect 9606 190294 9662 190350
rect 9234 190170 9290 190226
rect 9358 190170 9414 190226
rect 9482 190170 9538 190226
rect 9606 190170 9662 190226
rect 9234 190046 9290 190102
rect 9358 190046 9414 190102
rect 9482 190046 9538 190102
rect 9606 190046 9662 190102
rect 9234 189922 9290 189978
rect 9358 189922 9414 189978
rect 9482 189922 9538 189978
rect 9606 189922 9662 189978
rect 20076 186362 20132 186418
rect 24518 184294 24574 184350
rect 24642 184294 24698 184350
rect 24518 184170 24574 184226
rect 24642 184170 24698 184226
rect 24518 184046 24574 184102
rect 24642 184046 24698 184102
rect 24518 183922 24574 183978
rect 24642 183922 24698 183978
rect 55238 202294 55294 202350
rect 55362 202294 55418 202350
rect 55238 202170 55294 202226
rect 55362 202170 55418 202226
rect 55238 202046 55294 202102
rect 55362 202046 55418 202102
rect 55238 201922 55294 201978
rect 55362 201922 55418 201978
rect 64204 196622 64260 196678
rect 64204 195188 64260 195238
rect 64204 195182 64260 195188
rect 39878 190294 39934 190350
rect 40002 190294 40058 190350
rect 39878 190170 39934 190226
rect 40002 190170 40058 190226
rect 39878 190046 39934 190102
rect 40002 190046 40058 190102
rect 39878 189922 39934 189978
rect 40002 189922 40058 189978
rect 66954 202294 67010 202350
rect 67078 202294 67134 202350
rect 67202 202294 67258 202350
rect 67326 202294 67382 202350
rect 66954 202170 67010 202226
rect 67078 202170 67134 202226
rect 67202 202170 67258 202226
rect 67326 202170 67382 202226
rect 66954 202046 67010 202102
rect 67078 202046 67134 202102
rect 67202 202046 67258 202102
rect 67326 202046 67382 202102
rect 66954 201922 67010 201978
rect 67078 201922 67134 201978
rect 67202 201922 67258 201978
rect 67326 201922 67382 201978
rect 36234 184294 36290 184350
rect 36358 184294 36414 184350
rect 36482 184294 36538 184350
rect 36606 184294 36662 184350
rect 36234 184170 36290 184226
rect 36358 184170 36414 184226
rect 36482 184170 36538 184226
rect 36606 184170 36662 184226
rect 36234 184046 36290 184102
rect 36358 184046 36414 184102
rect 36482 184046 36538 184102
rect 36606 184046 36662 184102
rect 36234 183922 36290 183978
rect 36358 183922 36414 183978
rect 36482 183922 36538 183978
rect 36606 183922 36662 183978
rect 9234 172294 9290 172350
rect 9358 172294 9414 172350
rect 9482 172294 9538 172350
rect 9606 172294 9662 172350
rect 9234 172170 9290 172226
rect 9358 172170 9414 172226
rect 9482 172170 9538 172226
rect 9606 172170 9662 172226
rect 9234 172046 9290 172102
rect 9358 172046 9414 172102
rect 9482 172046 9538 172102
rect 9606 172046 9662 172102
rect 9234 171922 9290 171978
rect 9358 171922 9414 171978
rect 9482 171922 9538 171978
rect 9606 171922 9662 171978
rect 55238 184294 55294 184350
rect 55362 184294 55418 184350
rect 55238 184170 55294 184226
rect 55362 184170 55418 184226
rect 55238 184046 55294 184102
rect 55362 184046 55418 184102
rect 55238 183922 55294 183978
rect 55362 183922 55418 183978
rect 66954 184294 67010 184350
rect 67078 184294 67134 184350
rect 67202 184294 67258 184350
rect 67326 184294 67382 184350
rect 66954 184170 67010 184226
rect 67078 184170 67134 184226
rect 67202 184170 67258 184226
rect 67326 184170 67382 184226
rect 66954 184046 67010 184102
rect 67078 184046 67134 184102
rect 67202 184046 67258 184102
rect 67326 184046 67382 184102
rect 66954 183922 67010 183978
rect 67078 183922 67134 183978
rect 67202 183922 67258 183978
rect 67326 183922 67382 183978
rect 36234 166294 36290 166350
rect 36358 166294 36414 166350
rect 36482 166294 36538 166350
rect 36606 166294 36662 166350
rect 36234 166170 36290 166226
rect 36358 166170 36414 166226
rect 36482 166170 36538 166226
rect 36606 166170 36662 166226
rect 36234 166046 36290 166102
rect 36358 166046 36414 166102
rect 36482 166046 36538 166102
rect 36606 166046 36662 166102
rect 36234 165922 36290 165978
rect 36358 165922 36414 165978
rect 36482 165922 36538 165978
rect 36606 165922 36662 165978
rect 9234 154294 9290 154350
rect 9358 154294 9414 154350
rect 9482 154294 9538 154350
rect 9606 154294 9662 154350
rect 9234 154170 9290 154226
rect 9358 154170 9414 154226
rect 9482 154170 9538 154226
rect 9606 154170 9662 154226
rect 9234 154046 9290 154102
rect 9358 154046 9414 154102
rect 9482 154046 9538 154102
rect 9606 154046 9662 154102
rect 9234 153922 9290 153978
rect 9358 153922 9414 153978
rect 9482 153922 9538 153978
rect 9606 153922 9662 153978
rect 9234 136294 9290 136350
rect 9358 136294 9414 136350
rect 9482 136294 9538 136350
rect 9606 136294 9662 136350
rect 9234 136170 9290 136226
rect 9358 136170 9414 136226
rect 9482 136170 9538 136226
rect 9606 136170 9662 136226
rect 9234 136046 9290 136102
rect 9358 136046 9414 136102
rect 9482 136046 9538 136102
rect 9606 136046 9662 136102
rect 9234 135922 9290 135978
rect 9358 135922 9414 135978
rect 9482 135922 9538 135978
rect 9606 135922 9662 135978
rect 36234 148294 36290 148350
rect 36358 148294 36414 148350
rect 36482 148294 36538 148350
rect 36606 148294 36662 148350
rect 36234 148170 36290 148226
rect 36358 148170 36414 148226
rect 36482 148170 36538 148226
rect 36606 148170 36662 148226
rect 36234 148046 36290 148102
rect 36358 148046 36414 148102
rect 36482 148046 36538 148102
rect 36606 148046 36662 148102
rect 36234 147922 36290 147978
rect 36358 147922 36414 147978
rect 36482 147922 36538 147978
rect 36606 147922 36662 147978
rect 20076 131282 20132 131338
rect 18396 131102 18452 131158
rect 18284 128582 18340 128638
rect 24518 130294 24574 130350
rect 24642 130294 24698 130350
rect 24518 130170 24574 130226
rect 24642 130170 24698 130226
rect 24518 130046 24574 130102
rect 24642 130046 24698 130102
rect 24518 129922 24574 129978
rect 24642 129922 24698 129978
rect 39954 172294 40010 172350
rect 40078 172294 40134 172350
rect 40202 172294 40258 172350
rect 40326 172294 40382 172350
rect 39954 172170 40010 172226
rect 40078 172170 40134 172226
rect 40202 172170 40258 172226
rect 40326 172170 40382 172226
rect 39954 172046 40010 172102
rect 40078 172046 40134 172102
rect 40202 172046 40258 172102
rect 40326 172046 40382 172102
rect 39954 171922 40010 171978
rect 40078 171922 40134 171978
rect 40202 171922 40258 171978
rect 40326 171922 40382 171978
rect 66954 166294 67010 166350
rect 67078 166294 67134 166350
rect 67202 166294 67258 166350
rect 67326 166294 67382 166350
rect 66954 166170 67010 166226
rect 67078 166170 67134 166226
rect 67202 166170 67258 166226
rect 67326 166170 67382 166226
rect 66954 166046 67010 166102
rect 67078 166046 67134 166102
rect 67202 166046 67258 166102
rect 67326 166046 67382 166102
rect 66954 165922 67010 165978
rect 67078 165922 67134 165978
rect 67202 165922 67258 165978
rect 67326 165922 67382 165978
rect 39954 154294 40010 154350
rect 40078 154294 40134 154350
rect 40202 154294 40258 154350
rect 40326 154294 40382 154350
rect 39954 154170 40010 154226
rect 40078 154170 40134 154226
rect 40202 154170 40258 154226
rect 40326 154170 40382 154226
rect 39954 154046 40010 154102
rect 40078 154046 40134 154102
rect 40202 154046 40258 154102
rect 40326 154046 40382 154102
rect 39954 153922 40010 153978
rect 40078 153922 40134 153978
rect 40202 153922 40258 153978
rect 40326 153922 40382 153978
rect 39878 136294 39934 136350
rect 40002 136294 40058 136350
rect 39878 136170 39934 136226
rect 40002 136170 40058 136226
rect 39878 136046 39934 136102
rect 40002 136046 40058 136102
rect 39878 135922 39934 135978
rect 40002 135922 40058 135978
rect 36234 130294 36290 130350
rect 36358 130294 36414 130350
rect 36482 130294 36538 130350
rect 36606 130294 36662 130350
rect 36234 130170 36290 130226
rect 36358 130170 36414 130226
rect 36482 130170 36538 130226
rect 36606 130170 36662 130226
rect 36234 130046 36290 130102
rect 36358 130046 36414 130102
rect 36482 130046 36538 130102
rect 36606 130046 36662 130102
rect 36234 129922 36290 129978
rect 36358 129922 36414 129978
rect 36482 129922 36538 129978
rect 36606 129922 36662 129978
rect 55238 130294 55294 130350
rect 55362 130294 55418 130350
rect 55238 130170 55294 130226
rect 55362 130170 55418 130226
rect 55238 130046 55294 130102
rect 55362 130046 55418 130102
rect 55238 129922 55294 129978
rect 55362 129922 55418 129978
rect 20076 127862 20132 127918
rect 37772 127862 37828 127918
rect 20636 127502 20692 127558
rect 37772 127502 37828 127558
rect 64204 124262 64260 124318
rect 64204 120842 64260 120898
rect 9234 118294 9290 118350
rect 9358 118294 9414 118350
rect 9482 118294 9538 118350
rect 9606 118294 9662 118350
rect 9234 118170 9290 118226
rect 9358 118170 9414 118226
rect 9482 118170 9538 118226
rect 9606 118170 9662 118226
rect 9234 118046 9290 118102
rect 9358 118046 9414 118102
rect 9482 118046 9538 118102
rect 9606 118046 9662 118102
rect 9234 117922 9290 117978
rect 9358 117922 9414 117978
rect 9482 117922 9538 117978
rect 9606 117922 9662 117978
rect 39878 118294 39934 118350
rect 40002 118294 40058 118350
rect 39878 118170 39934 118226
rect 40002 118170 40058 118226
rect 39878 118046 39934 118102
rect 40002 118046 40058 118102
rect 39878 117922 39934 117978
rect 40002 117922 40058 117978
rect 66954 148294 67010 148350
rect 67078 148294 67134 148350
rect 67202 148294 67258 148350
rect 67326 148294 67382 148350
rect 66954 148170 67010 148226
rect 67078 148170 67134 148226
rect 67202 148170 67258 148226
rect 67326 148170 67382 148226
rect 66954 148046 67010 148102
rect 67078 148046 67134 148102
rect 67202 148046 67258 148102
rect 67326 148046 67382 148102
rect 66954 147922 67010 147978
rect 67078 147922 67134 147978
rect 67202 147922 67258 147978
rect 67326 147922 67382 147978
rect 86518 274294 86574 274350
rect 86642 274294 86698 274350
rect 86518 274170 86574 274226
rect 86642 274170 86698 274226
rect 86518 274046 86574 274102
rect 86642 274046 86698 274102
rect 86518 273922 86574 273978
rect 86642 273922 86698 273978
rect 128394 310294 128450 310350
rect 128518 310294 128574 310350
rect 128642 310294 128698 310350
rect 128766 310294 128822 310350
rect 128394 310170 128450 310226
rect 128518 310170 128574 310226
rect 128642 310170 128698 310226
rect 128766 310170 128822 310226
rect 128394 310046 128450 310102
rect 128518 310046 128574 310102
rect 128642 310046 128698 310102
rect 128766 310046 128822 310102
rect 128394 309922 128450 309978
rect 128518 309922 128574 309978
rect 128642 309922 128698 309978
rect 128766 309922 128822 309978
rect 128394 292294 128450 292350
rect 128518 292294 128574 292350
rect 128642 292294 128698 292350
rect 128766 292294 128822 292350
rect 128394 292170 128450 292226
rect 128518 292170 128574 292226
rect 128642 292170 128698 292226
rect 128766 292170 128822 292226
rect 128394 292046 128450 292102
rect 128518 292046 128574 292102
rect 128642 292046 128698 292102
rect 128766 292046 128822 292102
rect 128394 291922 128450 291978
rect 128518 291922 128574 291978
rect 128642 291922 128698 291978
rect 128766 291922 128822 291978
rect 101878 280294 101934 280350
rect 102002 280294 102058 280350
rect 101878 280170 101934 280226
rect 102002 280170 102058 280226
rect 101878 280046 101934 280102
rect 102002 280046 102058 280102
rect 101878 279922 101934 279978
rect 102002 279922 102058 279978
rect 126812 277982 126868 278038
rect 124348 275642 124404 275698
rect 97674 274294 97730 274350
rect 97798 274294 97854 274350
rect 97922 274294 97978 274350
rect 98046 274294 98102 274350
rect 97674 274170 97730 274226
rect 97798 274170 97854 274226
rect 97922 274170 97978 274226
rect 98046 274170 98102 274226
rect 97674 274046 97730 274102
rect 97798 274046 97854 274102
rect 97922 274046 97978 274102
rect 98046 274046 98102 274102
rect 97674 273922 97730 273978
rect 97798 273922 97854 273978
rect 97922 273922 97978 273978
rect 98046 273922 98102 273978
rect 82460 270602 82516 270658
rect 82460 267002 82516 267058
rect 82684 259442 82740 259498
rect 86518 256294 86574 256350
rect 86642 256294 86698 256350
rect 86518 256170 86574 256226
rect 86642 256170 86698 256226
rect 86518 256046 86574 256102
rect 86642 256046 86698 256102
rect 86518 255922 86574 255978
rect 86642 255922 86698 255978
rect 117238 274294 117294 274350
rect 117362 274294 117418 274350
rect 117238 274170 117294 274226
rect 117362 274170 117418 274226
rect 117238 274046 117294 274102
rect 117362 274046 117418 274102
rect 117238 273922 117294 273978
rect 117362 273922 117418 273978
rect 124348 268442 124404 268498
rect 127596 276362 127652 276418
rect 159114 364046 159170 364102
rect 159238 364046 159294 364102
rect 159362 364046 159418 364102
rect 159486 364046 159542 364102
rect 159114 363922 159170 363978
rect 159238 363922 159294 363978
rect 159362 363922 159418 363978
rect 159486 363922 159542 363978
rect 148518 346294 148574 346350
rect 148642 346294 148698 346350
rect 148518 346170 148574 346226
rect 148642 346170 148698 346226
rect 148518 346046 148574 346102
rect 148642 346046 148698 346102
rect 148518 345922 148574 345978
rect 148642 345922 148698 345978
rect 159114 346294 159170 346350
rect 159238 346294 159294 346350
rect 159362 346294 159418 346350
rect 159486 346294 159542 346350
rect 159114 346170 159170 346226
rect 159238 346170 159294 346226
rect 159362 346170 159418 346226
rect 159486 346170 159542 346226
rect 159114 346046 159170 346102
rect 159238 346046 159294 346102
rect 159362 346046 159418 346102
rect 159486 346046 159542 346102
rect 159114 345922 159170 345978
rect 159238 345922 159294 345978
rect 159362 345922 159418 345978
rect 159486 345922 159542 345978
rect 144060 341522 144116 341578
rect 141036 341162 141092 341218
rect 132114 334294 132170 334350
rect 132238 334294 132294 334350
rect 132362 334294 132418 334350
rect 132486 334294 132542 334350
rect 132114 334170 132170 334226
rect 132238 334170 132294 334226
rect 132362 334170 132418 334226
rect 132486 334170 132542 334226
rect 132114 334046 132170 334102
rect 132238 334046 132294 334102
rect 132362 334046 132418 334102
rect 132486 334046 132542 334102
rect 132114 333922 132170 333978
rect 132238 333922 132294 333978
rect 132362 333922 132418 333978
rect 132486 333922 132542 333978
rect 132114 316294 132170 316350
rect 132238 316294 132294 316350
rect 132362 316294 132418 316350
rect 132486 316294 132542 316350
rect 132114 316170 132170 316226
rect 132238 316170 132294 316226
rect 132362 316170 132418 316226
rect 132486 316170 132542 316226
rect 132114 316046 132170 316102
rect 132238 316046 132294 316102
rect 132362 316046 132418 316102
rect 132486 316046 132542 316102
rect 132114 315922 132170 315978
rect 132238 315922 132294 315978
rect 132362 315922 132418 315978
rect 132486 315922 132542 315978
rect 148518 328294 148574 328350
rect 148642 328294 148698 328350
rect 148518 328170 148574 328226
rect 148642 328170 148698 328226
rect 148518 328046 148574 328102
rect 148642 328046 148698 328102
rect 148518 327922 148574 327978
rect 148642 327922 148698 327978
rect 163878 460294 163934 460350
rect 164002 460294 164058 460350
rect 163878 460170 163934 460226
rect 164002 460170 164058 460226
rect 163878 460046 163934 460102
rect 164002 460046 164058 460102
rect 163878 459922 163934 459978
rect 164002 459922 164058 459978
rect 162834 442294 162890 442350
rect 162958 442294 163014 442350
rect 163082 442294 163138 442350
rect 163206 442294 163262 442350
rect 162834 442170 162890 442226
rect 162958 442170 163014 442226
rect 163082 442170 163138 442226
rect 163206 442170 163262 442226
rect 162834 442046 162890 442102
rect 162958 442046 163014 442102
rect 163082 442046 163138 442102
rect 163206 442046 163262 442102
rect 162834 441922 162890 441978
rect 162958 441922 163014 441978
rect 163082 441922 163138 441978
rect 163206 441922 163262 441978
rect 193554 598116 193610 598172
rect 193678 598116 193734 598172
rect 193802 598116 193858 598172
rect 193926 598116 193982 598172
rect 193554 597992 193610 598048
rect 193678 597992 193734 598048
rect 193802 597992 193858 598048
rect 193926 597992 193982 598048
rect 193554 597868 193610 597924
rect 193678 597868 193734 597924
rect 193802 597868 193858 597924
rect 193926 597868 193982 597924
rect 193554 597744 193610 597800
rect 193678 597744 193734 597800
rect 193802 597744 193858 597800
rect 193926 597744 193982 597800
rect 193554 586294 193610 586350
rect 193678 586294 193734 586350
rect 193802 586294 193858 586350
rect 193926 586294 193982 586350
rect 193554 586170 193610 586226
rect 193678 586170 193734 586226
rect 193802 586170 193858 586226
rect 193926 586170 193982 586226
rect 193554 586046 193610 586102
rect 193678 586046 193734 586102
rect 193802 586046 193858 586102
rect 193926 586046 193982 586102
rect 193554 585922 193610 585978
rect 193678 585922 193734 585978
rect 193802 585922 193858 585978
rect 193926 585922 193982 585978
rect 220554 597156 220610 597212
rect 220678 597156 220734 597212
rect 220802 597156 220858 597212
rect 220926 597156 220982 597212
rect 220554 597032 220610 597088
rect 220678 597032 220734 597088
rect 220802 597032 220858 597088
rect 220926 597032 220982 597088
rect 220554 596908 220610 596964
rect 220678 596908 220734 596964
rect 220802 596908 220858 596964
rect 220926 596908 220982 596964
rect 220554 596784 220610 596840
rect 220678 596784 220734 596840
rect 220802 596784 220858 596840
rect 220926 596784 220982 596840
rect 220554 580294 220610 580350
rect 220678 580294 220734 580350
rect 220802 580294 220858 580350
rect 220926 580294 220982 580350
rect 220554 580170 220610 580226
rect 220678 580170 220734 580226
rect 220802 580170 220858 580226
rect 220926 580170 220982 580226
rect 220554 580046 220610 580102
rect 220678 580046 220734 580102
rect 220802 580046 220858 580102
rect 220926 580046 220982 580102
rect 220554 579922 220610 579978
rect 220678 579922 220734 579978
rect 220802 579922 220858 579978
rect 220926 579922 220982 579978
rect 193554 568294 193610 568350
rect 193678 568294 193734 568350
rect 193802 568294 193858 568350
rect 193926 568294 193982 568350
rect 193554 568170 193610 568226
rect 193678 568170 193734 568226
rect 193802 568170 193858 568226
rect 193926 568170 193982 568226
rect 193554 568046 193610 568102
rect 193678 568046 193734 568102
rect 193802 568046 193858 568102
rect 193926 568046 193982 568102
rect 193554 567922 193610 567978
rect 193678 567922 193734 567978
rect 193802 567922 193858 567978
rect 193926 567922 193982 567978
rect 193554 550294 193610 550350
rect 193678 550294 193734 550350
rect 193802 550294 193858 550350
rect 193926 550294 193982 550350
rect 193554 550170 193610 550226
rect 193678 550170 193734 550226
rect 193802 550170 193858 550226
rect 193926 550170 193982 550226
rect 193554 550046 193610 550102
rect 193678 550046 193734 550102
rect 193802 550046 193858 550102
rect 193926 550046 193982 550102
rect 193554 549922 193610 549978
rect 193678 549922 193734 549978
rect 193802 549922 193858 549978
rect 193926 549922 193982 549978
rect 200844 571202 200900 571258
rect 193554 532294 193610 532350
rect 193678 532294 193734 532350
rect 193802 532294 193858 532350
rect 193926 532294 193982 532350
rect 193554 532170 193610 532226
rect 193678 532170 193734 532226
rect 193802 532170 193858 532226
rect 193926 532170 193982 532226
rect 193554 532046 193610 532102
rect 193678 532046 193734 532102
rect 193802 532046 193858 532102
rect 193926 532046 193982 532102
rect 193554 531922 193610 531978
rect 193678 531922 193734 531978
rect 193802 531922 193858 531978
rect 193926 531922 193982 531978
rect 193554 514294 193610 514350
rect 193678 514294 193734 514350
rect 193802 514294 193858 514350
rect 193926 514294 193982 514350
rect 193554 514170 193610 514226
rect 193678 514170 193734 514226
rect 193802 514170 193858 514226
rect 193926 514170 193982 514226
rect 193554 514046 193610 514102
rect 193678 514046 193734 514102
rect 193802 514046 193858 514102
rect 193926 514046 193982 514102
rect 193554 513922 193610 513978
rect 193678 513922 193734 513978
rect 193802 513922 193858 513978
rect 193926 513922 193982 513978
rect 193554 496294 193610 496350
rect 193678 496294 193734 496350
rect 193802 496294 193858 496350
rect 193926 496294 193982 496350
rect 193554 496170 193610 496226
rect 193678 496170 193734 496226
rect 193802 496170 193858 496226
rect 193926 496170 193982 496226
rect 193554 496046 193610 496102
rect 193678 496046 193734 496102
rect 193802 496046 193858 496102
rect 193926 496046 193982 496102
rect 193554 495922 193610 495978
rect 193678 495922 193734 495978
rect 193802 495922 193858 495978
rect 193926 495922 193982 495978
rect 193554 478294 193610 478350
rect 193678 478294 193734 478350
rect 193802 478294 193858 478350
rect 193926 478294 193982 478350
rect 193554 478170 193610 478226
rect 193678 478170 193734 478226
rect 193802 478170 193858 478226
rect 193926 478170 193982 478226
rect 193554 478046 193610 478102
rect 193678 478046 193734 478102
rect 193802 478046 193858 478102
rect 193926 478046 193982 478102
rect 193554 477922 193610 477978
rect 193678 477922 193734 477978
rect 193802 477922 193858 477978
rect 193926 477922 193982 477978
rect 193116 469502 193172 469558
rect 193116 465182 193172 465238
rect 189834 454294 189890 454350
rect 189958 454294 190014 454350
rect 190082 454294 190138 454350
rect 190206 454294 190262 454350
rect 189834 454170 189890 454226
rect 189958 454170 190014 454226
rect 190082 454170 190138 454226
rect 190206 454170 190262 454226
rect 189834 454046 189890 454102
rect 189958 454046 190014 454102
rect 190082 454046 190138 454102
rect 190206 454046 190262 454102
rect 189834 453922 189890 453978
rect 189958 453922 190014 453978
rect 190082 453922 190138 453978
rect 190206 453922 190262 453978
rect 189834 436294 189890 436350
rect 189958 436294 190014 436350
rect 190082 436294 190138 436350
rect 190206 436294 190262 436350
rect 189834 436170 189890 436226
rect 189958 436170 190014 436226
rect 190082 436170 190138 436226
rect 190206 436170 190262 436226
rect 189834 436046 189890 436102
rect 189958 436046 190014 436102
rect 190082 436046 190138 436102
rect 190206 436046 190262 436102
rect 189834 435922 189890 435978
rect 189958 435922 190014 435978
rect 190082 435922 190138 435978
rect 190206 435922 190262 435978
rect 162834 424294 162890 424350
rect 162958 424294 163014 424350
rect 163082 424294 163138 424350
rect 163206 424294 163262 424350
rect 162834 424170 162890 424226
rect 162958 424170 163014 424226
rect 163082 424170 163138 424226
rect 163206 424170 163262 424226
rect 162834 424046 162890 424102
rect 162958 424046 163014 424102
rect 163082 424046 163138 424102
rect 163206 424046 163262 424102
rect 162834 423922 162890 423978
rect 162958 423922 163014 423978
rect 163082 423922 163138 423978
rect 163206 423922 163262 423978
rect 179238 418294 179294 418350
rect 179362 418294 179418 418350
rect 179238 418170 179294 418226
rect 179362 418170 179418 418226
rect 179238 418046 179294 418102
rect 179362 418046 179418 418102
rect 179238 417922 179294 417978
rect 179362 417922 179418 417978
rect 189834 418294 189890 418350
rect 189958 418294 190014 418350
rect 190082 418294 190138 418350
rect 190206 418294 190262 418350
rect 189834 418170 189890 418226
rect 189958 418170 190014 418226
rect 190082 418170 190138 418226
rect 190206 418170 190262 418226
rect 189834 418046 189890 418102
rect 189958 418046 190014 418102
rect 190082 418046 190138 418102
rect 190206 418046 190262 418102
rect 189834 417922 189890 417978
rect 189958 417922 190014 417978
rect 190082 417922 190138 417978
rect 190206 417922 190262 417978
rect 162834 406294 162890 406350
rect 162958 406294 163014 406350
rect 163082 406294 163138 406350
rect 163206 406294 163262 406350
rect 162834 406170 162890 406226
rect 162958 406170 163014 406226
rect 163082 406170 163138 406226
rect 163206 406170 163262 406226
rect 162834 406046 162890 406102
rect 162958 406046 163014 406102
rect 163082 406046 163138 406102
rect 163206 406046 163262 406102
rect 162834 405922 162890 405978
rect 162958 405922 163014 405978
rect 163082 405922 163138 405978
rect 163206 405922 163262 405978
rect 163878 406294 163934 406350
rect 164002 406294 164058 406350
rect 163878 406170 163934 406226
rect 164002 406170 164058 406226
rect 163878 406046 163934 406102
rect 164002 406046 164058 406102
rect 163878 405922 163934 405978
rect 164002 405922 164058 405978
rect 179238 400294 179294 400350
rect 179362 400294 179418 400350
rect 179238 400170 179294 400226
rect 179362 400170 179418 400226
rect 179238 400046 179294 400102
rect 179362 400046 179418 400102
rect 179238 399922 179294 399978
rect 179362 399922 179418 399978
rect 189308 404702 189364 404758
rect 189420 403982 189476 404038
rect 189532 404522 189588 404578
rect 189532 399482 189588 399538
rect 197372 469502 197428 469558
rect 194908 467882 194964 467938
rect 199052 463562 199108 463618
rect 193554 460294 193610 460350
rect 193678 460294 193734 460350
rect 193802 460294 193858 460350
rect 193926 460294 193982 460350
rect 193554 460170 193610 460226
rect 193678 460170 193734 460226
rect 193802 460170 193858 460226
rect 193926 460170 193982 460226
rect 193554 460046 193610 460102
rect 193678 460046 193734 460102
rect 193802 460046 193858 460102
rect 193926 460046 193982 460102
rect 193554 459922 193610 459978
rect 193678 459922 193734 459978
rect 193802 459922 193858 459978
rect 193926 459922 193982 459978
rect 193554 442294 193610 442350
rect 193678 442294 193734 442350
rect 193802 442294 193858 442350
rect 193926 442294 193982 442350
rect 193554 442170 193610 442226
rect 193678 442170 193734 442226
rect 193802 442170 193858 442226
rect 193926 442170 193982 442226
rect 193554 442046 193610 442102
rect 193678 442046 193734 442102
rect 193802 442046 193858 442102
rect 193926 442046 193982 442102
rect 193554 441922 193610 441978
rect 193678 441922 193734 441978
rect 193802 441922 193858 441978
rect 193926 441922 193982 441978
rect 193554 424294 193610 424350
rect 193678 424294 193734 424350
rect 193802 424294 193858 424350
rect 193926 424294 193982 424350
rect 193554 424170 193610 424226
rect 193678 424170 193734 424226
rect 193802 424170 193858 424226
rect 193926 424170 193982 424226
rect 193554 424046 193610 424102
rect 193678 424046 193734 424102
rect 193802 424046 193858 424102
rect 193926 424046 193982 424102
rect 193554 423922 193610 423978
rect 193678 423922 193734 423978
rect 193802 423922 193858 423978
rect 193926 423922 193982 423978
rect 191548 406862 191604 406918
rect 193554 406294 193610 406350
rect 193678 406294 193734 406350
rect 193802 406294 193858 406350
rect 193926 406294 193982 406350
rect 193554 406170 193610 406226
rect 193678 406170 193734 406226
rect 193802 406170 193858 406226
rect 193926 406170 193982 406226
rect 193554 406046 193610 406102
rect 193678 406046 193734 406102
rect 193802 406046 193858 406102
rect 193926 406046 193982 406102
rect 193554 405922 193610 405978
rect 193678 405922 193734 405978
rect 193802 405922 193858 405978
rect 193926 405922 193982 405978
rect 189834 400294 189890 400350
rect 189958 400294 190014 400350
rect 190082 400294 190138 400350
rect 190206 400294 190262 400350
rect 189834 400170 189890 400226
rect 189958 400170 190014 400226
rect 190082 400170 190138 400226
rect 190206 400170 190262 400226
rect 189834 400046 189890 400102
rect 189958 400046 190014 400102
rect 190082 400046 190138 400102
rect 190206 400046 190262 400102
rect 189834 399922 189890 399978
rect 189958 399922 190014 399978
rect 190082 399922 190138 399978
rect 190206 399922 190262 399978
rect 162834 388294 162890 388350
rect 162958 388294 163014 388350
rect 163082 388294 163138 388350
rect 163206 388294 163262 388350
rect 163836 388333 163892 388389
rect 163940 388333 163996 388389
rect 164044 388333 164100 388389
rect 162834 388170 162890 388226
rect 162958 388170 163014 388226
rect 163082 388170 163138 388226
rect 163206 388170 163262 388226
rect 162834 388046 162890 388102
rect 162958 388046 163014 388102
rect 163082 388046 163138 388102
rect 163206 388046 163262 388102
rect 162834 387922 162890 387978
rect 162958 387922 163014 387978
rect 163082 387922 163138 387978
rect 163206 387922 163262 387978
rect 162834 370294 162890 370350
rect 162958 370294 163014 370350
rect 163082 370294 163138 370350
rect 163206 370294 163262 370350
rect 162834 370170 162890 370226
rect 162958 370170 163014 370226
rect 163082 370170 163138 370226
rect 163206 370170 163262 370226
rect 162834 370046 162890 370102
rect 162958 370046 163014 370102
rect 163082 370046 163138 370102
rect 163206 370046 163262 370102
rect 162834 369922 162890 369978
rect 162958 369922 163014 369978
rect 163082 369922 163138 369978
rect 163206 369922 163262 369978
rect 189834 382294 189890 382350
rect 189958 382294 190014 382350
rect 190082 382294 190138 382350
rect 190206 382294 190262 382350
rect 189834 382170 189890 382226
rect 189958 382170 190014 382226
rect 190082 382170 190138 382226
rect 190206 382170 190262 382226
rect 189834 382046 189890 382102
rect 189958 382046 190014 382102
rect 190082 382046 190138 382102
rect 190206 382046 190262 382102
rect 189834 381922 189890 381978
rect 189958 381922 190014 381978
rect 190082 381922 190138 381978
rect 190206 381922 190262 381978
rect 199836 403082 199892 403138
rect 199052 402362 199108 402418
rect 199052 396242 199108 396298
rect 193554 388294 193610 388350
rect 193678 388294 193734 388350
rect 193802 388294 193858 388350
rect 193926 388294 193982 388350
rect 193554 388170 193610 388226
rect 193678 388170 193734 388226
rect 193802 388170 193858 388226
rect 193926 388170 193982 388226
rect 193554 388046 193610 388102
rect 193678 388046 193734 388102
rect 193802 388046 193858 388102
rect 193926 388046 193982 388102
rect 193554 387922 193610 387978
rect 193678 387922 193734 387978
rect 193802 387922 193858 387978
rect 193926 387922 193982 387978
rect 189834 364294 189890 364350
rect 189958 364294 190014 364350
rect 190082 364294 190138 364350
rect 190206 364294 190262 364350
rect 189834 364170 189890 364226
rect 189958 364170 190014 364226
rect 190082 364170 190138 364226
rect 190206 364170 190262 364226
rect 189834 364046 189890 364102
rect 189958 364046 190014 364102
rect 190082 364046 190138 364102
rect 190206 364046 190262 364102
rect 189834 363922 189890 363978
rect 189958 363922 190014 363978
rect 190082 363922 190138 363978
rect 190206 363922 190262 363978
rect 162834 352294 162890 352350
rect 162958 352294 163014 352350
rect 163082 352294 163138 352350
rect 163206 352294 163262 352350
rect 162834 352170 162890 352226
rect 162958 352170 163014 352226
rect 163082 352170 163138 352226
rect 163206 352170 163262 352226
rect 162834 352046 162890 352102
rect 162958 352046 163014 352102
rect 163082 352046 163138 352102
rect 163206 352046 163262 352102
rect 162834 351922 162890 351978
rect 162958 351922 163014 351978
rect 163082 351922 163138 351978
rect 163206 351922 163262 351978
rect 160524 342782 160580 342838
rect 159740 341522 159796 341578
rect 159740 339182 159796 339238
rect 163878 352294 163934 352350
rect 164002 352294 164058 352350
rect 163878 352170 163934 352226
rect 164002 352170 164058 352226
rect 163878 352046 163934 352102
rect 164002 352046 164058 352102
rect 163878 351922 163934 351978
rect 164002 351922 164058 351978
rect 179238 346294 179294 346350
rect 179362 346294 179418 346350
rect 179238 346170 179294 346226
rect 179362 346170 179418 346226
rect 179238 346046 179294 346102
rect 179362 346046 179418 346102
rect 179238 345922 179294 345978
rect 179362 345922 179418 345978
rect 189834 346294 189890 346350
rect 189958 346294 190014 346350
rect 190082 346294 190138 346350
rect 190206 346294 190262 346350
rect 189834 346170 189890 346226
rect 189958 346170 190014 346226
rect 190082 346170 190138 346226
rect 190206 346170 190262 346226
rect 189834 346046 189890 346102
rect 189958 346046 190014 346102
rect 190082 346046 190138 346102
rect 190206 346046 190262 346102
rect 189834 345922 189890 345978
rect 189958 345922 190014 345978
rect 190082 345922 190138 345978
rect 190206 345922 190262 345978
rect 189084 343502 189140 343558
rect 160524 337562 160580 337618
rect 159114 328294 159170 328350
rect 159238 328294 159294 328350
rect 159362 328294 159418 328350
rect 159486 328294 159542 328350
rect 159114 328170 159170 328226
rect 159238 328170 159294 328226
rect 159362 328170 159418 328226
rect 159486 328170 159542 328226
rect 159114 328046 159170 328102
rect 159238 328046 159294 328102
rect 159362 328046 159418 328102
rect 159486 328046 159542 328102
rect 159114 327922 159170 327978
rect 159238 327922 159294 327978
rect 159362 327922 159418 327978
rect 159486 327922 159542 327978
rect 160412 336122 160468 336178
rect 163878 334294 163934 334350
rect 164002 334294 164058 334350
rect 163878 334170 163934 334226
rect 164002 334170 164058 334226
rect 163878 334046 163934 334102
rect 164002 334046 164058 334102
rect 163878 333922 163934 333978
rect 164002 333922 164058 333978
rect 160412 325862 160468 325918
rect 160524 332702 160580 332758
rect 162540 331802 162596 331858
rect 162540 330542 162596 330598
rect 166236 331082 166292 331138
rect 166236 330362 166292 330418
rect 160524 325682 160580 325738
rect 179238 328294 179294 328350
rect 179362 328294 179418 328350
rect 179238 328170 179294 328226
rect 179362 328170 179418 328226
rect 179238 328046 179294 328102
rect 179362 328046 179418 328102
rect 179238 327922 179294 327978
rect 179362 327922 179418 327978
rect 189420 338462 189476 338518
rect 193554 370294 193610 370350
rect 193678 370294 193734 370350
rect 193802 370294 193858 370350
rect 193926 370294 193982 370350
rect 193554 370170 193610 370226
rect 193678 370170 193734 370226
rect 193802 370170 193858 370226
rect 193926 370170 193982 370226
rect 193554 370046 193610 370102
rect 193678 370046 193734 370102
rect 193802 370046 193858 370102
rect 193926 370046 193982 370102
rect 193554 369922 193610 369978
rect 193678 369922 193734 369978
rect 193802 369922 193858 369978
rect 193926 369922 193982 369978
rect 193554 352294 193610 352350
rect 193678 352294 193734 352350
rect 193802 352294 193858 352350
rect 193926 352294 193982 352350
rect 193554 352170 193610 352226
rect 193678 352170 193734 352226
rect 193802 352170 193858 352226
rect 193926 352170 193982 352226
rect 193554 352046 193610 352102
rect 193678 352046 193734 352102
rect 193802 352046 193858 352102
rect 193926 352046 193982 352102
rect 193554 351922 193610 351978
rect 193678 351922 193734 351978
rect 193802 351922 193858 351978
rect 193926 351922 193982 351978
rect 192444 344402 192500 344458
rect 192332 341702 192388 341758
rect 197372 347822 197428 347878
rect 195692 344582 195748 344638
rect 195804 342962 195860 343018
rect 193554 334294 193610 334350
rect 193678 334294 193734 334350
rect 193802 334294 193858 334350
rect 193926 334294 193982 334350
rect 193554 334170 193610 334226
rect 193678 334170 193734 334226
rect 193802 334170 193858 334226
rect 193926 334170 193982 334226
rect 193554 334046 193610 334102
rect 193678 334046 193734 334102
rect 193802 334046 193858 334102
rect 193926 334046 193982 334102
rect 193554 333922 193610 333978
rect 193678 333922 193734 333978
rect 193802 333922 193858 333978
rect 193926 333922 193982 333978
rect 189834 328294 189890 328350
rect 189958 328294 190014 328350
rect 190082 328294 190138 328350
rect 190206 328294 190262 328350
rect 189834 328170 189890 328226
rect 189958 328170 190014 328226
rect 190082 328170 190138 328226
rect 190206 328170 190262 328226
rect 189834 328046 189890 328102
rect 189958 328046 190014 328102
rect 190082 328046 190138 328102
rect 190206 328046 190262 328102
rect 189834 327922 189890 327978
rect 189958 327922 190014 327978
rect 190082 327922 190138 327978
rect 190206 327922 190262 327978
rect 162834 316294 162890 316350
rect 162958 316294 163014 316350
rect 163082 316294 163138 316350
rect 163206 316294 163262 316350
rect 162834 316170 162890 316226
rect 162958 316170 163014 316226
rect 163082 316170 163138 316226
rect 163206 316170 163262 316226
rect 162834 316046 162890 316102
rect 162958 316046 163014 316102
rect 163082 316046 163138 316102
rect 163206 316046 163262 316102
rect 162834 315922 162890 315978
rect 162958 315922 163014 315978
rect 163082 315922 163138 315978
rect 163206 315922 163262 315978
rect 159114 310294 159170 310350
rect 159238 310294 159294 310350
rect 159362 310294 159418 310350
rect 159486 310294 159542 310350
rect 159114 310170 159170 310226
rect 159238 310170 159294 310226
rect 159362 310170 159418 310226
rect 159486 310170 159542 310226
rect 159114 310046 159170 310102
rect 159238 310046 159294 310102
rect 159362 310046 159418 310102
rect 159486 310046 159542 310102
rect 159114 309922 159170 309978
rect 159238 309922 159294 309978
rect 159362 309922 159418 309978
rect 159486 309922 159542 309978
rect 132114 298294 132170 298350
rect 132238 298294 132294 298350
rect 132362 298294 132418 298350
rect 132486 298294 132542 298350
rect 132114 298170 132170 298226
rect 132238 298170 132294 298226
rect 132362 298170 132418 298226
rect 132486 298170 132542 298226
rect 132114 298046 132170 298102
rect 132238 298046 132294 298102
rect 132362 298046 132418 298102
rect 132486 298046 132542 298102
rect 132114 297922 132170 297978
rect 132238 297922 132294 297978
rect 132362 297922 132418 297978
rect 132486 297922 132542 297978
rect 128394 274294 128450 274350
rect 128518 274294 128574 274350
rect 128642 274294 128698 274350
rect 128766 274294 128822 274350
rect 128394 274170 128450 274226
rect 128518 274170 128574 274226
rect 128642 274170 128698 274226
rect 128766 274170 128822 274226
rect 128394 274046 128450 274102
rect 128518 274046 128574 274102
rect 128642 274046 128698 274102
rect 128766 274046 128822 274102
rect 128394 273922 128450 273978
rect 128518 273922 128574 273978
rect 128642 273922 128698 273978
rect 128766 273922 128822 273978
rect 127596 272942 127652 272998
rect 101878 262294 101934 262350
rect 102002 262294 102058 262350
rect 101878 262170 101934 262226
rect 102002 262170 102058 262226
rect 101878 262046 101934 262102
rect 102002 262046 102058 262102
rect 101878 261922 101934 261978
rect 102002 261922 102058 261978
rect 125132 259442 125188 259498
rect 97674 256294 97730 256350
rect 97798 256294 97854 256350
rect 97922 256294 97978 256350
rect 98046 256294 98102 256350
rect 97674 256170 97730 256226
rect 97798 256170 97854 256226
rect 97922 256170 97978 256226
rect 98046 256170 98102 256226
rect 97674 256046 97730 256102
rect 97798 256046 97854 256102
rect 97922 256046 97978 256102
rect 98046 256046 98102 256102
rect 97674 255922 97730 255978
rect 97798 255922 97854 255978
rect 97922 255922 97978 255978
rect 98046 255922 98102 255978
rect 70674 226294 70730 226350
rect 70798 226294 70854 226350
rect 70922 226294 70978 226350
rect 71046 226294 71102 226350
rect 70674 226170 70730 226226
rect 70798 226170 70854 226226
rect 70922 226170 70978 226226
rect 71046 226170 71102 226226
rect 70674 226046 70730 226102
rect 70798 226046 70854 226102
rect 70922 226046 70978 226102
rect 71046 226046 71102 226102
rect 70674 225922 70730 225978
rect 70798 225922 70854 225978
rect 70922 225922 70978 225978
rect 71046 225922 71102 225978
rect 117238 256294 117294 256350
rect 117362 256294 117418 256350
rect 117238 256170 117294 256226
rect 117362 256170 117418 256226
rect 117238 256046 117294 256102
rect 117362 256046 117418 256102
rect 117238 255922 117294 255978
rect 117362 255922 117418 255978
rect 126812 254402 126868 254458
rect 128394 256294 128450 256350
rect 128518 256294 128574 256350
rect 128642 256294 128698 256350
rect 128766 256294 128822 256350
rect 128394 256170 128450 256226
rect 128518 256170 128574 256226
rect 128642 256170 128698 256226
rect 128766 256170 128822 256226
rect 128394 256046 128450 256102
rect 128518 256046 128574 256102
rect 128642 256046 128698 256102
rect 128766 256046 128822 256102
rect 128394 255922 128450 255978
rect 128518 255922 128574 255978
rect 128642 255922 128698 255978
rect 128766 255922 128822 255978
rect 125132 253322 125188 253378
rect 97674 238294 97730 238350
rect 97798 238294 97854 238350
rect 97922 238294 97978 238350
rect 98046 238294 98102 238350
rect 97674 238170 97730 238226
rect 97798 238170 97854 238226
rect 97922 238170 97978 238226
rect 98046 238170 98102 238226
rect 97674 238046 97730 238102
rect 97798 238046 97854 238102
rect 97922 238046 97978 238102
rect 98046 238046 98102 238102
rect 97674 237922 97730 237978
rect 97798 237922 97854 237978
rect 97922 237922 97978 237978
rect 98046 237922 98102 237978
rect 70674 208294 70730 208350
rect 70798 208294 70854 208350
rect 70922 208294 70978 208350
rect 71046 208294 71102 208350
rect 70674 208170 70730 208226
rect 70798 208170 70854 208226
rect 70922 208170 70978 208226
rect 71046 208170 71102 208226
rect 70674 208046 70730 208102
rect 70798 208046 70854 208102
rect 70922 208046 70978 208102
rect 71046 208046 71102 208102
rect 70674 207922 70730 207978
rect 70798 207922 70854 207978
rect 70922 207922 70978 207978
rect 71046 207922 71102 207978
rect 70674 190294 70730 190350
rect 70798 190294 70854 190350
rect 70922 190294 70978 190350
rect 71046 190294 71102 190350
rect 70674 190170 70730 190226
rect 70798 190170 70854 190226
rect 70922 190170 70978 190226
rect 71046 190170 71102 190226
rect 70674 190046 70730 190102
rect 70798 190046 70854 190102
rect 70922 190046 70978 190102
rect 71046 190046 71102 190102
rect 70674 189922 70730 189978
rect 70798 189922 70854 189978
rect 70922 189922 70978 189978
rect 71046 189922 71102 189978
rect 159114 292294 159170 292350
rect 159238 292294 159294 292350
rect 159362 292294 159418 292350
rect 159486 292294 159542 292350
rect 159114 292170 159170 292226
rect 159238 292170 159294 292226
rect 159362 292170 159418 292226
rect 159486 292170 159542 292226
rect 159114 292046 159170 292102
rect 159238 292046 159294 292102
rect 159362 292046 159418 292102
rect 159486 292046 159542 292102
rect 159114 291922 159170 291978
rect 159238 291922 159294 291978
rect 159362 291922 159418 291978
rect 159486 291922 159542 291978
rect 132114 280294 132170 280350
rect 132238 280294 132294 280350
rect 132362 280294 132418 280350
rect 132486 280294 132542 280350
rect 132114 280170 132170 280226
rect 132238 280170 132294 280226
rect 132362 280170 132418 280226
rect 132486 280170 132542 280226
rect 132114 280046 132170 280102
rect 132238 280046 132294 280102
rect 132362 280046 132418 280102
rect 132486 280046 132542 280102
rect 132114 279922 132170 279978
rect 132238 279922 132294 279978
rect 132362 279922 132418 279978
rect 132486 279922 132542 279978
rect 130172 250262 130228 250318
rect 133532 275642 133588 275698
rect 132114 262294 132170 262350
rect 132238 262294 132294 262350
rect 132362 262294 132418 262350
rect 132486 262294 132542 262350
rect 132114 262170 132170 262226
rect 132238 262170 132294 262226
rect 132362 262170 132418 262226
rect 132486 262170 132542 262226
rect 132114 262046 132170 262102
rect 132238 262046 132294 262102
rect 132362 262046 132418 262102
rect 132486 262046 132542 262102
rect 132114 261922 132170 261978
rect 132238 261922 132294 261978
rect 132362 261922 132418 261978
rect 132486 261922 132542 261978
rect 128394 238294 128450 238350
rect 128518 238294 128574 238350
rect 128642 238294 128698 238350
rect 128766 238294 128822 238350
rect 128394 238170 128450 238226
rect 128518 238170 128574 238226
rect 128642 238170 128698 238226
rect 128766 238170 128822 238226
rect 128394 238046 128450 238102
rect 128518 238046 128574 238102
rect 128642 238046 128698 238102
rect 128766 238046 128822 238102
rect 128394 237922 128450 237978
rect 128518 237922 128574 237978
rect 128642 237922 128698 237978
rect 128766 237922 128822 237978
rect 97674 220294 97730 220350
rect 97798 220294 97854 220350
rect 97922 220294 97978 220350
rect 98046 220294 98102 220350
rect 97674 220170 97730 220226
rect 97798 220170 97854 220226
rect 97922 220170 97978 220226
rect 98046 220170 98102 220226
rect 97674 220046 97730 220102
rect 97798 220046 97854 220102
rect 97922 220046 97978 220102
rect 98046 220046 98102 220102
rect 97674 219922 97730 219978
rect 97798 219922 97854 219978
rect 97922 219922 97978 219978
rect 98046 219922 98102 219978
rect 86518 202294 86574 202350
rect 86642 202294 86698 202350
rect 86518 202170 86574 202226
rect 86642 202170 86698 202226
rect 86518 202046 86574 202102
rect 86642 202046 86698 202102
rect 86518 201922 86574 201978
rect 86642 201922 86698 201978
rect 101878 208294 101934 208350
rect 102002 208294 102058 208350
rect 101878 208170 101934 208226
rect 102002 208170 102058 208226
rect 101878 208046 101934 208102
rect 102002 208046 102058 208102
rect 101878 207922 101934 207978
rect 102002 207922 102058 207978
rect 97674 202294 97730 202350
rect 97798 202294 97854 202350
rect 97922 202294 97978 202350
rect 98046 202294 98102 202350
rect 97674 202170 97730 202226
rect 97798 202170 97854 202226
rect 97922 202170 97978 202226
rect 98046 202170 98102 202226
rect 97674 202046 97730 202102
rect 97798 202046 97854 202102
rect 97922 202046 97978 202102
rect 98046 202046 98102 202102
rect 97674 201922 97730 201978
rect 97798 201922 97854 201978
rect 97922 201922 97978 201978
rect 98046 201922 98102 201978
rect 82684 198962 82740 199018
rect 82684 186002 82740 186058
rect 86518 184294 86574 184350
rect 86642 184294 86698 184350
rect 86518 184170 86574 184226
rect 86642 184170 86698 184226
rect 86518 184046 86574 184102
rect 86642 184046 86698 184102
rect 86518 183922 86574 183978
rect 86642 183922 86698 183978
rect 117238 202294 117294 202350
rect 117362 202294 117418 202350
rect 117238 202170 117294 202226
rect 117362 202170 117418 202226
rect 117238 202046 117294 202102
rect 117362 202046 117418 202102
rect 117238 201922 117294 201978
rect 117362 201922 117418 201978
rect 101878 190294 101934 190350
rect 102002 190294 102058 190350
rect 101878 190170 101934 190226
rect 102002 190170 102058 190226
rect 101878 190046 101934 190102
rect 102002 190046 102058 190102
rect 101878 189922 101934 189978
rect 102002 189922 102058 189978
rect 141036 270602 141092 270658
rect 141036 264662 141092 264718
rect 148518 274294 148574 274350
rect 148642 274294 148698 274350
rect 148518 274170 148574 274226
rect 148642 274170 148698 274226
rect 148518 274046 148574 274102
rect 148642 274046 148698 274102
rect 148518 273922 148574 273978
rect 148642 273922 148698 273978
rect 159114 274294 159170 274350
rect 159238 274294 159294 274350
rect 159362 274294 159418 274350
rect 159486 274294 159542 274350
rect 159114 274170 159170 274226
rect 159238 274170 159294 274226
rect 159362 274170 159418 274226
rect 159486 274170 159542 274226
rect 159114 274046 159170 274102
rect 159238 274046 159294 274102
rect 159362 274046 159418 274102
rect 159486 274046 159542 274102
rect 159114 273922 159170 273978
rect 159238 273922 159294 273978
rect 159362 273922 159418 273978
rect 159486 273922 159542 273978
rect 144060 271142 144116 271198
rect 144284 260342 144340 260398
rect 142716 258542 142772 258598
rect 148518 256294 148574 256350
rect 148642 256294 148698 256350
rect 148518 256170 148574 256226
rect 148642 256170 148698 256226
rect 148518 256046 148574 256102
rect 148642 256046 148698 256102
rect 148518 255922 148574 255978
rect 148642 255922 148698 255978
rect 162834 298294 162890 298350
rect 162958 298294 163014 298350
rect 163082 298294 163138 298350
rect 163206 298294 163262 298350
rect 162834 298170 162890 298226
rect 162958 298170 163014 298226
rect 163082 298170 163138 298226
rect 163206 298170 163262 298226
rect 162834 298046 162890 298102
rect 162958 298046 163014 298102
rect 163082 298046 163138 298102
rect 163206 298046 163262 298102
rect 162834 297922 162890 297978
rect 162958 297922 163014 297978
rect 163082 297922 163138 297978
rect 163206 297922 163262 297978
rect 189834 310294 189890 310350
rect 189958 310294 190014 310350
rect 190082 310294 190138 310350
rect 190206 310294 190262 310350
rect 189834 310170 189890 310226
rect 189958 310170 190014 310226
rect 190082 310170 190138 310226
rect 190206 310170 190262 310226
rect 189834 310046 189890 310102
rect 189958 310046 190014 310102
rect 190082 310046 190138 310102
rect 190206 310046 190262 310102
rect 189834 309922 189890 309978
rect 189958 309922 190014 309978
rect 190082 309922 190138 309978
rect 190206 309922 190262 309978
rect 189834 292294 189890 292350
rect 189958 292294 190014 292350
rect 190082 292294 190138 292350
rect 190206 292294 190262 292350
rect 189834 292170 189890 292226
rect 189958 292170 190014 292226
rect 190082 292170 190138 292226
rect 190206 292170 190262 292226
rect 189834 292046 189890 292102
rect 189958 292046 190014 292102
rect 190082 292046 190138 292102
rect 190206 292046 190262 292102
rect 189834 291922 189890 291978
rect 189958 291922 190014 291978
rect 190082 291922 190138 291978
rect 190206 291922 190262 291978
rect 162834 280294 162890 280350
rect 162958 280294 163014 280350
rect 163082 280294 163138 280350
rect 163206 280294 163262 280350
rect 162834 280170 162890 280226
rect 162958 280170 163014 280226
rect 163082 280170 163138 280226
rect 163206 280170 163262 280226
rect 162834 280046 162890 280102
rect 162958 280046 163014 280102
rect 163082 280046 163138 280102
rect 163206 280046 163262 280102
rect 162834 279922 162890 279978
rect 162958 279922 163014 279978
rect 163082 279922 163138 279978
rect 163206 279922 163262 279978
rect 163878 280294 163934 280350
rect 164002 280294 164058 280350
rect 163878 280170 163934 280226
rect 164002 280170 164058 280226
rect 163878 280046 163934 280102
rect 164002 280046 164058 280102
rect 163878 279922 163934 279978
rect 164002 279922 164058 279978
rect 179238 274294 179294 274350
rect 179362 274294 179418 274350
rect 179238 274170 179294 274226
rect 179362 274170 179418 274226
rect 179238 274046 179294 274102
rect 179362 274046 179418 274102
rect 179238 273922 179294 273978
rect 179362 273922 179418 273978
rect 163878 262294 163934 262350
rect 164002 262294 164058 262350
rect 163878 262170 163934 262226
rect 164002 262170 164058 262226
rect 159114 256294 159170 256350
rect 159238 256294 159294 256350
rect 159362 256294 159418 256350
rect 159486 256294 159542 256350
rect 159114 256170 159170 256226
rect 159238 256170 159294 256226
rect 159362 256170 159418 256226
rect 159486 256170 159542 256226
rect 159114 256046 159170 256102
rect 159238 256046 159294 256102
rect 159362 256046 159418 256102
rect 159486 256046 159542 256102
rect 159114 255922 159170 255978
rect 159238 255922 159294 255978
rect 159362 255922 159418 255978
rect 159486 255922 159542 255978
rect 135212 255302 135268 255358
rect 133532 251882 133588 251938
rect 132114 244294 132170 244350
rect 132238 244294 132294 244350
rect 132362 244294 132418 244350
rect 132486 244294 132542 244350
rect 132114 244170 132170 244226
rect 132238 244170 132294 244226
rect 132362 244170 132418 244226
rect 132486 244170 132542 244226
rect 132114 244046 132170 244102
rect 132238 244046 132294 244102
rect 132362 244046 132418 244102
rect 132486 244046 132542 244102
rect 132114 243922 132170 243978
rect 132238 243922 132294 243978
rect 132362 243922 132418 243978
rect 132486 243922 132542 243978
rect 159114 238294 159170 238350
rect 159238 238294 159294 238350
rect 159362 238294 159418 238350
rect 159486 238294 159542 238350
rect 159114 238170 159170 238226
rect 159238 238170 159294 238226
rect 159362 238170 159418 238226
rect 159486 238170 159542 238226
rect 159114 238046 159170 238102
rect 159238 238046 159294 238102
rect 159362 238046 159418 238102
rect 159486 238046 159542 238102
rect 159114 237922 159170 237978
rect 159238 237922 159294 237978
rect 159362 237922 159418 237978
rect 159486 237922 159542 237978
rect 132114 226294 132170 226350
rect 132238 226294 132294 226350
rect 132362 226294 132418 226350
rect 132486 226294 132542 226350
rect 132114 226170 132170 226226
rect 132238 226170 132294 226226
rect 132362 226170 132418 226226
rect 132486 226170 132542 226226
rect 132114 226046 132170 226102
rect 132238 226046 132294 226102
rect 132362 226046 132418 226102
rect 132486 226046 132542 226102
rect 132114 225922 132170 225978
rect 132238 225922 132294 225978
rect 132362 225922 132418 225978
rect 132486 225922 132542 225978
rect 128394 220294 128450 220350
rect 128518 220294 128574 220350
rect 128642 220294 128698 220350
rect 128766 220294 128822 220350
rect 128394 220170 128450 220226
rect 128518 220170 128574 220226
rect 128642 220170 128698 220226
rect 128766 220170 128822 220226
rect 128394 220046 128450 220102
rect 128518 220046 128574 220102
rect 128642 220046 128698 220102
rect 128766 220046 128822 220102
rect 128394 219922 128450 219978
rect 128518 219922 128574 219978
rect 128642 219922 128698 219978
rect 128766 219922 128822 219978
rect 128394 202294 128450 202350
rect 128518 202294 128574 202350
rect 128642 202294 128698 202350
rect 128766 202294 128822 202350
rect 128394 202170 128450 202226
rect 128518 202170 128574 202226
rect 128642 202170 128698 202226
rect 128766 202170 128822 202226
rect 128394 202046 128450 202102
rect 128518 202046 128574 202102
rect 128642 202046 128698 202102
rect 128766 202046 128822 202102
rect 128394 201922 128450 201978
rect 128518 201922 128574 201978
rect 128642 201922 128698 201978
rect 128766 201922 128822 201978
rect 127484 193922 127540 193978
rect 127596 193202 127652 193258
rect 127596 186182 127652 186238
rect 97674 184294 97730 184350
rect 97798 184294 97854 184350
rect 97922 184294 97978 184350
rect 98046 184294 98102 184350
rect 97674 184170 97730 184226
rect 97798 184170 97854 184226
rect 97922 184170 97978 184226
rect 98046 184170 98102 184226
rect 97674 184046 97730 184102
rect 97798 184046 97854 184102
rect 97922 184046 97978 184102
rect 98046 184046 98102 184102
rect 97674 183922 97730 183978
rect 97798 183922 97854 183978
rect 97922 183922 97978 183978
rect 98046 183922 98102 183978
rect 70674 172294 70730 172350
rect 70798 172294 70854 172350
rect 70922 172294 70978 172350
rect 71046 172294 71102 172350
rect 70674 172170 70730 172226
rect 70798 172170 70854 172226
rect 70922 172170 70978 172226
rect 71046 172170 71102 172226
rect 70674 172046 70730 172102
rect 70798 172046 70854 172102
rect 70922 172046 70978 172102
rect 71046 172046 71102 172102
rect 70674 171922 70730 171978
rect 70798 171922 70854 171978
rect 70922 171922 70978 171978
rect 71046 171922 71102 171978
rect 70674 154294 70730 154350
rect 70798 154294 70854 154350
rect 70922 154294 70978 154350
rect 71046 154294 71102 154350
rect 70674 154170 70730 154226
rect 70798 154170 70854 154226
rect 70922 154170 70978 154226
rect 71046 154170 71102 154226
rect 70674 154046 70730 154102
rect 70798 154046 70854 154102
rect 70922 154046 70978 154102
rect 71046 154046 71102 154102
rect 70674 153922 70730 153978
rect 70798 153922 70854 153978
rect 70922 153922 70978 153978
rect 71046 153922 71102 153978
rect 66954 130294 67010 130350
rect 67078 130294 67134 130350
rect 67202 130294 67258 130350
rect 67326 130294 67382 130350
rect 66954 130170 67010 130226
rect 67078 130170 67134 130226
rect 67202 130170 67258 130226
rect 67326 130170 67382 130226
rect 66954 130046 67010 130102
rect 67078 130046 67134 130102
rect 67202 130046 67258 130102
rect 67326 130046 67382 130102
rect 66954 129922 67010 129978
rect 67078 129922 67134 129978
rect 67202 129922 67258 129978
rect 67326 129922 67382 129978
rect 64204 117422 64260 117478
rect 24518 112294 24574 112350
rect 24642 112294 24698 112350
rect 24518 112170 24574 112226
rect 24642 112170 24698 112226
rect 24518 112046 24574 112102
rect 24642 112046 24698 112102
rect 24518 111922 24574 111978
rect 24642 111922 24698 111978
rect 36234 112294 36290 112350
rect 36358 112294 36414 112350
rect 36482 112294 36538 112350
rect 36606 112294 36662 112350
rect 36234 112170 36290 112226
rect 36358 112170 36414 112226
rect 36482 112170 36538 112226
rect 36606 112170 36662 112226
rect 36234 112046 36290 112102
rect 36358 112046 36414 112102
rect 36482 112046 36538 112102
rect 36606 112046 36662 112102
rect 36234 111922 36290 111978
rect 36358 111922 36414 111978
rect 36482 111922 36538 111978
rect 36606 111922 36662 111978
rect 9234 100294 9290 100350
rect 9358 100294 9414 100350
rect 9482 100294 9538 100350
rect 9606 100294 9662 100350
rect 9234 100170 9290 100226
rect 9358 100170 9414 100226
rect 9482 100170 9538 100226
rect 9606 100170 9662 100226
rect 9234 100046 9290 100102
rect 9358 100046 9414 100102
rect 9482 100046 9538 100102
rect 9606 100046 9662 100102
rect 9234 99922 9290 99978
rect 9358 99922 9414 99978
rect 9482 99922 9538 99978
rect 9606 99922 9662 99978
rect 9234 82294 9290 82350
rect 9358 82294 9414 82350
rect 9482 82294 9538 82350
rect 9606 82294 9662 82350
rect 9234 82170 9290 82226
rect 9358 82170 9414 82226
rect 9482 82170 9538 82226
rect 9606 82170 9662 82226
rect 9234 82046 9290 82102
rect 9358 82046 9414 82102
rect 9482 82046 9538 82102
rect 9606 82046 9662 82102
rect 9234 81922 9290 81978
rect 9358 81922 9414 81978
rect 9482 81922 9538 81978
rect 9606 81922 9662 81978
rect 55238 112294 55294 112350
rect 55362 112294 55418 112350
rect 55238 112170 55294 112226
rect 55362 112170 55418 112226
rect 55238 112046 55294 112102
rect 55362 112046 55418 112102
rect 55238 111922 55294 111978
rect 55362 111922 55418 111978
rect 117238 184294 117294 184350
rect 117362 184294 117418 184350
rect 117238 184170 117294 184226
rect 117362 184170 117418 184226
rect 117238 184046 117294 184102
rect 117362 184046 117418 184102
rect 117238 183922 117294 183978
rect 117362 183922 117418 183978
rect 128394 184294 128450 184350
rect 128518 184294 128574 184350
rect 128642 184294 128698 184350
rect 128766 184294 128822 184350
rect 128394 184170 128450 184226
rect 128518 184170 128574 184226
rect 128642 184170 128698 184226
rect 128766 184170 128822 184226
rect 128394 184046 128450 184102
rect 128518 184046 128574 184102
rect 128642 184046 128698 184102
rect 128766 184046 128822 184102
rect 128394 183922 128450 183978
rect 128518 183922 128574 183978
rect 128642 183922 128698 183978
rect 128766 183922 128822 183978
rect 97674 166294 97730 166350
rect 97798 166294 97854 166350
rect 97922 166294 97978 166350
rect 98046 166294 98102 166350
rect 97674 166170 97730 166226
rect 97798 166170 97854 166226
rect 97922 166170 97978 166226
rect 98046 166170 98102 166226
rect 97674 166046 97730 166102
rect 97798 166046 97854 166102
rect 97922 166046 97978 166102
rect 98046 166046 98102 166102
rect 97674 165922 97730 165978
rect 97798 165922 97854 165978
rect 97922 165922 97978 165978
rect 98046 165922 98102 165978
rect 70674 136294 70730 136350
rect 70798 136294 70854 136350
rect 70922 136294 70978 136350
rect 71046 136294 71102 136350
rect 70674 136170 70730 136226
rect 70798 136170 70854 136226
rect 70922 136170 70978 136226
rect 71046 136170 71102 136226
rect 70674 136046 70730 136102
rect 70798 136046 70854 136102
rect 70922 136046 70978 136102
rect 71046 136046 71102 136102
rect 70674 135922 70730 135978
rect 70798 135922 70854 135978
rect 70922 135922 70978 135978
rect 71046 135922 71102 135978
rect 66954 112294 67010 112350
rect 67078 112294 67134 112350
rect 67202 112294 67258 112350
rect 67326 112294 67382 112350
rect 66954 112170 67010 112226
rect 67078 112170 67134 112226
rect 67202 112170 67258 112226
rect 67326 112170 67382 112226
rect 66954 112046 67010 112102
rect 67078 112046 67134 112102
rect 67202 112046 67258 112102
rect 67326 112046 67382 112102
rect 66954 111922 67010 111978
rect 67078 111922 67134 111978
rect 67202 111922 67258 111978
rect 67326 111922 67382 111978
rect 36234 94294 36290 94350
rect 36358 94294 36414 94350
rect 36482 94294 36538 94350
rect 36606 94294 36662 94350
rect 36234 94170 36290 94226
rect 36358 94170 36414 94226
rect 36482 94170 36538 94226
rect 36606 94170 36662 94226
rect 36234 94046 36290 94102
rect 36358 94046 36414 94102
rect 36482 94046 36538 94102
rect 36606 94046 36662 94102
rect 36234 93922 36290 93978
rect 36358 93922 36414 93978
rect 36482 93922 36538 93978
rect 36606 93922 36662 93978
rect 36234 76294 36290 76350
rect 36358 76294 36414 76350
rect 36482 76294 36538 76350
rect 36606 76294 36662 76350
rect 36234 76170 36290 76226
rect 36358 76170 36414 76226
rect 36482 76170 36538 76226
rect 36606 76170 36662 76226
rect 36234 76046 36290 76102
rect 36358 76046 36414 76102
rect 36482 76046 36538 76102
rect 36606 76046 36662 76102
rect 36234 75922 36290 75978
rect 36358 75922 36414 75978
rect 36482 75922 36538 75978
rect 36606 75922 36662 75978
rect 9234 64294 9290 64350
rect 9358 64294 9414 64350
rect 9482 64294 9538 64350
rect 9606 64294 9662 64350
rect 9234 64170 9290 64226
rect 9358 64170 9414 64226
rect 9482 64170 9538 64226
rect 9606 64170 9662 64226
rect 9234 64046 9290 64102
rect 9358 64046 9414 64102
rect 9482 64046 9538 64102
rect 9606 64046 9662 64102
rect 9234 63922 9290 63978
rect 9358 63922 9414 63978
rect 9482 63922 9538 63978
rect 9606 63922 9662 63978
rect 9234 46294 9290 46350
rect 9358 46294 9414 46350
rect 9482 46294 9538 46350
rect 9606 46294 9662 46350
rect 9234 46170 9290 46226
rect 9358 46170 9414 46226
rect 9482 46170 9538 46226
rect 9606 46170 9662 46226
rect 9234 46046 9290 46102
rect 9358 46046 9414 46102
rect 9482 46046 9538 46102
rect 9606 46046 9662 46102
rect 9234 45922 9290 45978
rect 9358 45922 9414 45978
rect 9482 45922 9538 45978
rect 9606 45922 9662 45978
rect 18396 55502 18452 55558
rect 9234 28294 9290 28350
rect 9358 28294 9414 28350
rect 9482 28294 9538 28350
rect 9606 28294 9662 28350
rect 9234 28170 9290 28226
rect 9358 28170 9414 28226
rect 9482 28170 9538 28226
rect 9606 28170 9662 28226
rect 9234 28046 9290 28102
rect 9358 28046 9414 28102
rect 9482 28046 9538 28102
rect 9606 28046 9662 28102
rect 9234 27922 9290 27978
rect 9358 27922 9414 27978
rect 9482 27922 9538 27978
rect 9606 27922 9662 27978
rect 9234 10294 9290 10350
rect 9358 10294 9414 10350
rect 9482 10294 9538 10350
rect 9606 10294 9662 10350
rect 9234 10170 9290 10226
rect 9358 10170 9414 10226
rect 9482 10170 9538 10226
rect 9606 10170 9662 10226
rect 9234 10046 9290 10102
rect 9358 10046 9414 10102
rect 9482 10046 9538 10102
rect 9606 10046 9662 10102
rect 9234 9922 9290 9978
rect 9358 9922 9414 9978
rect 9482 9922 9538 9978
rect 9606 9922 9662 9978
rect 24518 58294 24574 58350
rect 24642 58294 24698 58350
rect 24518 58170 24574 58226
rect 24642 58170 24698 58226
rect 24518 58046 24574 58102
rect 24642 58046 24698 58102
rect 24518 57922 24574 57978
rect 24642 57922 24698 57978
rect 39954 100294 40010 100350
rect 40078 100294 40134 100350
rect 40202 100294 40258 100350
rect 40326 100294 40382 100350
rect 39954 100170 40010 100226
rect 40078 100170 40134 100226
rect 40202 100170 40258 100226
rect 40326 100170 40382 100226
rect 39954 100046 40010 100102
rect 40078 100046 40134 100102
rect 40202 100046 40258 100102
rect 40326 100046 40382 100102
rect 39954 99922 40010 99978
rect 40078 99922 40134 99978
rect 40202 99922 40258 99978
rect 40326 99922 40382 99978
rect 39954 82294 40010 82350
rect 40078 82294 40134 82350
rect 40202 82294 40258 82350
rect 40326 82294 40382 82350
rect 39954 82170 40010 82226
rect 40078 82170 40134 82226
rect 40202 82170 40258 82226
rect 40326 82170 40382 82226
rect 39954 82046 40010 82102
rect 40078 82046 40134 82102
rect 40202 82046 40258 82102
rect 40326 82046 40382 82102
rect 39954 81922 40010 81978
rect 40078 81922 40134 81978
rect 40202 81922 40258 81978
rect 40326 81922 40382 81978
rect 73836 126062 73892 126118
rect 80444 132722 80500 132778
rect 97674 148294 97730 148350
rect 97798 148294 97854 148350
rect 97922 148294 97978 148350
rect 98046 148294 98102 148350
rect 97674 148170 97730 148226
rect 97798 148170 97854 148226
rect 97922 148170 97978 148226
rect 98046 148170 98102 148226
rect 97674 148046 97730 148102
rect 97798 148046 97854 148102
rect 97922 148046 97978 148102
rect 98046 148046 98102 148102
rect 97674 147922 97730 147978
rect 97798 147922 97854 147978
rect 97922 147922 97978 147978
rect 98046 147922 98102 147978
rect 86518 130294 86574 130350
rect 86642 130294 86698 130350
rect 86518 130170 86574 130226
rect 86642 130170 86698 130226
rect 86518 130046 86574 130102
rect 86642 130046 86698 130102
rect 86518 129922 86574 129978
rect 86642 129922 86698 129978
rect 101394 172294 101450 172350
rect 101518 172294 101574 172350
rect 101642 172294 101698 172350
rect 101766 172294 101822 172350
rect 101394 172170 101450 172226
rect 101518 172170 101574 172226
rect 101642 172170 101698 172226
rect 101766 172170 101822 172226
rect 101394 172046 101450 172102
rect 101518 172046 101574 172102
rect 101642 172046 101698 172102
rect 101766 172046 101822 172102
rect 101394 171922 101450 171978
rect 101518 171922 101574 171978
rect 101642 171922 101698 171978
rect 101766 171922 101822 171978
rect 128394 166294 128450 166350
rect 128518 166294 128574 166350
rect 128642 166294 128698 166350
rect 128766 166294 128822 166350
rect 128394 166170 128450 166226
rect 128518 166170 128574 166226
rect 128642 166170 128698 166226
rect 128766 166170 128822 166226
rect 128394 166046 128450 166102
rect 128518 166046 128574 166102
rect 128642 166046 128698 166102
rect 128766 166046 128822 166102
rect 128394 165922 128450 165978
rect 128518 165922 128574 165978
rect 128642 165922 128698 165978
rect 128766 165922 128822 165978
rect 101394 154294 101450 154350
rect 101518 154294 101574 154350
rect 101642 154294 101698 154350
rect 101766 154294 101822 154350
rect 101394 154170 101450 154226
rect 101518 154170 101574 154226
rect 101642 154170 101698 154226
rect 101766 154170 101822 154226
rect 101394 154046 101450 154102
rect 101518 154046 101574 154102
rect 101642 154046 101698 154102
rect 101766 154046 101822 154102
rect 101394 153922 101450 153978
rect 101518 153922 101574 153978
rect 101642 153922 101698 153978
rect 101766 153922 101822 153978
rect 101878 136294 101934 136350
rect 102002 136294 102058 136350
rect 101878 136170 101934 136226
rect 102002 136170 102058 136226
rect 101878 136046 101934 136102
rect 102002 136046 102058 136102
rect 101878 135922 101934 135978
rect 102002 135922 102058 135978
rect 97674 130294 97730 130350
rect 97798 130294 97854 130350
rect 97922 130294 97978 130350
rect 98046 130294 98102 130350
rect 97674 130170 97730 130226
rect 97798 130170 97854 130226
rect 97922 130170 97978 130226
rect 98046 130170 98102 130226
rect 97674 130046 97730 130102
rect 97798 130046 97854 130102
rect 97922 130046 97978 130102
rect 98046 130046 98102 130102
rect 97674 129922 97730 129978
rect 97798 129922 97854 129978
rect 97922 129922 97978 129978
rect 98046 129922 98102 129978
rect 82684 127682 82740 127738
rect 82460 125882 82516 125938
rect 70674 118294 70730 118350
rect 70798 118294 70854 118350
rect 70922 118294 70978 118350
rect 71046 118294 71102 118350
rect 70674 118170 70730 118226
rect 70798 118170 70854 118226
rect 70922 118170 70978 118226
rect 71046 118170 71102 118226
rect 70674 118046 70730 118102
rect 70798 118046 70854 118102
rect 70922 118046 70978 118102
rect 71046 118046 71102 118102
rect 70674 117922 70730 117978
rect 70798 117922 70854 117978
rect 70922 117922 70978 117978
rect 71046 117922 71102 117978
rect 86518 112294 86574 112350
rect 86642 112294 86698 112350
rect 86518 112170 86574 112226
rect 86642 112170 86698 112226
rect 86518 112046 86574 112102
rect 86642 112046 86698 112102
rect 86518 111922 86574 111978
rect 86642 111922 86698 111978
rect 117238 130294 117294 130350
rect 117362 130294 117418 130350
rect 117238 130170 117294 130226
rect 117362 130170 117418 130226
rect 117238 130046 117294 130102
rect 117362 130046 117418 130102
rect 117238 129922 117294 129978
rect 117362 129922 117418 129978
rect 128394 148294 128450 148350
rect 128518 148294 128574 148350
rect 128642 148294 128698 148350
rect 128766 148294 128822 148350
rect 128394 148170 128450 148226
rect 128518 148170 128574 148226
rect 128642 148170 128698 148226
rect 128766 148170 128822 148226
rect 128394 148046 128450 148102
rect 128518 148046 128574 148102
rect 128642 148046 128698 148102
rect 128766 148046 128822 148102
rect 128394 147922 128450 147978
rect 128518 147922 128574 147978
rect 128642 147922 128698 147978
rect 128766 147922 128822 147978
rect 128394 130294 128450 130350
rect 128518 130294 128574 130350
rect 128642 130294 128698 130350
rect 128766 130294 128822 130350
rect 128394 130170 128450 130226
rect 128518 130170 128574 130226
rect 128642 130170 128698 130226
rect 128766 130170 128822 130226
rect 128394 130046 128450 130102
rect 128518 130046 128574 130102
rect 128642 130046 128698 130102
rect 128766 130046 128822 130102
rect 128394 129922 128450 129978
rect 128518 129922 128574 129978
rect 128642 129922 128698 129978
rect 128766 129922 128822 129978
rect 101878 118294 101934 118350
rect 102002 118294 102058 118350
rect 101878 118170 101934 118226
rect 102002 118170 102058 118226
rect 101878 118046 101934 118102
rect 102002 118046 102058 118102
rect 101878 117922 101934 117978
rect 102002 117922 102058 117978
rect 97674 112294 97730 112350
rect 97798 112294 97854 112350
rect 97922 112294 97978 112350
rect 98046 112294 98102 112350
rect 97674 112170 97730 112226
rect 97798 112170 97854 112226
rect 97922 112170 97978 112226
rect 98046 112170 98102 112226
rect 97674 112046 97730 112102
rect 97798 112046 97854 112102
rect 97922 112046 97978 112102
rect 98046 112046 98102 112102
rect 97674 111922 97730 111978
rect 97798 111922 97854 111978
rect 97922 111922 97978 111978
rect 98046 111922 98102 111978
rect 70674 100294 70730 100350
rect 70798 100294 70854 100350
rect 70922 100294 70978 100350
rect 71046 100294 71102 100350
rect 70674 100170 70730 100226
rect 70798 100170 70854 100226
rect 70922 100170 70978 100226
rect 71046 100170 71102 100226
rect 70674 100046 70730 100102
rect 70798 100046 70854 100102
rect 70922 100046 70978 100102
rect 71046 100046 71102 100102
rect 70674 99922 70730 99978
rect 70798 99922 70854 99978
rect 70922 99922 70978 99978
rect 71046 99922 71102 99978
rect 66954 94294 67010 94350
rect 67078 94294 67134 94350
rect 67202 94294 67258 94350
rect 67326 94294 67382 94350
rect 66954 94170 67010 94226
rect 67078 94170 67134 94226
rect 67202 94170 67258 94226
rect 67326 94170 67382 94226
rect 66954 94046 67010 94102
rect 67078 94046 67134 94102
rect 67202 94046 67258 94102
rect 67326 94046 67382 94102
rect 66954 93922 67010 93978
rect 67078 93922 67134 93978
rect 67202 93922 67258 93978
rect 67326 93922 67382 93978
rect 66954 76294 67010 76350
rect 67078 76294 67134 76350
rect 67202 76294 67258 76350
rect 67326 76294 67382 76350
rect 66954 76170 67010 76226
rect 67078 76170 67134 76226
rect 67202 76170 67258 76226
rect 67326 76170 67382 76226
rect 66954 76046 67010 76102
rect 67078 76046 67134 76102
rect 67202 76046 67258 76102
rect 67326 76046 67382 76102
rect 66954 75922 67010 75978
rect 67078 75922 67134 75978
rect 67202 75922 67258 75978
rect 67326 75922 67382 75978
rect 39878 64294 39934 64350
rect 40002 64294 40058 64350
rect 39878 64170 39934 64226
rect 40002 64170 40058 64226
rect 39878 64046 39934 64102
rect 40002 64046 40058 64102
rect 39878 63922 39934 63978
rect 40002 63922 40058 63978
rect 36234 58294 36290 58350
rect 36358 58294 36414 58350
rect 36482 58294 36538 58350
rect 36606 58294 36662 58350
rect 36234 58170 36290 58226
rect 36358 58170 36414 58226
rect 36482 58170 36538 58226
rect 36606 58170 36662 58226
rect 36234 58046 36290 58102
rect 36358 58046 36414 58102
rect 36482 58046 36538 58102
rect 36606 58046 36662 58102
rect 36234 57922 36290 57978
rect 36358 57922 36414 57978
rect 36482 57922 36538 57978
rect 36606 57922 36662 57978
rect 24518 40294 24574 40350
rect 24642 40294 24698 40350
rect 24518 40170 24574 40226
rect 24642 40170 24698 40226
rect 24518 40046 24574 40102
rect 24642 40046 24698 40102
rect 24518 39922 24574 39978
rect 24642 39922 24698 39978
rect 55238 58294 55294 58350
rect 55362 58294 55418 58350
rect 55238 58170 55294 58226
rect 55362 58170 55418 58226
rect 55238 58046 55294 58102
rect 55362 58046 55418 58102
rect 55238 57922 55294 57978
rect 55362 57922 55418 57978
rect 66954 58294 67010 58350
rect 67078 58294 67134 58350
rect 67202 58294 67258 58350
rect 67326 58294 67382 58350
rect 66954 58170 67010 58226
rect 67078 58170 67134 58226
rect 67202 58170 67258 58226
rect 67326 58170 67382 58226
rect 66954 58046 67010 58102
rect 67078 58046 67134 58102
rect 67202 58046 67258 58102
rect 67326 58046 67382 58102
rect 66954 57922 67010 57978
rect 67078 57922 67134 57978
rect 67202 57922 67258 57978
rect 67326 57922 67382 57978
rect 39878 46294 39934 46350
rect 40002 46294 40058 46350
rect 39878 46170 39934 46226
rect 40002 46170 40058 46226
rect 39878 46046 39934 46102
rect 40002 46046 40058 46102
rect 39878 45922 39934 45978
rect 40002 45922 40058 45978
rect 36234 40294 36290 40350
rect 36358 40294 36414 40350
rect 36482 40294 36538 40350
rect 36606 40294 36662 40350
rect 36234 40170 36290 40226
rect 36358 40170 36414 40226
rect 36482 40170 36538 40226
rect 36606 40170 36662 40226
rect 36234 40046 36290 40102
rect 36358 40046 36414 40102
rect 36482 40046 36538 40102
rect 36606 40046 36662 40102
rect 36234 39922 36290 39978
rect 36358 39922 36414 39978
rect 36482 39922 36538 39978
rect 36606 39922 36662 39978
rect 55238 40294 55294 40350
rect 55362 40294 55418 40350
rect 55238 40170 55294 40226
rect 55362 40170 55418 40226
rect 55238 40046 55294 40102
rect 55362 40046 55418 40102
rect 55238 39922 55294 39978
rect 55362 39922 55418 39978
rect 70674 82294 70730 82350
rect 70798 82294 70854 82350
rect 70922 82294 70978 82350
rect 71046 82294 71102 82350
rect 70674 82170 70730 82226
rect 70798 82170 70854 82226
rect 70922 82170 70978 82226
rect 71046 82170 71102 82226
rect 70674 82046 70730 82102
rect 70798 82046 70854 82102
rect 70922 82046 70978 82102
rect 71046 82046 71102 82102
rect 70674 81922 70730 81978
rect 70798 81922 70854 81978
rect 70922 81922 70978 81978
rect 71046 81922 71102 81978
rect 70674 64294 70730 64350
rect 70798 64294 70854 64350
rect 70922 64294 70978 64350
rect 71046 64294 71102 64350
rect 70674 64170 70730 64226
rect 70798 64170 70854 64226
rect 70922 64170 70978 64226
rect 71046 64170 71102 64226
rect 70674 64046 70730 64102
rect 70798 64046 70854 64102
rect 70922 64046 70978 64102
rect 71046 64046 71102 64102
rect 70674 63922 70730 63978
rect 70798 63922 70854 63978
rect 70922 63922 70978 63978
rect 71046 63922 71102 63978
rect 70674 46294 70730 46350
rect 70798 46294 70854 46350
rect 70922 46294 70978 46350
rect 71046 46294 71102 46350
rect 70674 46170 70730 46226
rect 70798 46170 70854 46226
rect 70922 46170 70978 46226
rect 71046 46170 71102 46226
rect 70674 46046 70730 46102
rect 70798 46046 70854 46102
rect 70922 46046 70978 46102
rect 71046 46046 71102 46102
rect 117238 112294 117294 112350
rect 117362 112294 117418 112350
rect 117238 112170 117294 112226
rect 117362 112170 117418 112226
rect 117238 112046 117294 112102
rect 117362 112046 117418 112102
rect 117238 111922 117294 111978
rect 117362 111922 117418 111978
rect 128394 112294 128450 112350
rect 128518 112294 128574 112350
rect 128642 112294 128698 112350
rect 128766 112294 128822 112350
rect 128394 112170 128450 112226
rect 128518 112170 128574 112226
rect 128642 112170 128698 112226
rect 128766 112170 128822 112226
rect 128394 112046 128450 112102
rect 128518 112046 128574 112102
rect 128642 112046 128698 112102
rect 128766 112046 128822 112102
rect 128394 111922 128450 111978
rect 128518 111922 128574 111978
rect 128642 111922 128698 111978
rect 128766 111922 128822 111978
rect 97674 94294 97730 94350
rect 97798 94294 97854 94350
rect 97922 94294 97978 94350
rect 98046 94294 98102 94350
rect 97674 94170 97730 94226
rect 97798 94170 97854 94226
rect 97922 94170 97978 94226
rect 98046 94170 98102 94226
rect 97674 94046 97730 94102
rect 97798 94046 97854 94102
rect 97922 94046 97978 94102
rect 98046 94046 98102 94102
rect 97674 93922 97730 93978
rect 97798 93922 97854 93978
rect 97922 93922 97978 93978
rect 98046 93922 98102 93978
rect 97674 76294 97730 76350
rect 97798 76294 97854 76350
rect 97922 76294 97978 76350
rect 98046 76294 98102 76350
rect 97674 76170 97730 76226
rect 97798 76170 97854 76226
rect 97922 76170 97978 76226
rect 98046 76170 98102 76226
rect 97674 76046 97730 76102
rect 97798 76046 97854 76102
rect 97922 76046 97978 76102
rect 98046 76046 98102 76102
rect 97674 75922 97730 75978
rect 97798 75922 97854 75978
rect 97922 75922 97978 75978
rect 98046 75922 98102 75978
rect 86518 58294 86574 58350
rect 86642 58294 86698 58350
rect 86518 58170 86574 58226
rect 86642 58170 86698 58226
rect 86518 58046 86574 58102
rect 86642 58046 86698 58102
rect 86518 57922 86574 57978
rect 86642 57922 86698 57978
rect 101394 100294 101450 100350
rect 101518 100294 101574 100350
rect 101642 100294 101698 100350
rect 101766 100294 101822 100350
rect 101394 100170 101450 100226
rect 101518 100170 101574 100226
rect 101642 100170 101698 100226
rect 101766 100170 101822 100226
rect 101394 100046 101450 100102
rect 101518 100046 101574 100102
rect 101642 100046 101698 100102
rect 101766 100046 101822 100102
rect 101394 99922 101450 99978
rect 101518 99922 101574 99978
rect 101642 99922 101698 99978
rect 101766 99922 101822 99978
rect 128394 94294 128450 94350
rect 128518 94294 128574 94350
rect 128642 94294 128698 94350
rect 128766 94294 128822 94350
rect 128394 94170 128450 94226
rect 128518 94170 128574 94226
rect 128642 94170 128698 94226
rect 128766 94170 128822 94226
rect 128394 94046 128450 94102
rect 128518 94046 128574 94102
rect 128642 94046 128698 94102
rect 128766 94046 128822 94102
rect 128394 93922 128450 93978
rect 128518 93922 128574 93978
rect 128642 93922 128698 93978
rect 128766 93922 128822 93978
rect 101394 82294 101450 82350
rect 101518 82294 101574 82350
rect 101642 82294 101698 82350
rect 101766 82294 101822 82350
rect 101394 82170 101450 82226
rect 101518 82170 101574 82226
rect 101642 82170 101698 82226
rect 101766 82170 101822 82226
rect 101394 82046 101450 82102
rect 101518 82046 101574 82102
rect 101642 82046 101698 82102
rect 101766 82046 101822 82102
rect 101394 81922 101450 81978
rect 101518 81922 101574 81978
rect 101642 81922 101698 81978
rect 101766 81922 101822 81978
rect 101878 64294 101934 64350
rect 102002 64294 102058 64350
rect 101878 64170 101934 64226
rect 102002 64170 102058 64226
rect 101878 64046 101934 64102
rect 102002 64046 102058 64102
rect 101878 63922 101934 63978
rect 102002 63922 102058 63978
rect 97674 58294 97730 58350
rect 97798 58294 97854 58350
rect 97922 58294 97978 58350
rect 98046 58294 98102 58350
rect 97674 58170 97730 58226
rect 97798 58170 97854 58226
rect 97922 58170 97978 58226
rect 98046 58170 98102 58226
rect 97674 58046 97730 58102
rect 97798 58046 97854 58102
rect 97922 58046 97978 58102
rect 98046 58046 98102 58102
rect 97674 57922 97730 57978
rect 97798 57922 97854 57978
rect 97922 57922 97978 57978
rect 98046 57922 98102 57978
rect 82684 56222 82740 56278
rect 117238 58294 117294 58350
rect 117362 58294 117418 58350
rect 117238 58170 117294 58226
rect 117362 58170 117418 58226
rect 117238 58046 117294 58102
rect 117362 58046 117418 58102
rect 117238 57922 117294 57978
rect 117362 57922 117418 57978
rect 132114 208294 132170 208350
rect 132238 208294 132294 208350
rect 132362 208294 132418 208350
rect 132486 208294 132542 208350
rect 132114 208170 132170 208226
rect 132238 208170 132294 208226
rect 132362 208170 132418 208226
rect 132486 208170 132542 208226
rect 132114 208046 132170 208102
rect 132238 208046 132294 208102
rect 132362 208046 132418 208102
rect 132486 208046 132542 208102
rect 132114 207922 132170 207978
rect 132238 207922 132294 207978
rect 132362 207922 132418 207978
rect 132486 207922 132542 207978
rect 132114 190294 132170 190350
rect 132238 190294 132294 190350
rect 132362 190294 132418 190350
rect 132486 190294 132542 190350
rect 132114 190170 132170 190226
rect 132238 190170 132294 190226
rect 132362 190170 132418 190226
rect 132486 190170 132542 190226
rect 132114 190046 132170 190102
rect 132238 190046 132294 190102
rect 132362 190046 132418 190102
rect 132486 190046 132542 190102
rect 132114 189922 132170 189978
rect 132238 189922 132294 189978
rect 132362 189922 132418 189978
rect 132486 189922 132542 189978
rect 134428 192122 134484 192178
rect 159114 220294 159170 220350
rect 159238 220294 159294 220350
rect 159362 220294 159418 220350
rect 159486 220294 159542 220350
rect 159114 220170 159170 220226
rect 159238 220170 159294 220226
rect 159362 220170 159418 220226
rect 159486 220170 159542 220226
rect 159114 220046 159170 220102
rect 159238 220046 159294 220102
rect 159362 220046 159418 220102
rect 159486 220046 159542 220102
rect 159114 219922 159170 219978
rect 159238 219922 159294 219978
rect 159362 219922 159418 219978
rect 159486 219922 159542 219978
rect 148518 202294 148574 202350
rect 148642 202294 148698 202350
rect 148518 202170 148574 202226
rect 148642 202170 148698 202226
rect 148518 202046 148574 202102
rect 148642 202046 148698 202102
rect 148518 201922 148574 201978
rect 148642 201922 148698 201978
rect 162834 261996 162890 262052
rect 162958 261996 163014 262052
rect 163082 261996 163138 262052
rect 163206 261996 163262 262052
rect 162834 261872 162890 261928
rect 162958 261872 163014 261928
rect 163082 261872 163138 261928
rect 163206 261872 163262 261928
rect 163878 262046 163934 262102
rect 164002 262046 164058 262102
rect 163878 261922 163934 261978
rect 164002 261922 164058 261978
rect 189834 274294 189890 274350
rect 189958 274294 190014 274350
rect 190082 274294 190138 274350
rect 190206 274294 190262 274350
rect 189834 274170 189890 274226
rect 189958 274170 190014 274226
rect 190082 274170 190138 274226
rect 190206 274170 190262 274226
rect 189834 274046 189890 274102
rect 189958 274046 190014 274102
rect 190082 274046 190138 274102
rect 190206 274046 190262 274102
rect 189834 273922 189890 273978
rect 189958 273922 190014 273978
rect 190082 273922 190138 273978
rect 190206 273922 190262 273978
rect 189532 264842 189588 264898
rect 179238 256294 179294 256350
rect 179362 256294 179418 256350
rect 179238 256170 179294 256226
rect 179362 256170 179418 256226
rect 179238 256046 179294 256102
rect 179362 256046 179418 256102
rect 179238 255922 179294 255978
rect 179362 255922 179418 255978
rect 189834 256294 189890 256350
rect 189958 256294 190014 256350
rect 190082 256294 190138 256350
rect 190206 256294 190262 256350
rect 189834 256170 189890 256226
rect 189958 256170 190014 256226
rect 190082 256170 190138 256226
rect 190206 256170 190262 256226
rect 189834 256046 189890 256102
rect 189958 256046 190014 256102
rect 190082 256046 190138 256102
rect 190206 256046 190262 256102
rect 189834 255922 189890 255978
rect 189958 255922 190014 255978
rect 190082 255922 190138 255978
rect 190206 255922 190262 255978
rect 162834 244294 162890 244350
rect 162958 244294 163014 244350
rect 163082 244294 163138 244350
rect 163206 244294 163262 244350
rect 162834 244170 162890 244226
rect 162958 244170 163014 244226
rect 163082 244170 163138 244226
rect 163206 244170 163262 244226
rect 162834 244046 162890 244102
rect 162958 244046 163014 244102
rect 163082 244046 163138 244102
rect 163206 244046 163262 244102
rect 162834 243922 162890 243978
rect 162958 243922 163014 243978
rect 163082 243922 163138 243978
rect 163206 243922 163262 243978
rect 189834 238294 189890 238350
rect 189958 238294 190014 238350
rect 190082 238294 190138 238350
rect 190206 238294 190262 238350
rect 189834 238170 189890 238226
rect 189958 238170 190014 238226
rect 190082 238170 190138 238226
rect 190206 238170 190262 238226
rect 189834 238046 189890 238102
rect 189958 238046 190014 238102
rect 190082 238046 190138 238102
rect 190206 238046 190262 238102
rect 189834 237922 189890 237978
rect 189958 237922 190014 237978
rect 190082 237922 190138 237978
rect 190206 237922 190262 237978
rect 162834 226294 162890 226350
rect 162958 226294 163014 226350
rect 163082 226294 163138 226350
rect 163206 226294 163262 226350
rect 162834 226170 162890 226226
rect 162958 226170 163014 226226
rect 163082 226170 163138 226226
rect 163206 226170 163262 226226
rect 162834 226046 162890 226102
rect 162958 226046 163014 226102
rect 163082 226046 163138 226102
rect 163206 226046 163262 226102
rect 162834 225922 162890 225978
rect 162958 225922 163014 225978
rect 163082 225922 163138 225978
rect 163206 225922 163262 225978
rect 159114 202294 159170 202350
rect 159238 202294 159294 202350
rect 159362 202294 159418 202350
rect 159486 202294 159542 202350
rect 159114 202170 159170 202226
rect 159238 202170 159294 202226
rect 159362 202170 159418 202226
rect 159486 202170 159542 202226
rect 159114 202046 159170 202102
rect 159238 202046 159294 202102
rect 159362 202046 159418 202102
rect 159486 202046 159542 202102
rect 159114 201922 159170 201978
rect 159238 201922 159294 201978
rect 159362 201922 159418 201978
rect 159486 201922 159542 201978
rect 141036 198962 141092 199018
rect 148518 184294 148574 184350
rect 148642 184294 148698 184350
rect 148518 184170 148574 184226
rect 148642 184170 148698 184226
rect 148518 184046 148574 184102
rect 148642 184046 148698 184102
rect 148518 183922 148574 183978
rect 148642 183922 148698 183978
rect 162834 208294 162890 208350
rect 162958 208294 163014 208350
rect 163082 208294 163138 208350
rect 163206 208294 163262 208350
rect 162834 208170 162890 208226
rect 162958 208170 163014 208226
rect 163082 208170 163138 208226
rect 163206 208170 163262 208226
rect 162834 208046 162890 208102
rect 162958 208046 163014 208102
rect 163082 208046 163138 208102
rect 163206 208046 163262 208102
rect 162834 207922 162890 207978
rect 162958 207922 163014 207978
rect 163082 207922 163138 207978
rect 163206 207922 163262 207978
rect 163878 208294 163934 208350
rect 164002 208294 164058 208350
rect 163878 208170 163934 208226
rect 164002 208170 164058 208226
rect 163878 208046 163934 208102
rect 164002 208046 164058 208102
rect 163878 207922 163934 207978
rect 164002 207922 164058 207978
rect 179238 202294 179294 202350
rect 179362 202294 179418 202350
rect 179238 202170 179294 202226
rect 179362 202170 179418 202226
rect 179238 202046 179294 202102
rect 179362 202046 179418 202102
rect 179238 201922 179294 201978
rect 179362 201922 179418 201978
rect 187292 196622 187348 196678
rect 169708 193922 169764 193978
rect 163878 190294 163934 190350
rect 164002 190294 164058 190350
rect 163878 190170 163934 190226
rect 164002 190170 164058 190226
rect 163878 190046 163934 190102
rect 164002 190046 164058 190102
rect 163878 189922 163934 189978
rect 164002 189922 164058 189978
rect 169708 189602 169764 189658
rect 188076 195182 188132 195238
rect 193554 316294 193610 316350
rect 193678 316294 193734 316350
rect 193802 316294 193858 316350
rect 193926 316294 193982 316350
rect 193554 316170 193610 316226
rect 193678 316170 193734 316226
rect 193802 316170 193858 316226
rect 193926 316170 193982 316226
rect 193554 316046 193610 316102
rect 193678 316046 193734 316102
rect 193802 316046 193858 316102
rect 193926 316046 193982 316102
rect 193554 315922 193610 315978
rect 193678 315922 193734 315978
rect 193802 315922 193858 315978
rect 193926 315922 193982 315978
rect 193554 298294 193610 298350
rect 193678 298294 193734 298350
rect 193802 298294 193858 298350
rect 193926 298294 193982 298350
rect 193554 298170 193610 298226
rect 193678 298170 193734 298226
rect 193802 298170 193858 298226
rect 193926 298170 193982 298226
rect 193554 298046 193610 298102
rect 193678 298046 193734 298102
rect 193802 298046 193858 298102
rect 193926 298046 193982 298102
rect 193554 297922 193610 297978
rect 193678 297922 193734 297978
rect 193802 297922 193858 297978
rect 193926 297922 193982 297978
rect 193554 280294 193610 280350
rect 193678 280294 193734 280350
rect 193802 280294 193858 280350
rect 193926 280294 193982 280350
rect 193554 280170 193610 280226
rect 193678 280170 193734 280226
rect 193802 280170 193858 280226
rect 193926 280170 193982 280226
rect 193554 280046 193610 280102
rect 193678 280046 193734 280102
rect 193802 280046 193858 280102
rect 193926 280046 193982 280102
rect 193554 279922 193610 279978
rect 193678 279922 193734 279978
rect 193802 279922 193858 279978
rect 193926 279922 193982 279978
rect 195692 278162 195748 278218
rect 194908 271502 194964 271558
rect 194908 270062 194964 270118
rect 195692 267002 195748 267058
rect 198268 268802 198324 268858
rect 198268 264482 198324 264538
rect 193554 262294 193610 262350
rect 193678 262294 193734 262350
rect 193802 262294 193858 262350
rect 193926 262294 193982 262350
rect 193554 262170 193610 262226
rect 193678 262170 193734 262226
rect 193802 262170 193858 262226
rect 193926 262170 193982 262226
rect 193554 262046 193610 262102
rect 193678 262046 193734 262102
rect 193802 262046 193858 262102
rect 193926 262046 193982 262102
rect 193554 261922 193610 261978
rect 193678 261922 193734 261978
rect 193802 261922 193858 261978
rect 193926 261922 193982 261978
rect 199836 260162 199892 260218
rect 194908 258362 194964 258418
rect 193554 244294 193610 244350
rect 193678 244294 193734 244350
rect 193802 244294 193858 244350
rect 193926 244294 193982 244350
rect 193554 244170 193610 244226
rect 193678 244170 193734 244226
rect 193802 244170 193858 244226
rect 193926 244170 193982 244226
rect 193554 244046 193610 244102
rect 193678 244046 193734 244102
rect 193802 244046 193858 244102
rect 193926 244046 193982 244102
rect 193554 243922 193610 243978
rect 193678 243922 193734 243978
rect 193802 243922 193858 243978
rect 193926 243922 193982 243978
rect 193554 226294 193610 226350
rect 193678 226294 193734 226350
rect 193802 226294 193858 226350
rect 193926 226294 193982 226350
rect 193554 226170 193610 226226
rect 193678 226170 193734 226226
rect 193802 226170 193858 226226
rect 193926 226170 193982 226226
rect 193554 226046 193610 226102
rect 193678 226046 193734 226102
rect 193802 226046 193858 226102
rect 193926 226046 193982 226102
rect 193554 225922 193610 225978
rect 193678 225922 193734 225978
rect 193802 225922 193858 225978
rect 193926 225922 193982 225978
rect 189834 220294 189890 220350
rect 189958 220294 190014 220350
rect 190082 220294 190138 220350
rect 190206 220294 190262 220350
rect 189834 220170 189890 220226
rect 189958 220170 190014 220226
rect 190082 220170 190138 220226
rect 190206 220170 190262 220226
rect 189834 220046 189890 220102
rect 189958 220046 190014 220102
rect 190082 220046 190138 220102
rect 190206 220046 190262 220102
rect 189834 219922 189890 219978
rect 189958 219922 190014 219978
rect 190082 219922 190138 219978
rect 190206 219922 190262 219978
rect 189834 202294 189890 202350
rect 189958 202294 190014 202350
rect 190082 202294 190138 202350
rect 190206 202294 190262 202350
rect 189834 202170 189890 202226
rect 189958 202170 190014 202226
rect 190082 202170 190138 202226
rect 190206 202170 190262 202226
rect 189834 202046 189890 202102
rect 189958 202046 190014 202102
rect 190082 202046 190138 202102
rect 190206 202046 190262 202102
rect 189834 201922 189890 201978
rect 189958 201922 190014 201978
rect 190082 201922 190138 201978
rect 190206 201922 190262 201978
rect 189532 196442 189588 196498
rect 188076 189422 188132 189478
rect 187292 187442 187348 187498
rect 169708 187262 169764 187318
rect 169708 186002 169764 186058
rect 159114 184294 159170 184350
rect 159238 184294 159294 184350
rect 159362 184294 159418 184350
rect 159486 184294 159542 184350
rect 159114 184170 159170 184226
rect 159238 184170 159294 184226
rect 159362 184170 159418 184226
rect 159486 184170 159542 184226
rect 159114 184046 159170 184102
rect 159238 184046 159294 184102
rect 159362 184046 159418 184102
rect 159486 184046 159542 184102
rect 159114 183922 159170 183978
rect 159238 183922 159294 183978
rect 159362 183922 159418 183978
rect 159486 183922 159542 183978
rect 132114 172294 132170 172350
rect 132238 172294 132294 172350
rect 132362 172294 132418 172350
rect 132486 172294 132542 172350
rect 132114 172170 132170 172226
rect 132238 172170 132294 172226
rect 132362 172170 132418 172226
rect 132486 172170 132542 172226
rect 132114 172046 132170 172102
rect 132238 172046 132294 172102
rect 132362 172046 132418 172102
rect 132486 172046 132542 172102
rect 132114 171922 132170 171978
rect 132238 171922 132294 171978
rect 132362 171922 132418 171978
rect 132486 171922 132542 171978
rect 132114 154294 132170 154350
rect 132238 154294 132294 154350
rect 132362 154294 132418 154350
rect 132486 154294 132542 154350
rect 132114 154170 132170 154226
rect 132238 154170 132294 154226
rect 132362 154170 132418 154226
rect 132486 154170 132542 154226
rect 132114 154046 132170 154102
rect 132238 154046 132294 154102
rect 132362 154046 132418 154102
rect 132486 154046 132542 154102
rect 132114 153922 132170 153978
rect 132238 153922 132294 153978
rect 132362 153922 132418 153978
rect 132486 153922 132542 153978
rect 132114 136294 132170 136350
rect 132238 136294 132294 136350
rect 132362 136294 132418 136350
rect 132486 136294 132542 136350
rect 132114 136170 132170 136226
rect 132238 136170 132294 136226
rect 132362 136170 132418 136226
rect 132486 136170 132542 136226
rect 132114 136046 132170 136102
rect 132238 136046 132294 136102
rect 132362 136046 132418 136102
rect 132486 136046 132542 136102
rect 132114 135922 132170 135978
rect 132238 135922 132294 135978
rect 132362 135922 132418 135978
rect 132486 135922 132542 135978
rect 138572 132902 138628 132958
rect 138572 125882 138628 125938
rect 159114 166294 159170 166350
rect 159238 166294 159294 166350
rect 159362 166294 159418 166350
rect 159486 166294 159542 166350
rect 159114 166170 159170 166226
rect 159238 166170 159294 166226
rect 159362 166170 159418 166226
rect 159486 166170 159542 166226
rect 159114 166046 159170 166102
rect 159238 166046 159294 166102
rect 159362 166046 159418 166102
rect 159486 166046 159542 166102
rect 159114 165922 159170 165978
rect 159238 165922 159294 165978
rect 159362 165922 159418 165978
rect 159486 165922 159542 165978
rect 159114 148294 159170 148350
rect 159238 148294 159294 148350
rect 159362 148294 159418 148350
rect 159486 148294 159542 148350
rect 159114 148170 159170 148226
rect 159238 148170 159294 148226
rect 159362 148170 159418 148226
rect 159486 148170 159542 148226
rect 159114 148046 159170 148102
rect 159238 148046 159294 148102
rect 159362 148046 159418 148102
rect 159486 148046 159542 148102
rect 159114 147922 159170 147978
rect 159238 147922 159294 147978
rect 159362 147922 159418 147978
rect 159486 147922 159542 147978
rect 141932 137762 141988 137818
rect 141036 127682 141092 127738
rect 132114 118294 132170 118350
rect 132238 118294 132294 118350
rect 132362 118294 132418 118350
rect 132486 118294 132542 118350
rect 132114 118170 132170 118226
rect 132238 118170 132294 118226
rect 132362 118170 132418 118226
rect 132486 118170 132542 118226
rect 132114 118046 132170 118102
rect 132238 118046 132294 118102
rect 132362 118046 132418 118102
rect 132486 118046 132542 118102
rect 132114 117922 132170 117978
rect 132238 117922 132294 117978
rect 132362 117922 132418 117978
rect 132486 117922 132542 117978
rect 148518 130294 148574 130350
rect 148642 130294 148698 130350
rect 148518 130170 148574 130226
rect 148642 130170 148698 130226
rect 148518 130046 148574 130102
rect 148642 130046 148698 130102
rect 148518 129922 148574 129978
rect 148642 129922 148698 129978
rect 159114 130294 159170 130350
rect 159238 130294 159294 130350
rect 159362 130294 159418 130350
rect 159486 130294 159542 130350
rect 159114 130170 159170 130226
rect 159238 130170 159294 130226
rect 159362 130170 159418 130226
rect 159486 130170 159542 130226
rect 159114 130046 159170 130102
rect 159238 130046 159294 130102
rect 159362 130046 159418 130102
rect 159486 130046 159542 130102
rect 159114 129922 159170 129978
rect 159238 129922 159294 129978
rect 159362 129922 159418 129978
rect 159486 129922 159542 129978
rect 144060 128042 144116 128098
rect 148518 112294 148574 112350
rect 148642 112294 148698 112350
rect 148518 112170 148574 112226
rect 148642 112170 148698 112226
rect 148518 112046 148574 112102
rect 148642 112046 148698 112102
rect 148518 111922 148574 111978
rect 148642 111922 148698 111978
rect 179238 184294 179294 184350
rect 179362 184294 179418 184350
rect 179238 184170 179294 184226
rect 179362 184170 179418 184226
rect 179238 184046 179294 184102
rect 179362 184046 179418 184102
rect 179238 183922 179294 183978
rect 179362 183922 179418 183978
rect 191548 195002 191604 195058
rect 193554 208294 193610 208350
rect 193678 208294 193734 208350
rect 193802 208294 193858 208350
rect 193926 208294 193982 208350
rect 193554 208170 193610 208226
rect 193678 208170 193734 208226
rect 193802 208170 193858 208226
rect 193926 208170 193982 208226
rect 193554 208046 193610 208102
rect 193678 208046 193734 208102
rect 193802 208046 193858 208102
rect 193926 208046 193982 208102
rect 193554 207922 193610 207978
rect 193678 207922 193734 207978
rect 193802 207922 193858 207978
rect 193926 207922 193982 207978
rect 191548 186002 191604 186058
rect 196588 196802 196644 196858
rect 197484 196622 197540 196678
rect 193554 190294 193610 190350
rect 193678 190294 193734 190350
rect 193802 190294 193858 190350
rect 193926 190294 193982 190350
rect 193554 190170 193610 190226
rect 193678 190170 193734 190226
rect 193802 190170 193858 190226
rect 193926 190170 193982 190226
rect 193554 190046 193610 190102
rect 193678 190046 193734 190102
rect 193802 190046 193858 190102
rect 193926 190046 193982 190102
rect 193554 189922 193610 189978
rect 193678 189922 193734 189978
rect 193802 189922 193858 189978
rect 193926 189922 193982 189978
rect 189834 184294 189890 184350
rect 189958 184294 190014 184350
rect 190082 184294 190138 184350
rect 190206 184294 190262 184350
rect 189834 184170 189890 184226
rect 189958 184170 190014 184226
rect 190082 184170 190138 184226
rect 190206 184170 190262 184226
rect 189834 184046 189890 184102
rect 189958 184046 190014 184102
rect 190082 184046 190138 184102
rect 190206 184046 190262 184102
rect 189834 183922 189890 183978
rect 189958 183922 190014 183978
rect 190082 183922 190138 183978
rect 190206 183922 190262 183978
rect 162834 172294 162890 172350
rect 162958 172294 163014 172350
rect 163082 172294 163138 172350
rect 163206 172294 163262 172350
rect 162834 172170 162890 172226
rect 162958 172170 163014 172226
rect 163082 172170 163138 172226
rect 163206 172170 163262 172226
rect 162834 172046 162890 172102
rect 162958 172046 163014 172102
rect 163082 172046 163138 172102
rect 163206 172046 163262 172102
rect 162834 171922 162890 171978
rect 162958 171922 163014 171978
rect 163082 171922 163138 171978
rect 163206 171922 163262 171978
rect 162834 154294 162890 154350
rect 162958 154294 163014 154350
rect 163082 154294 163138 154350
rect 163206 154294 163262 154350
rect 162834 154170 162890 154226
rect 162958 154170 163014 154226
rect 163082 154170 163138 154226
rect 163206 154170 163262 154226
rect 162834 154046 162890 154102
rect 162958 154046 163014 154102
rect 163082 154046 163138 154102
rect 163206 154046 163262 154102
rect 162834 153922 162890 153978
rect 162958 153922 163014 153978
rect 163082 153922 163138 153978
rect 163206 153922 163262 153978
rect 162834 136294 162890 136350
rect 162958 136294 163014 136350
rect 163082 136294 163138 136350
rect 163206 136294 163262 136350
rect 162834 136170 162890 136226
rect 162958 136170 163014 136226
rect 163082 136170 163138 136226
rect 163206 136170 163262 136226
rect 162834 136046 162890 136102
rect 162958 136046 163014 136102
rect 163082 136046 163138 136102
rect 163206 136046 163262 136102
rect 162834 135922 162890 135978
rect 162958 135922 163014 135978
rect 163082 135922 163138 135978
rect 163206 135922 163262 135978
rect 163878 136294 163934 136350
rect 164002 136294 164058 136350
rect 163878 136170 163934 136226
rect 164002 136170 164058 136226
rect 163878 136046 163934 136102
rect 164002 136046 164058 136102
rect 163878 135922 163934 135978
rect 164002 135922 164058 135978
rect 179238 130294 179294 130350
rect 179362 130294 179418 130350
rect 179238 130170 179294 130226
rect 179362 130170 179418 130226
rect 179238 130046 179294 130102
rect 179362 130046 179418 130102
rect 179238 129922 179294 129978
rect 179362 129922 179418 129978
rect 189834 166294 189890 166350
rect 189958 166294 190014 166350
rect 190082 166294 190138 166350
rect 190206 166294 190262 166350
rect 189834 166170 189890 166226
rect 189958 166170 190014 166226
rect 190082 166170 190138 166226
rect 190206 166170 190262 166226
rect 189834 166046 189890 166102
rect 189958 166046 190014 166102
rect 190082 166046 190138 166102
rect 190206 166046 190262 166102
rect 189834 165922 189890 165978
rect 189958 165922 190014 165978
rect 190082 165922 190138 165978
rect 190206 165922 190262 165978
rect 193554 172294 193610 172350
rect 193678 172294 193734 172350
rect 193802 172294 193858 172350
rect 193926 172294 193982 172350
rect 193554 172170 193610 172226
rect 193678 172170 193734 172226
rect 193802 172170 193858 172226
rect 193926 172170 193982 172226
rect 193554 172046 193610 172102
rect 193678 172046 193734 172102
rect 193802 172046 193858 172102
rect 193926 172046 193982 172102
rect 193554 171922 193610 171978
rect 193678 171922 193734 171978
rect 193802 171922 193858 171978
rect 193926 171922 193982 171978
rect 189834 148294 189890 148350
rect 189958 148294 190014 148350
rect 190082 148294 190138 148350
rect 190206 148294 190262 148350
rect 189834 148170 189890 148226
rect 189958 148170 190014 148226
rect 190082 148170 190138 148226
rect 190206 148170 190262 148226
rect 189834 148046 189890 148102
rect 189958 148046 190014 148102
rect 190082 148046 190138 148102
rect 190206 148046 190262 148102
rect 189834 147922 189890 147978
rect 189958 147922 190014 147978
rect 190082 147922 190138 147978
rect 190206 147922 190262 147978
rect 189834 130294 189890 130350
rect 189958 130294 190014 130350
rect 190082 130294 190138 130350
rect 190206 130294 190262 130350
rect 189834 130170 189890 130226
rect 189958 130170 190014 130226
rect 190082 130170 190138 130226
rect 190206 130170 190262 130226
rect 189834 130046 189890 130102
rect 189958 130046 190014 130102
rect 190082 130046 190138 130102
rect 190206 130046 190262 130102
rect 189834 129922 189890 129978
rect 189958 129922 190014 129978
rect 190082 129922 190138 129978
rect 190206 129922 190262 129978
rect 159114 112294 159170 112350
rect 159238 112294 159294 112350
rect 159362 112294 159418 112350
rect 159486 112294 159542 112350
rect 159114 112170 159170 112226
rect 159238 112170 159294 112226
rect 159362 112170 159418 112226
rect 159486 112170 159542 112226
rect 159114 112046 159170 112102
rect 159238 112046 159294 112102
rect 159362 112046 159418 112102
rect 159486 112046 159542 112102
rect 159114 111922 159170 111978
rect 159238 111922 159294 111978
rect 159362 111922 159418 111978
rect 159486 111922 159542 111978
rect 132114 100294 132170 100350
rect 132238 100294 132294 100350
rect 132362 100294 132418 100350
rect 132486 100294 132542 100350
rect 132114 100170 132170 100226
rect 132238 100170 132294 100226
rect 132362 100170 132418 100226
rect 132486 100170 132542 100226
rect 132114 100046 132170 100102
rect 132238 100046 132294 100102
rect 132362 100046 132418 100102
rect 132486 100046 132542 100102
rect 132114 99922 132170 99978
rect 132238 99922 132294 99978
rect 132362 99922 132418 99978
rect 132486 99922 132542 99978
rect 132114 82294 132170 82350
rect 132238 82294 132294 82350
rect 132362 82294 132418 82350
rect 132486 82294 132542 82350
rect 132114 82170 132170 82226
rect 132238 82170 132294 82226
rect 132362 82170 132418 82226
rect 132486 82170 132542 82226
rect 132114 82046 132170 82102
rect 132238 82046 132294 82102
rect 132362 82046 132418 82102
rect 132486 82046 132542 82102
rect 132114 81922 132170 81978
rect 132238 81922 132294 81978
rect 132362 81922 132418 81978
rect 132486 81922 132542 81978
rect 128394 76294 128450 76350
rect 128518 76294 128574 76350
rect 128642 76294 128698 76350
rect 128766 76294 128822 76350
rect 128394 76170 128450 76226
rect 128518 76170 128574 76226
rect 128642 76170 128698 76226
rect 128766 76170 128822 76226
rect 128394 76046 128450 76102
rect 128518 76046 128574 76102
rect 128642 76046 128698 76102
rect 128766 76046 128822 76102
rect 128394 75922 128450 75978
rect 128518 75922 128574 75978
rect 128642 75922 128698 75978
rect 128766 75922 128822 75978
rect 128394 58294 128450 58350
rect 128518 58294 128574 58350
rect 128642 58294 128698 58350
rect 128766 58294 128822 58350
rect 128394 58170 128450 58226
rect 128518 58170 128574 58226
rect 128642 58170 128698 58226
rect 128766 58170 128822 58226
rect 128394 58046 128450 58102
rect 128518 58046 128574 58102
rect 128642 58046 128698 58102
rect 128766 58046 128822 58102
rect 128394 57922 128450 57978
rect 128518 57922 128574 57978
rect 128642 57922 128698 57978
rect 128766 57922 128822 57978
rect 101878 46294 101934 46350
rect 102002 46294 102058 46350
rect 101878 46170 101934 46226
rect 102002 46170 102058 46226
rect 70674 45922 70730 45978
rect 70798 45922 70854 45978
rect 70922 45922 70978 45978
rect 71046 45922 71102 45978
rect 66954 40294 67010 40350
rect 67078 40294 67134 40350
rect 67202 40294 67258 40350
rect 67326 40294 67382 40350
rect 66954 40170 67010 40226
rect 67078 40170 67134 40226
rect 67202 40170 67258 40226
rect 67326 40170 67382 40226
rect 66954 40046 67010 40102
rect 67078 40046 67134 40102
rect 67202 40046 67258 40102
rect 67326 40046 67382 40102
rect 66954 39922 67010 39978
rect 67078 39922 67134 39978
rect 67202 39922 67258 39978
rect 67326 39922 67382 39978
rect 36234 22294 36290 22350
rect 36358 22294 36414 22350
rect 36482 22294 36538 22350
rect 36606 22294 36662 22350
rect 36234 22170 36290 22226
rect 36358 22170 36414 22226
rect 36482 22170 36538 22226
rect 36606 22170 36662 22226
rect 36234 22046 36290 22102
rect 36358 22046 36414 22102
rect 36482 22046 36538 22102
rect 36606 22046 36662 22102
rect 36234 21922 36290 21978
rect 36358 21922 36414 21978
rect 36482 21922 36538 21978
rect 36606 21922 36662 21978
rect 9234 -1176 9290 -1120
rect 9358 -1176 9414 -1120
rect 9482 -1176 9538 -1120
rect 9606 -1176 9662 -1120
rect 9234 -1300 9290 -1244
rect 9358 -1300 9414 -1244
rect 9482 -1300 9538 -1244
rect 9606 -1300 9662 -1244
rect 9234 -1424 9290 -1368
rect 9358 -1424 9414 -1368
rect 9482 -1424 9538 -1368
rect 9606 -1424 9662 -1368
rect 9234 -1548 9290 -1492
rect 9358 -1548 9414 -1492
rect 9482 -1548 9538 -1492
rect 9606 -1548 9662 -1492
rect 36234 4294 36290 4350
rect 36358 4294 36414 4350
rect 36482 4294 36538 4350
rect 36606 4294 36662 4350
rect 36234 4170 36290 4226
rect 36358 4170 36414 4226
rect 36482 4170 36538 4226
rect 36606 4170 36662 4226
rect 36234 4046 36290 4102
rect 36358 4046 36414 4102
rect 36482 4046 36538 4102
rect 36606 4046 36662 4102
rect 36234 3922 36290 3978
rect 36358 3922 36414 3978
rect 36482 3922 36538 3978
rect 36606 3922 36662 3978
rect 36234 -216 36290 -160
rect 36358 -216 36414 -160
rect 36482 -216 36538 -160
rect 36606 -216 36662 -160
rect 36234 -340 36290 -284
rect 36358 -340 36414 -284
rect 36482 -340 36538 -284
rect 36606 -340 36662 -284
rect 36234 -464 36290 -408
rect 36358 -464 36414 -408
rect 36482 -464 36538 -408
rect 36606 -464 36662 -408
rect 36234 -588 36290 -532
rect 36358 -588 36414 -532
rect 36482 -588 36538 -532
rect 36606 -588 36662 -532
rect 39954 28294 40010 28350
rect 40078 28294 40134 28350
rect 40202 28294 40258 28350
rect 40326 28294 40382 28350
rect 39954 28170 40010 28226
rect 40078 28170 40134 28226
rect 40202 28170 40258 28226
rect 40326 28170 40382 28226
rect 39954 28046 40010 28102
rect 40078 28046 40134 28102
rect 40202 28046 40258 28102
rect 40326 28046 40382 28102
rect 39954 27922 40010 27978
rect 40078 27922 40134 27978
rect 40202 27922 40258 27978
rect 40326 27922 40382 27978
rect 39954 10294 40010 10350
rect 40078 10294 40134 10350
rect 40202 10294 40258 10350
rect 40326 10294 40382 10350
rect 39954 10170 40010 10226
rect 40078 10170 40134 10226
rect 40202 10170 40258 10226
rect 40326 10170 40382 10226
rect 39954 10046 40010 10102
rect 40078 10046 40134 10102
rect 40202 10046 40258 10102
rect 40326 10046 40382 10102
rect 39954 9922 40010 9978
rect 40078 9922 40134 9978
rect 40202 9922 40258 9978
rect 40326 9922 40382 9978
rect 39954 -1176 40010 -1120
rect 40078 -1176 40134 -1120
rect 40202 -1176 40258 -1120
rect 40326 -1176 40382 -1120
rect 39954 -1300 40010 -1244
rect 40078 -1300 40134 -1244
rect 40202 -1300 40258 -1244
rect 40326 -1300 40382 -1244
rect 39954 -1424 40010 -1368
rect 40078 -1424 40134 -1368
rect 40202 -1424 40258 -1368
rect 40326 -1424 40382 -1368
rect 39954 -1548 40010 -1492
rect 40078 -1548 40134 -1492
rect 40202 -1548 40258 -1492
rect 40326 -1548 40382 -1492
rect 66954 22294 67010 22350
rect 67078 22294 67134 22350
rect 67202 22294 67258 22350
rect 67326 22294 67382 22350
rect 66954 22170 67010 22226
rect 67078 22170 67134 22226
rect 67202 22170 67258 22226
rect 67326 22170 67382 22226
rect 66954 22046 67010 22102
rect 67078 22046 67134 22102
rect 67202 22046 67258 22102
rect 67326 22046 67382 22102
rect 66954 21922 67010 21978
rect 67078 21922 67134 21978
rect 67202 21922 67258 21978
rect 67326 21922 67382 21978
rect 66954 4294 67010 4350
rect 67078 4294 67134 4350
rect 67202 4294 67258 4350
rect 67326 4294 67382 4350
rect 66954 4170 67010 4226
rect 67078 4170 67134 4226
rect 67202 4170 67258 4226
rect 67326 4170 67382 4226
rect 66954 4046 67010 4102
rect 67078 4046 67134 4102
rect 67202 4046 67258 4102
rect 67326 4046 67382 4102
rect 66954 3922 67010 3978
rect 67078 3922 67134 3978
rect 67202 3922 67258 3978
rect 67326 3922 67382 3978
rect 66954 -216 67010 -160
rect 67078 -216 67134 -160
rect 67202 -216 67258 -160
rect 67326 -216 67382 -160
rect 66954 -340 67010 -284
rect 67078 -340 67134 -284
rect 67202 -340 67258 -284
rect 67326 -340 67382 -284
rect 66954 -464 67010 -408
rect 67078 -464 67134 -408
rect 67202 -464 67258 -408
rect 67326 -464 67382 -408
rect 66954 -588 67010 -532
rect 67078 -588 67134 -532
rect 67202 -588 67258 -532
rect 67326 -588 67382 -532
rect 101878 46046 101934 46102
rect 102002 46046 102058 46102
rect 101878 45922 101934 45978
rect 102002 45922 102058 45978
rect 86518 40294 86574 40350
rect 86642 40294 86698 40350
rect 86518 40170 86574 40226
rect 86642 40170 86698 40226
rect 86518 40046 86574 40102
rect 86642 40046 86698 40102
rect 86518 39922 86574 39978
rect 86642 39922 86698 39978
rect 97674 40294 97730 40350
rect 97798 40294 97854 40350
rect 97922 40294 97978 40350
rect 98046 40294 98102 40350
rect 97674 40170 97730 40226
rect 97798 40170 97854 40226
rect 97922 40170 97978 40226
rect 98046 40170 98102 40226
rect 97674 40046 97730 40102
rect 97798 40046 97854 40102
rect 97922 40046 97978 40102
rect 98046 40046 98102 40102
rect 97674 39922 97730 39978
rect 97798 39922 97854 39978
rect 97922 39922 97978 39978
rect 98046 39922 98102 39978
rect 70674 28294 70730 28350
rect 70798 28294 70854 28350
rect 70922 28294 70978 28350
rect 71046 28294 71102 28350
rect 70674 28170 70730 28226
rect 70798 28170 70854 28226
rect 70922 28170 70978 28226
rect 71046 28170 71102 28226
rect 70674 28046 70730 28102
rect 70798 28046 70854 28102
rect 70922 28046 70978 28102
rect 71046 28046 71102 28102
rect 70674 27922 70730 27978
rect 70798 27922 70854 27978
rect 70922 27922 70978 27978
rect 71046 27922 71102 27978
rect 70674 10294 70730 10350
rect 70798 10294 70854 10350
rect 70922 10294 70978 10350
rect 71046 10294 71102 10350
rect 70674 10170 70730 10226
rect 70798 10170 70854 10226
rect 70922 10170 70978 10226
rect 71046 10170 71102 10226
rect 70674 10046 70730 10102
rect 70798 10046 70854 10102
rect 70922 10046 70978 10102
rect 71046 10046 71102 10102
rect 70674 9922 70730 9978
rect 70798 9922 70854 9978
rect 70922 9922 70978 9978
rect 71046 9922 71102 9978
rect 70674 -1176 70730 -1120
rect 70798 -1176 70854 -1120
rect 70922 -1176 70978 -1120
rect 71046 -1176 71102 -1120
rect 70674 -1300 70730 -1244
rect 70798 -1300 70854 -1244
rect 70922 -1300 70978 -1244
rect 71046 -1300 71102 -1244
rect 70674 -1424 70730 -1368
rect 70798 -1424 70854 -1368
rect 70922 -1424 70978 -1368
rect 71046 -1424 71102 -1368
rect 70674 -1548 70730 -1492
rect 70798 -1548 70854 -1492
rect 70922 -1548 70978 -1492
rect 71046 -1548 71102 -1492
rect 117238 40294 117294 40350
rect 117362 40294 117418 40350
rect 117238 40170 117294 40226
rect 117362 40170 117418 40226
rect 117238 40046 117294 40102
rect 117362 40046 117418 40102
rect 117238 39922 117294 39978
rect 117362 39922 117418 39978
rect 132114 64294 132170 64350
rect 132238 64294 132294 64350
rect 132362 64294 132418 64350
rect 132486 64294 132542 64350
rect 132114 64170 132170 64226
rect 132238 64170 132294 64226
rect 132362 64170 132418 64226
rect 132486 64170 132542 64226
rect 132114 64046 132170 64102
rect 132238 64046 132294 64102
rect 132362 64046 132418 64102
rect 132486 64046 132542 64102
rect 132114 63922 132170 63978
rect 132238 63922 132294 63978
rect 132362 63922 132418 63978
rect 132486 63922 132542 63978
rect 128394 40294 128450 40350
rect 128518 40294 128574 40350
rect 128642 40294 128698 40350
rect 128766 40294 128822 40350
rect 128394 40170 128450 40226
rect 128518 40170 128574 40226
rect 128642 40170 128698 40226
rect 128766 40170 128822 40226
rect 128394 40046 128450 40102
rect 128518 40046 128574 40102
rect 128642 40046 128698 40102
rect 128766 40046 128822 40102
rect 128394 39922 128450 39978
rect 128518 39922 128574 39978
rect 128642 39922 128698 39978
rect 128766 39922 128822 39978
rect 97674 22294 97730 22350
rect 97798 22294 97854 22350
rect 97922 22294 97978 22350
rect 98046 22294 98102 22350
rect 97674 22170 97730 22226
rect 97798 22170 97854 22226
rect 97922 22170 97978 22226
rect 98046 22170 98102 22226
rect 97674 22046 97730 22102
rect 97798 22046 97854 22102
rect 97922 22046 97978 22102
rect 98046 22046 98102 22102
rect 97674 21922 97730 21978
rect 97798 21922 97854 21978
rect 97922 21922 97978 21978
rect 98046 21922 98102 21978
rect 97674 4294 97730 4350
rect 97798 4294 97854 4350
rect 97922 4294 97978 4350
rect 98046 4294 98102 4350
rect 97674 4170 97730 4226
rect 97798 4170 97854 4226
rect 97922 4170 97978 4226
rect 98046 4170 98102 4226
rect 97674 4046 97730 4102
rect 97798 4046 97854 4102
rect 97922 4046 97978 4102
rect 98046 4046 98102 4102
rect 97674 3922 97730 3978
rect 97798 3922 97854 3978
rect 97922 3922 97978 3978
rect 98046 3922 98102 3978
rect 97674 -216 97730 -160
rect 97798 -216 97854 -160
rect 97922 -216 97978 -160
rect 98046 -216 98102 -160
rect 97674 -340 97730 -284
rect 97798 -340 97854 -284
rect 97922 -340 97978 -284
rect 98046 -340 98102 -284
rect 97674 -464 97730 -408
rect 97798 -464 97854 -408
rect 97922 -464 97978 -408
rect 98046 -464 98102 -408
rect 97674 -588 97730 -532
rect 97798 -588 97854 -532
rect 97922 -588 97978 -532
rect 98046 -588 98102 -532
rect 101394 28294 101450 28350
rect 101518 28294 101574 28350
rect 101642 28294 101698 28350
rect 101766 28294 101822 28350
rect 101394 28170 101450 28226
rect 101518 28170 101574 28226
rect 101642 28170 101698 28226
rect 101766 28170 101822 28226
rect 101394 28046 101450 28102
rect 101518 28046 101574 28102
rect 101642 28046 101698 28102
rect 101766 28046 101822 28102
rect 101394 27922 101450 27978
rect 101518 27922 101574 27978
rect 101642 27922 101698 27978
rect 101766 27922 101822 27978
rect 101394 10294 101450 10350
rect 101518 10294 101574 10350
rect 101642 10294 101698 10350
rect 101766 10294 101822 10350
rect 101394 10170 101450 10226
rect 101518 10170 101574 10226
rect 101642 10170 101698 10226
rect 101766 10170 101822 10226
rect 101394 10046 101450 10102
rect 101518 10046 101574 10102
rect 101642 10046 101698 10102
rect 101766 10046 101822 10102
rect 101394 9922 101450 9978
rect 101518 9922 101574 9978
rect 101642 9922 101698 9978
rect 101766 9922 101822 9978
rect 101394 -1176 101450 -1120
rect 101518 -1176 101574 -1120
rect 101642 -1176 101698 -1120
rect 101766 -1176 101822 -1120
rect 101394 -1300 101450 -1244
rect 101518 -1300 101574 -1244
rect 101642 -1300 101698 -1244
rect 101766 -1300 101822 -1244
rect 101394 -1424 101450 -1368
rect 101518 -1424 101574 -1368
rect 101642 -1424 101698 -1368
rect 101766 -1424 101822 -1368
rect 101394 -1548 101450 -1492
rect 101518 -1548 101574 -1492
rect 101642 -1548 101698 -1492
rect 101766 -1548 101822 -1492
rect 128394 22294 128450 22350
rect 128518 22294 128574 22350
rect 128642 22294 128698 22350
rect 128766 22294 128822 22350
rect 128394 22170 128450 22226
rect 128518 22170 128574 22226
rect 128642 22170 128698 22226
rect 128766 22170 128822 22226
rect 128394 22046 128450 22102
rect 128518 22046 128574 22102
rect 128642 22046 128698 22102
rect 128766 22046 128822 22102
rect 128394 21922 128450 21978
rect 128518 21922 128574 21978
rect 128642 21922 128698 21978
rect 128766 21922 128822 21978
rect 128394 4294 128450 4350
rect 128518 4294 128574 4350
rect 128642 4294 128698 4350
rect 128766 4294 128822 4350
rect 128394 4170 128450 4226
rect 128518 4170 128574 4226
rect 128642 4170 128698 4226
rect 128766 4170 128822 4226
rect 128394 4046 128450 4102
rect 128518 4046 128574 4102
rect 128642 4046 128698 4102
rect 128766 4046 128822 4102
rect 128394 3922 128450 3978
rect 128518 3922 128574 3978
rect 128642 3922 128698 3978
rect 128766 3922 128822 3978
rect 128394 -216 128450 -160
rect 128518 -216 128574 -160
rect 128642 -216 128698 -160
rect 128766 -216 128822 -160
rect 128394 -340 128450 -284
rect 128518 -340 128574 -284
rect 128642 -340 128698 -284
rect 128766 -340 128822 -284
rect 128394 -464 128450 -408
rect 128518 -464 128574 -408
rect 128642 -464 128698 -408
rect 128766 -464 128822 -408
rect 128394 -588 128450 -532
rect 128518 -588 128574 -532
rect 128642 -588 128698 -532
rect 128766 -588 128822 -532
rect 132114 46294 132170 46350
rect 132238 46294 132294 46350
rect 132362 46294 132418 46350
rect 132486 46294 132542 46350
rect 132114 46170 132170 46226
rect 132238 46170 132294 46226
rect 132362 46170 132418 46226
rect 132486 46170 132542 46226
rect 132114 46046 132170 46102
rect 132238 46046 132294 46102
rect 132362 46046 132418 46102
rect 132486 46046 132542 46102
rect 132114 45922 132170 45978
rect 132238 45922 132294 45978
rect 132362 45922 132418 45978
rect 132486 45922 132542 45978
rect 141036 56222 141092 56278
rect 162834 118294 162890 118350
rect 162958 118294 163014 118350
rect 163082 118294 163138 118350
rect 163206 118294 163262 118350
rect 162834 118170 162890 118226
rect 162958 118170 163014 118226
rect 163082 118170 163138 118226
rect 163206 118170 163262 118226
rect 162834 118046 162890 118102
rect 162958 118046 163014 118102
rect 163082 118046 163138 118102
rect 163206 118046 163262 118102
rect 162834 117922 162890 117978
rect 162958 117922 163014 117978
rect 163082 117922 163138 117978
rect 163206 117922 163262 117978
rect 159114 94294 159170 94350
rect 159238 94294 159294 94350
rect 159362 94294 159418 94350
rect 159486 94294 159542 94350
rect 159114 94170 159170 94226
rect 159238 94170 159294 94226
rect 159362 94170 159418 94226
rect 159486 94170 159542 94226
rect 159114 94046 159170 94102
rect 159238 94046 159294 94102
rect 159362 94046 159418 94102
rect 159486 94046 159542 94102
rect 159114 93922 159170 93978
rect 159238 93922 159294 93978
rect 159362 93922 159418 93978
rect 159486 93922 159542 93978
rect 144060 56222 144116 56278
rect 159114 76294 159170 76350
rect 159238 76294 159294 76350
rect 159362 76294 159418 76350
rect 159486 76294 159542 76350
rect 159114 76170 159170 76226
rect 159238 76170 159294 76226
rect 159362 76170 159418 76226
rect 159486 76170 159542 76226
rect 159114 76046 159170 76102
rect 159238 76046 159294 76102
rect 159362 76046 159418 76102
rect 159486 76046 159542 76102
rect 159114 75922 159170 75978
rect 159238 75922 159294 75978
rect 159362 75922 159418 75978
rect 159486 75922 159542 75978
rect 148518 58294 148574 58350
rect 148642 58294 148698 58350
rect 148518 58170 148574 58226
rect 148642 58170 148698 58226
rect 148518 58046 148574 58102
rect 148642 58046 148698 58102
rect 148518 57922 148574 57978
rect 148642 57922 148698 57978
rect 159114 58294 159170 58350
rect 159238 58294 159294 58350
rect 159362 58294 159418 58350
rect 159486 58294 159542 58350
rect 159114 58170 159170 58226
rect 159238 58170 159294 58226
rect 159362 58170 159418 58226
rect 159486 58170 159542 58226
rect 159114 58046 159170 58102
rect 159238 58046 159294 58102
rect 159362 58046 159418 58102
rect 159486 58046 159542 58102
rect 159114 57922 159170 57978
rect 159238 57922 159294 57978
rect 159362 57922 159418 57978
rect 159486 57922 159542 57978
rect 148518 40294 148574 40350
rect 148642 40294 148698 40350
rect 148518 40170 148574 40226
rect 148642 40170 148698 40226
rect 148518 40046 148574 40102
rect 148642 40046 148698 40102
rect 148518 39922 148574 39978
rect 148642 39922 148698 39978
rect 163878 118294 163934 118350
rect 164002 118294 164058 118350
rect 163878 118170 163934 118226
rect 164002 118170 164058 118226
rect 163878 118046 163934 118102
rect 164002 118046 164058 118102
rect 163878 117922 163934 117978
rect 164002 117922 164058 117978
rect 179238 112294 179294 112350
rect 179362 112294 179418 112350
rect 179238 112170 179294 112226
rect 179362 112170 179418 112226
rect 179238 112046 179294 112102
rect 179362 112046 179418 112102
rect 179238 111922 179294 111978
rect 179362 111922 179418 111978
rect 193554 154294 193610 154350
rect 193678 154294 193734 154350
rect 193802 154294 193858 154350
rect 193926 154294 193982 154350
rect 193554 154170 193610 154226
rect 193678 154170 193734 154226
rect 193802 154170 193858 154226
rect 193926 154170 193982 154226
rect 193554 154046 193610 154102
rect 193678 154046 193734 154102
rect 193802 154046 193858 154102
rect 193926 154046 193982 154102
rect 193554 153922 193610 153978
rect 193678 153922 193734 153978
rect 193802 153922 193858 153978
rect 193926 153922 193982 153978
rect 193554 136294 193610 136350
rect 193678 136294 193734 136350
rect 193802 136294 193858 136350
rect 193926 136294 193982 136350
rect 193554 136170 193610 136226
rect 193678 136170 193734 136226
rect 193802 136170 193858 136226
rect 193926 136170 193982 136226
rect 193554 136046 193610 136102
rect 193678 136046 193734 136102
rect 193802 136046 193858 136102
rect 193926 136046 193982 136102
rect 193554 135922 193610 135978
rect 193678 135922 193734 135978
rect 193802 135922 193858 135978
rect 193926 135922 193982 135978
rect 189834 112294 189890 112350
rect 189958 112294 190014 112350
rect 190082 112294 190138 112350
rect 190206 112294 190262 112350
rect 189834 112170 189890 112226
rect 189958 112170 190014 112226
rect 190082 112170 190138 112226
rect 190206 112170 190262 112226
rect 189834 112046 189890 112102
rect 189958 112046 190014 112102
rect 190082 112046 190138 112102
rect 190206 112046 190262 112102
rect 189834 111922 189890 111978
rect 189958 111922 190014 111978
rect 190082 111922 190138 111978
rect 190206 111922 190262 111978
rect 162834 100294 162890 100350
rect 162958 100294 163014 100350
rect 163082 100294 163138 100350
rect 163206 100294 163262 100350
rect 162834 100170 162890 100226
rect 162958 100170 163014 100226
rect 163082 100170 163138 100226
rect 163206 100170 163262 100226
rect 162834 100046 162890 100102
rect 162958 100046 163014 100102
rect 163082 100046 163138 100102
rect 163206 100046 163262 100102
rect 162834 99922 162890 99978
rect 162958 99922 163014 99978
rect 163082 99922 163138 99978
rect 163206 99922 163262 99978
rect 189834 94294 189890 94350
rect 189958 94294 190014 94350
rect 190082 94294 190138 94350
rect 190206 94294 190262 94350
rect 189834 94170 189890 94226
rect 189958 94170 190014 94226
rect 190082 94170 190138 94226
rect 190206 94170 190262 94226
rect 189834 94046 189890 94102
rect 189958 94046 190014 94102
rect 190082 94046 190138 94102
rect 190206 94046 190262 94102
rect 189834 93922 189890 93978
rect 189958 93922 190014 93978
rect 190082 93922 190138 93978
rect 190206 93922 190262 93978
rect 162834 82294 162890 82350
rect 162958 82294 163014 82350
rect 163082 82294 163138 82350
rect 163206 82294 163262 82350
rect 162834 82170 162890 82226
rect 162958 82170 163014 82226
rect 163082 82170 163138 82226
rect 163206 82170 163262 82226
rect 162834 82046 162890 82102
rect 162958 82046 163014 82102
rect 163082 82046 163138 82102
rect 163206 82046 163262 82102
rect 162834 81922 162890 81978
rect 162958 81922 163014 81978
rect 163082 81922 163138 81978
rect 163206 81922 163262 81978
rect 162834 64294 162890 64350
rect 162958 64294 163014 64350
rect 163082 64294 163138 64350
rect 163206 64294 163262 64350
rect 162834 64170 162890 64226
rect 162958 64170 163014 64226
rect 163082 64170 163138 64226
rect 163206 64170 163262 64226
rect 162834 64046 162890 64102
rect 162958 64046 163014 64102
rect 163082 64046 163138 64102
rect 163206 64046 163262 64102
rect 162834 63922 162890 63978
rect 162958 63922 163014 63978
rect 163082 63922 163138 63978
rect 163206 63922 163262 63978
rect 163878 64294 163934 64350
rect 164002 64294 164058 64350
rect 163878 64170 163934 64226
rect 164002 64170 164058 64226
rect 163878 64046 163934 64102
rect 164002 64046 164058 64102
rect 163878 63922 163934 63978
rect 164002 63922 164058 63978
rect 179238 58294 179294 58350
rect 179362 58294 179418 58350
rect 179238 58170 179294 58226
rect 179362 58170 179418 58226
rect 179238 58046 179294 58102
rect 179362 58046 179418 58102
rect 179238 57922 179294 57978
rect 179362 57922 179418 57978
rect 189834 76294 189890 76350
rect 189958 76294 190014 76350
rect 190082 76294 190138 76350
rect 190206 76294 190262 76350
rect 189834 76170 189890 76226
rect 189958 76170 190014 76226
rect 190082 76170 190138 76226
rect 190206 76170 190262 76226
rect 189834 76046 189890 76102
rect 189958 76046 190014 76102
rect 190082 76046 190138 76102
rect 190206 76046 190262 76102
rect 189834 75922 189890 75978
rect 189958 75922 190014 75978
rect 190082 75922 190138 75978
rect 190206 75922 190262 75978
rect 189834 58294 189890 58350
rect 189958 58294 190014 58350
rect 190082 58294 190138 58350
rect 190206 58294 190262 58350
rect 189834 58170 189890 58226
rect 189958 58170 190014 58226
rect 190082 58170 190138 58226
rect 190206 58170 190262 58226
rect 189834 58046 189890 58102
rect 189958 58046 190014 58102
rect 190082 58046 190138 58102
rect 190206 58046 190262 58102
rect 189834 57922 189890 57978
rect 189958 57922 190014 57978
rect 190082 57922 190138 57978
rect 190206 57922 190262 57978
rect 159114 40294 159170 40350
rect 159238 40294 159294 40350
rect 159362 40294 159418 40350
rect 159486 40294 159542 40350
rect 159114 40170 159170 40226
rect 159238 40170 159294 40226
rect 159362 40170 159418 40226
rect 159486 40170 159542 40226
rect 159114 40046 159170 40102
rect 159238 40046 159294 40102
rect 159362 40046 159418 40102
rect 159486 40046 159542 40102
rect 159114 39922 159170 39978
rect 159238 39922 159294 39978
rect 159362 39922 159418 39978
rect 159486 39922 159542 39978
rect 132114 28294 132170 28350
rect 132238 28294 132294 28350
rect 132362 28294 132418 28350
rect 132486 28294 132542 28350
rect 132114 28170 132170 28226
rect 132238 28170 132294 28226
rect 132362 28170 132418 28226
rect 132486 28170 132542 28226
rect 132114 28046 132170 28102
rect 132238 28046 132294 28102
rect 132362 28046 132418 28102
rect 132486 28046 132542 28102
rect 132114 27922 132170 27978
rect 132238 27922 132294 27978
rect 132362 27922 132418 27978
rect 132486 27922 132542 27978
rect 132114 10294 132170 10350
rect 132238 10294 132294 10350
rect 132362 10294 132418 10350
rect 132486 10294 132542 10350
rect 132114 10170 132170 10226
rect 132238 10170 132294 10226
rect 132362 10170 132418 10226
rect 132486 10170 132542 10226
rect 132114 10046 132170 10102
rect 132238 10046 132294 10102
rect 132362 10046 132418 10102
rect 132486 10046 132542 10102
rect 132114 9922 132170 9978
rect 132238 9922 132294 9978
rect 132362 9922 132418 9978
rect 132486 9922 132542 9978
rect 132114 -1176 132170 -1120
rect 132238 -1176 132294 -1120
rect 132362 -1176 132418 -1120
rect 132486 -1176 132542 -1120
rect 132114 -1300 132170 -1244
rect 132238 -1300 132294 -1244
rect 132362 -1300 132418 -1244
rect 132486 -1300 132542 -1244
rect 132114 -1424 132170 -1368
rect 132238 -1424 132294 -1368
rect 132362 -1424 132418 -1368
rect 132486 -1424 132542 -1368
rect 132114 -1548 132170 -1492
rect 132238 -1548 132294 -1492
rect 132362 -1548 132418 -1492
rect 132486 -1548 132542 -1492
rect 159114 22294 159170 22350
rect 159238 22294 159294 22350
rect 159362 22294 159418 22350
rect 159486 22294 159542 22350
rect 159114 22170 159170 22226
rect 159238 22170 159294 22226
rect 159362 22170 159418 22226
rect 159486 22170 159542 22226
rect 159114 22046 159170 22102
rect 159238 22046 159294 22102
rect 159362 22046 159418 22102
rect 159486 22046 159542 22102
rect 159114 21922 159170 21978
rect 159238 21922 159294 21978
rect 159362 21922 159418 21978
rect 159486 21922 159542 21978
rect 159114 4294 159170 4350
rect 159238 4294 159294 4350
rect 159362 4294 159418 4350
rect 159486 4294 159542 4350
rect 159114 4170 159170 4226
rect 159238 4170 159294 4226
rect 159362 4170 159418 4226
rect 159486 4170 159542 4226
rect 159114 4046 159170 4102
rect 159238 4046 159294 4102
rect 159362 4046 159418 4102
rect 159486 4046 159542 4102
rect 159114 3922 159170 3978
rect 159238 3922 159294 3978
rect 159362 3922 159418 3978
rect 159486 3922 159542 3978
rect 159114 -216 159170 -160
rect 159238 -216 159294 -160
rect 159362 -216 159418 -160
rect 159486 -216 159542 -160
rect 159114 -340 159170 -284
rect 159238 -340 159294 -284
rect 159362 -340 159418 -284
rect 159486 -340 159542 -284
rect 159114 -464 159170 -408
rect 159238 -464 159294 -408
rect 159362 -464 159418 -408
rect 159486 -464 159542 -408
rect 159114 -588 159170 -532
rect 159238 -588 159294 -532
rect 159362 -588 159418 -532
rect 159486 -588 159542 -532
rect 162834 46294 162890 46350
rect 162958 46294 163014 46350
rect 163082 46294 163138 46350
rect 163206 46294 163262 46350
rect 162834 46170 162890 46226
rect 162958 46170 163014 46226
rect 163082 46170 163138 46226
rect 163206 46170 163262 46226
rect 162834 46046 162890 46102
rect 162958 46046 163014 46102
rect 163082 46046 163138 46102
rect 163206 46046 163262 46102
rect 162834 45922 162890 45978
rect 162958 45922 163014 45978
rect 163082 45922 163138 45978
rect 163206 45922 163262 45978
rect 163878 46294 163934 46350
rect 164002 46294 164058 46350
rect 163878 46170 163934 46226
rect 164002 46170 164058 46226
rect 163878 46046 163934 46102
rect 164002 46046 164058 46102
rect 163878 45922 163934 45978
rect 164002 45922 164058 45978
rect 179238 40294 179294 40350
rect 179362 40294 179418 40350
rect 179238 40170 179294 40226
rect 179362 40170 179418 40226
rect 179238 40046 179294 40102
rect 179362 40046 179418 40102
rect 179238 39922 179294 39978
rect 179362 39922 179418 39978
rect 189834 40294 189890 40350
rect 189958 40294 190014 40350
rect 190082 40294 190138 40350
rect 190206 40294 190262 40350
rect 189834 40170 189890 40226
rect 189958 40170 190014 40226
rect 190082 40170 190138 40226
rect 190206 40170 190262 40226
rect 189834 40046 189890 40102
rect 189958 40046 190014 40102
rect 190082 40046 190138 40102
rect 190206 40046 190262 40102
rect 189834 39922 189890 39978
rect 189958 39922 190014 39978
rect 190082 39922 190138 39978
rect 190206 39922 190262 39978
rect 162834 28294 162890 28350
rect 162958 28294 163014 28350
rect 163082 28294 163138 28350
rect 163206 28294 163262 28350
rect 162834 28170 162890 28226
rect 162958 28170 163014 28226
rect 163082 28170 163138 28226
rect 163206 28170 163262 28226
rect 162834 28046 162890 28102
rect 162958 28046 163014 28102
rect 163082 28046 163138 28102
rect 163206 28046 163262 28102
rect 162834 27922 162890 27978
rect 162958 27922 163014 27978
rect 163082 27922 163138 27978
rect 163206 27922 163262 27978
rect 162834 10294 162890 10350
rect 162958 10294 163014 10350
rect 163082 10294 163138 10350
rect 163206 10294 163262 10350
rect 162834 10170 162890 10226
rect 162958 10170 163014 10226
rect 163082 10170 163138 10226
rect 163206 10170 163262 10226
rect 162834 10046 162890 10102
rect 162958 10046 163014 10102
rect 163082 10046 163138 10102
rect 163206 10046 163262 10102
rect 162834 9922 162890 9978
rect 162958 9922 163014 9978
rect 163082 9922 163138 9978
rect 163206 9922 163262 9978
rect 162834 -1176 162890 -1120
rect 162958 -1176 163014 -1120
rect 163082 -1176 163138 -1120
rect 163206 -1176 163262 -1120
rect 162834 -1300 162890 -1244
rect 162958 -1300 163014 -1244
rect 163082 -1300 163138 -1244
rect 163206 -1300 163262 -1244
rect 162834 -1424 162890 -1368
rect 162958 -1424 163014 -1368
rect 163082 -1424 163138 -1368
rect 163206 -1424 163262 -1368
rect 162834 -1548 162890 -1492
rect 162958 -1548 163014 -1492
rect 163082 -1548 163138 -1492
rect 163206 -1548 163262 -1492
rect 189834 22294 189890 22350
rect 189958 22294 190014 22350
rect 190082 22294 190138 22350
rect 190206 22294 190262 22350
rect 189834 22170 189890 22226
rect 189958 22170 190014 22226
rect 190082 22170 190138 22226
rect 190206 22170 190262 22226
rect 189834 22046 189890 22102
rect 189958 22046 190014 22102
rect 190082 22046 190138 22102
rect 190206 22046 190262 22102
rect 189834 21922 189890 21978
rect 189958 21922 190014 21978
rect 190082 21922 190138 21978
rect 190206 21922 190262 21978
rect 189834 4294 189890 4350
rect 189958 4294 190014 4350
rect 190082 4294 190138 4350
rect 190206 4294 190262 4350
rect 189834 4170 189890 4226
rect 189958 4170 190014 4226
rect 190082 4170 190138 4226
rect 190206 4170 190262 4226
rect 189834 4046 189890 4102
rect 189958 4046 190014 4102
rect 190082 4046 190138 4102
rect 190206 4046 190262 4102
rect 189834 3922 189890 3978
rect 189958 3922 190014 3978
rect 190082 3922 190138 3978
rect 190206 3922 190262 3978
rect 189834 -216 189890 -160
rect 189958 -216 190014 -160
rect 190082 -216 190138 -160
rect 190206 -216 190262 -160
rect 189834 -340 189890 -284
rect 189958 -340 190014 -284
rect 190082 -340 190138 -284
rect 190206 -340 190262 -284
rect 189834 -464 189890 -408
rect 189958 -464 190014 -408
rect 190082 -464 190138 -408
rect 190206 -464 190262 -408
rect 189834 -588 189890 -532
rect 189958 -588 190014 -532
rect 190082 -588 190138 -532
rect 190206 -588 190262 -532
rect 193554 118294 193610 118350
rect 193678 118294 193734 118350
rect 193802 118294 193858 118350
rect 193926 118294 193982 118350
rect 193554 118170 193610 118226
rect 193678 118170 193734 118226
rect 193802 118170 193858 118226
rect 193926 118170 193982 118226
rect 193554 118046 193610 118102
rect 193678 118046 193734 118102
rect 193802 118046 193858 118102
rect 193926 118046 193982 118102
rect 193554 117922 193610 117978
rect 193678 117922 193734 117978
rect 193802 117922 193858 117978
rect 193926 117922 193982 117978
rect 193554 100294 193610 100350
rect 193678 100294 193734 100350
rect 193802 100294 193858 100350
rect 193926 100294 193982 100350
rect 193554 100170 193610 100226
rect 193678 100170 193734 100226
rect 193802 100170 193858 100226
rect 193926 100170 193982 100226
rect 193554 100046 193610 100102
rect 193678 100046 193734 100102
rect 193802 100046 193858 100102
rect 193926 100046 193982 100102
rect 193554 99922 193610 99978
rect 193678 99922 193734 99978
rect 193802 99922 193858 99978
rect 193926 99922 193982 99978
rect 193554 82294 193610 82350
rect 193678 82294 193734 82350
rect 193802 82294 193858 82350
rect 193926 82294 193982 82350
rect 193554 82170 193610 82226
rect 193678 82170 193734 82226
rect 193802 82170 193858 82226
rect 193926 82170 193982 82226
rect 193554 82046 193610 82102
rect 193678 82046 193734 82102
rect 193802 82046 193858 82102
rect 193926 82046 193982 82102
rect 193554 81922 193610 81978
rect 193678 81922 193734 81978
rect 193802 81922 193858 81978
rect 193926 81922 193982 81978
rect 193554 64294 193610 64350
rect 193678 64294 193734 64350
rect 193802 64294 193858 64350
rect 193926 64294 193982 64350
rect 193554 64170 193610 64226
rect 193678 64170 193734 64226
rect 193802 64170 193858 64226
rect 193926 64170 193982 64226
rect 193554 64046 193610 64102
rect 193678 64046 193734 64102
rect 193802 64046 193858 64102
rect 193926 64046 193982 64102
rect 193554 63922 193610 63978
rect 193678 63922 193734 63978
rect 193802 63922 193858 63978
rect 193926 63922 193982 63978
rect 193554 46294 193610 46350
rect 193678 46294 193734 46350
rect 193802 46294 193858 46350
rect 193926 46294 193982 46350
rect 193554 46170 193610 46226
rect 193678 46170 193734 46226
rect 193802 46170 193858 46226
rect 193926 46170 193982 46226
rect 193554 46046 193610 46102
rect 193678 46046 193734 46102
rect 193802 46046 193858 46102
rect 193926 46046 193982 46102
rect 193554 45922 193610 45978
rect 193678 45922 193734 45978
rect 193802 45922 193858 45978
rect 193926 45922 193982 45978
rect 193554 28294 193610 28350
rect 193678 28294 193734 28350
rect 193802 28294 193858 28350
rect 193926 28294 193982 28350
rect 193554 28170 193610 28226
rect 193678 28170 193734 28226
rect 193802 28170 193858 28226
rect 193926 28170 193982 28226
rect 193554 28046 193610 28102
rect 193678 28046 193734 28102
rect 193802 28046 193858 28102
rect 193926 28046 193982 28102
rect 193554 27922 193610 27978
rect 193678 27922 193734 27978
rect 193802 27922 193858 27978
rect 193926 27922 193982 27978
rect 193554 10294 193610 10350
rect 193678 10294 193734 10350
rect 193802 10294 193858 10350
rect 193926 10294 193982 10350
rect 193554 10170 193610 10226
rect 193678 10170 193734 10226
rect 193802 10170 193858 10226
rect 193926 10170 193982 10226
rect 193554 10046 193610 10102
rect 193678 10046 193734 10102
rect 193802 10046 193858 10102
rect 193926 10046 193982 10102
rect 193554 9922 193610 9978
rect 193678 9922 193734 9978
rect 193802 9922 193858 9978
rect 193926 9922 193982 9978
rect 210518 562294 210574 562350
rect 210642 562294 210698 562350
rect 210518 562170 210574 562226
rect 210642 562170 210698 562226
rect 210518 562046 210574 562102
rect 210642 562046 210698 562102
rect 210518 561922 210574 561978
rect 210642 561922 210698 561978
rect 220554 562294 220610 562350
rect 220678 562294 220734 562350
rect 220802 562294 220858 562350
rect 220926 562294 220982 562350
rect 220554 562170 220610 562226
rect 220678 562170 220734 562226
rect 220802 562170 220858 562226
rect 220926 562170 220982 562226
rect 220554 562046 220610 562102
rect 220678 562046 220734 562102
rect 220802 562046 220858 562102
rect 220926 562046 220982 562102
rect 220554 561922 220610 561978
rect 220678 561922 220734 561978
rect 220802 561922 220858 561978
rect 220926 561922 220982 561978
rect 201628 555182 201684 555238
rect 204876 533402 204932 533458
rect 210518 544294 210574 544350
rect 210642 544294 210698 544350
rect 210518 544170 210574 544226
rect 210642 544170 210698 544226
rect 210518 544046 210574 544102
rect 210642 544046 210698 544102
rect 210518 543922 210574 543978
rect 210642 543922 210698 543978
rect 224274 598116 224330 598172
rect 224398 598116 224454 598172
rect 224522 598116 224578 598172
rect 224646 598116 224702 598172
rect 224274 597992 224330 598048
rect 224398 597992 224454 598048
rect 224522 597992 224578 598048
rect 224646 597992 224702 598048
rect 224274 597868 224330 597924
rect 224398 597868 224454 597924
rect 224522 597868 224578 597924
rect 224646 597868 224702 597924
rect 224274 597744 224330 597800
rect 224398 597744 224454 597800
rect 224522 597744 224578 597800
rect 224646 597744 224702 597800
rect 224274 586294 224330 586350
rect 224398 586294 224454 586350
rect 224522 586294 224578 586350
rect 224646 586294 224702 586350
rect 224274 586170 224330 586226
rect 224398 586170 224454 586226
rect 224522 586170 224578 586226
rect 224646 586170 224702 586226
rect 224274 586046 224330 586102
rect 224398 586046 224454 586102
rect 224522 586046 224578 586102
rect 224646 586046 224702 586102
rect 224274 585922 224330 585978
rect 224398 585922 224454 585978
rect 224522 585922 224578 585978
rect 224646 585922 224702 585978
rect 224274 568294 224330 568350
rect 224398 568294 224454 568350
rect 224522 568294 224578 568350
rect 224646 568294 224702 568350
rect 224274 568170 224330 568226
rect 224398 568170 224454 568226
rect 224522 568170 224578 568226
rect 224646 568170 224702 568226
rect 224274 568046 224330 568102
rect 224398 568046 224454 568102
rect 224522 568046 224578 568102
rect 224646 568046 224702 568102
rect 224274 567922 224330 567978
rect 224398 567922 224454 567978
rect 224522 567922 224578 567978
rect 224646 567922 224702 567978
rect 251274 597156 251330 597212
rect 251398 597156 251454 597212
rect 251522 597156 251578 597212
rect 251646 597156 251702 597212
rect 251274 597032 251330 597088
rect 251398 597032 251454 597088
rect 251522 597032 251578 597088
rect 251646 597032 251702 597088
rect 251274 596908 251330 596964
rect 251398 596908 251454 596964
rect 251522 596908 251578 596964
rect 251646 596908 251702 596964
rect 251274 596784 251330 596840
rect 251398 596784 251454 596840
rect 251522 596784 251578 596840
rect 251646 596784 251702 596840
rect 251274 580294 251330 580350
rect 251398 580294 251454 580350
rect 251522 580294 251578 580350
rect 251646 580294 251702 580350
rect 251274 580170 251330 580226
rect 251398 580170 251454 580226
rect 251522 580170 251578 580226
rect 251646 580170 251702 580226
rect 251274 580046 251330 580102
rect 251398 580046 251454 580102
rect 251522 580046 251578 580102
rect 251646 580046 251702 580102
rect 251274 579922 251330 579978
rect 251398 579922 251454 579978
rect 251522 579922 251578 579978
rect 251646 579922 251702 579978
rect 241238 562294 241294 562350
rect 241362 562294 241418 562350
rect 241238 562170 241294 562226
rect 241362 562170 241418 562226
rect 241238 562046 241294 562102
rect 241362 562046 241418 562102
rect 241238 561922 241294 561978
rect 241362 561922 241418 561978
rect 251274 562294 251330 562350
rect 251398 562294 251454 562350
rect 251522 562294 251578 562350
rect 251646 562294 251702 562350
rect 251274 562170 251330 562226
rect 251398 562170 251454 562226
rect 251522 562170 251578 562226
rect 251646 562170 251702 562226
rect 251274 562046 251330 562102
rect 251398 562046 251454 562102
rect 251522 562046 251578 562102
rect 251646 562046 251702 562102
rect 251274 561922 251330 561978
rect 251398 561922 251454 561978
rect 251522 561922 251578 561978
rect 251646 561922 251702 561978
rect 225878 550294 225934 550350
rect 226002 550294 226058 550350
rect 225878 550170 225934 550226
rect 226002 550170 226058 550226
rect 225878 550046 225934 550102
rect 226002 550046 226058 550102
rect 225878 549922 225934 549978
rect 226002 549922 226058 549978
rect 220554 544294 220610 544350
rect 220678 544294 220734 544350
rect 220802 544294 220858 544350
rect 220926 544294 220982 544350
rect 220554 544170 220610 544226
rect 220678 544170 220734 544226
rect 220802 544170 220858 544226
rect 220926 544170 220982 544226
rect 220554 544046 220610 544102
rect 220678 544046 220734 544102
rect 220802 544046 220858 544102
rect 220926 544046 220982 544102
rect 241238 544294 241294 544350
rect 241362 544294 241418 544350
rect 241238 544170 241294 544226
rect 241362 544170 241418 544226
rect 241238 544046 241294 544102
rect 241362 544046 241418 544102
rect 220554 543922 220610 543978
rect 220678 543922 220734 543978
rect 220802 543922 220858 543978
rect 220926 543922 220982 543978
rect 220554 526294 220610 526350
rect 220678 526294 220734 526350
rect 220802 526294 220858 526350
rect 220926 526294 220982 526350
rect 220554 526170 220610 526226
rect 220678 526170 220734 526226
rect 220802 526170 220858 526226
rect 220926 526170 220982 526226
rect 220554 526046 220610 526102
rect 220678 526046 220734 526102
rect 220802 526046 220858 526102
rect 220926 526046 220982 526102
rect 220554 525922 220610 525978
rect 220678 525922 220734 525978
rect 220802 525922 220858 525978
rect 220926 525922 220982 525978
rect 220554 508294 220610 508350
rect 220678 508294 220734 508350
rect 220802 508294 220858 508350
rect 220926 508294 220982 508350
rect 220554 508170 220610 508226
rect 220678 508170 220734 508226
rect 220802 508170 220858 508226
rect 220926 508170 220982 508226
rect 220554 508046 220610 508102
rect 220678 508046 220734 508102
rect 220802 508046 220858 508102
rect 220926 508046 220982 508102
rect 220554 507922 220610 507978
rect 220678 507922 220734 507978
rect 220802 507922 220858 507978
rect 220926 507922 220982 507978
rect 210518 490294 210574 490350
rect 210642 490294 210698 490350
rect 210518 490170 210574 490226
rect 210642 490170 210698 490226
rect 210518 490046 210574 490102
rect 210642 490046 210698 490102
rect 210518 489922 210574 489978
rect 210642 489922 210698 489978
rect 220554 490294 220610 490350
rect 220678 490294 220734 490350
rect 220802 490294 220858 490350
rect 220926 490294 220982 490350
rect 220554 490170 220610 490226
rect 220678 490170 220734 490226
rect 220802 490170 220858 490226
rect 220926 490170 220982 490226
rect 220554 490046 220610 490102
rect 220678 490046 220734 490102
rect 220802 490046 220858 490102
rect 220926 490046 220982 490102
rect 220554 489922 220610 489978
rect 220678 489922 220734 489978
rect 220802 489922 220858 489978
rect 220926 489922 220982 489978
rect 201628 483002 201684 483058
rect 206668 482300 206724 482338
rect 206668 482282 206724 482300
rect 206556 474542 206612 474598
rect 210518 472294 210574 472350
rect 210642 472294 210698 472350
rect 210518 472170 210574 472226
rect 210642 472170 210698 472226
rect 210518 472046 210574 472102
rect 210642 472046 210698 472102
rect 210518 471922 210574 471978
rect 210642 471922 210698 471978
rect 241238 543922 241294 543978
rect 241362 543922 241418 543978
rect 254994 598116 255050 598172
rect 255118 598116 255174 598172
rect 255242 598116 255298 598172
rect 255366 598116 255422 598172
rect 254994 597992 255050 598048
rect 255118 597992 255174 598048
rect 255242 597992 255298 598048
rect 255366 597992 255422 598048
rect 254994 597868 255050 597924
rect 255118 597868 255174 597924
rect 255242 597868 255298 597924
rect 255366 597868 255422 597924
rect 254994 597744 255050 597800
rect 255118 597744 255174 597800
rect 255242 597744 255298 597800
rect 255366 597744 255422 597800
rect 254994 586294 255050 586350
rect 255118 586294 255174 586350
rect 255242 586294 255298 586350
rect 255366 586294 255422 586350
rect 254994 586170 255050 586226
rect 255118 586170 255174 586226
rect 255242 586170 255298 586226
rect 255366 586170 255422 586226
rect 254994 586046 255050 586102
rect 255118 586046 255174 586102
rect 255242 586046 255298 586102
rect 255366 586046 255422 586102
rect 254994 585922 255050 585978
rect 255118 585922 255174 585978
rect 255242 585922 255298 585978
rect 255366 585922 255422 585978
rect 281994 597156 282050 597212
rect 282118 597156 282174 597212
rect 282242 597156 282298 597212
rect 282366 597156 282422 597212
rect 281994 597032 282050 597088
rect 282118 597032 282174 597088
rect 282242 597032 282298 597088
rect 282366 597032 282422 597088
rect 281994 596908 282050 596964
rect 282118 596908 282174 596964
rect 282242 596908 282298 596964
rect 282366 596908 282422 596964
rect 281994 596784 282050 596840
rect 282118 596784 282174 596840
rect 282242 596784 282298 596840
rect 282366 596784 282422 596840
rect 281994 580294 282050 580350
rect 282118 580294 282174 580350
rect 282242 580294 282298 580350
rect 282366 580294 282422 580350
rect 281994 580170 282050 580226
rect 282118 580170 282174 580226
rect 282242 580170 282298 580226
rect 282366 580170 282422 580226
rect 281994 580046 282050 580102
rect 282118 580046 282174 580102
rect 282242 580046 282298 580102
rect 282366 580046 282422 580102
rect 281994 579922 282050 579978
rect 282118 579922 282174 579978
rect 282242 579922 282298 579978
rect 282366 579922 282422 579978
rect 254994 568294 255050 568350
rect 255118 568294 255174 568350
rect 255242 568294 255298 568350
rect 255366 568294 255422 568350
rect 254994 568170 255050 568226
rect 255118 568170 255174 568226
rect 255242 568170 255298 568226
rect 255366 568170 255422 568226
rect 254994 568046 255050 568102
rect 255118 568046 255174 568102
rect 255242 568046 255298 568102
rect 255366 568046 255422 568102
rect 254994 567922 255050 567978
rect 255118 567922 255174 567978
rect 255242 567922 255298 567978
rect 255366 567922 255422 567978
rect 251274 544294 251330 544350
rect 251398 544294 251454 544350
rect 251522 544294 251578 544350
rect 251646 544294 251702 544350
rect 251274 544170 251330 544226
rect 251398 544170 251454 544226
rect 251522 544170 251578 544226
rect 251646 544170 251702 544226
rect 251274 544046 251330 544102
rect 251398 544046 251454 544102
rect 251522 544046 251578 544102
rect 251646 544046 251702 544102
rect 251274 543922 251330 543978
rect 251398 543922 251454 543978
rect 251522 543922 251578 543978
rect 251646 543922 251702 543978
rect 224274 532294 224330 532350
rect 224398 532294 224454 532350
rect 224522 532294 224578 532350
rect 224646 532294 224702 532350
rect 224274 532170 224330 532226
rect 224398 532170 224454 532226
rect 224522 532170 224578 532226
rect 224646 532170 224702 532226
rect 224274 532046 224330 532102
rect 224398 532046 224454 532102
rect 224522 532046 224578 532102
rect 224646 532046 224702 532102
rect 224274 531922 224330 531978
rect 224398 531922 224454 531978
rect 224522 531922 224578 531978
rect 224646 531922 224702 531978
rect 225878 532294 225934 532350
rect 226002 532294 226058 532350
rect 225878 532170 225934 532226
rect 226002 532170 226058 532226
rect 225878 532046 225934 532102
rect 226002 532046 226058 532102
rect 225878 531922 225934 531978
rect 226002 531922 226058 531978
rect 224274 514294 224330 514350
rect 224398 514294 224454 514350
rect 224522 514294 224578 514350
rect 224646 514294 224702 514350
rect 224274 514170 224330 514226
rect 224398 514170 224454 514226
rect 224522 514170 224578 514226
rect 224646 514170 224702 514226
rect 224274 514046 224330 514102
rect 224398 514046 224454 514102
rect 224522 514046 224578 514102
rect 224646 514046 224702 514102
rect 224274 513922 224330 513978
rect 224398 513922 224454 513978
rect 224522 513922 224578 513978
rect 224646 513922 224702 513978
rect 224274 496294 224330 496350
rect 224398 496294 224454 496350
rect 224522 496294 224578 496350
rect 224646 496294 224702 496350
rect 224274 496170 224330 496226
rect 224398 496170 224454 496226
rect 224522 496170 224578 496226
rect 224646 496170 224702 496226
rect 224274 496046 224330 496102
rect 224398 496046 224454 496102
rect 224522 496046 224578 496102
rect 224646 496046 224702 496102
rect 224274 495922 224330 495978
rect 224398 495922 224454 495978
rect 224522 495922 224578 495978
rect 224646 495922 224702 495978
rect 241238 490294 241294 490350
rect 241362 490294 241418 490350
rect 241238 490170 241294 490226
rect 241362 490170 241418 490226
rect 241238 490046 241294 490102
rect 241362 490046 241418 490102
rect 241238 489922 241294 489978
rect 241362 489922 241418 489978
rect 251274 526294 251330 526350
rect 251398 526294 251454 526350
rect 251522 526294 251578 526350
rect 251646 526294 251702 526350
rect 251274 526170 251330 526226
rect 251398 526170 251454 526226
rect 251522 526170 251578 526226
rect 251646 526170 251702 526226
rect 251274 526046 251330 526102
rect 251398 526046 251454 526102
rect 251522 526046 251578 526102
rect 251646 526046 251702 526102
rect 251274 525922 251330 525978
rect 251398 525922 251454 525978
rect 251522 525922 251578 525978
rect 251646 525922 251702 525978
rect 285714 598116 285770 598172
rect 285838 598116 285894 598172
rect 285962 598116 286018 598172
rect 286086 598116 286142 598172
rect 285714 597992 285770 598048
rect 285838 597992 285894 598048
rect 285962 597992 286018 598048
rect 286086 597992 286142 598048
rect 285714 597868 285770 597924
rect 285838 597868 285894 597924
rect 285962 597868 286018 597924
rect 286086 597868 286142 597924
rect 285714 597744 285770 597800
rect 285838 597744 285894 597800
rect 285962 597744 286018 597800
rect 286086 597744 286142 597800
rect 285714 586294 285770 586350
rect 285838 586294 285894 586350
rect 285962 586294 286018 586350
rect 286086 586294 286142 586350
rect 285714 586170 285770 586226
rect 285838 586170 285894 586226
rect 285962 586170 286018 586226
rect 286086 586170 286142 586226
rect 285714 586046 285770 586102
rect 285838 586046 285894 586102
rect 285962 586046 286018 586102
rect 286086 586046 286142 586102
rect 285714 585922 285770 585978
rect 285838 585922 285894 585978
rect 285962 585922 286018 585978
rect 286086 585922 286142 585978
rect 312714 597156 312770 597212
rect 312838 597156 312894 597212
rect 312962 597156 313018 597212
rect 313086 597156 313142 597212
rect 312714 597032 312770 597088
rect 312838 597032 312894 597088
rect 312962 597032 313018 597088
rect 313086 597032 313142 597088
rect 312714 596908 312770 596964
rect 312838 596908 312894 596964
rect 312962 596908 313018 596964
rect 313086 596908 313142 596964
rect 312714 596784 312770 596840
rect 312838 596784 312894 596840
rect 312962 596784 313018 596840
rect 313086 596784 313142 596840
rect 312714 580294 312770 580350
rect 312838 580294 312894 580350
rect 312962 580294 313018 580350
rect 313086 580294 313142 580350
rect 312714 580170 312770 580226
rect 312838 580170 312894 580226
rect 312962 580170 313018 580226
rect 313086 580170 313142 580226
rect 312714 580046 312770 580102
rect 312838 580046 312894 580102
rect 312962 580046 313018 580102
rect 313086 580046 313142 580102
rect 312714 579922 312770 579978
rect 312838 579922 312894 579978
rect 312962 579922 313018 579978
rect 313086 579922 313142 579978
rect 290444 569582 290500 569638
rect 285714 568294 285770 568350
rect 285838 568294 285894 568350
rect 285962 568294 286018 568350
rect 286086 568294 286142 568350
rect 285714 568170 285770 568226
rect 285838 568170 285894 568226
rect 285962 568170 286018 568226
rect 286086 568170 286142 568226
rect 285714 568046 285770 568102
rect 285838 568046 285894 568102
rect 285962 568046 286018 568102
rect 286086 568046 286142 568102
rect 285714 567922 285770 567978
rect 285838 567922 285894 567978
rect 285962 567922 286018 567978
rect 286086 567922 286142 567978
rect 316434 598116 316490 598172
rect 316558 598116 316614 598172
rect 316682 598116 316738 598172
rect 316806 598116 316862 598172
rect 316434 597992 316490 598048
rect 316558 597992 316614 598048
rect 316682 597992 316738 598048
rect 316806 597992 316862 598048
rect 316434 597868 316490 597924
rect 316558 597868 316614 597924
rect 316682 597868 316738 597924
rect 316806 597868 316862 597924
rect 316434 597744 316490 597800
rect 316558 597744 316614 597800
rect 316682 597744 316738 597800
rect 316806 597744 316862 597800
rect 316434 586294 316490 586350
rect 316558 586294 316614 586350
rect 316682 586294 316738 586350
rect 316806 586294 316862 586350
rect 316434 586170 316490 586226
rect 316558 586170 316614 586226
rect 316682 586170 316738 586226
rect 316806 586170 316862 586226
rect 316434 586046 316490 586102
rect 316558 586046 316614 586102
rect 316682 586046 316738 586102
rect 316806 586046 316862 586102
rect 316434 585922 316490 585978
rect 316558 585922 316614 585978
rect 316682 585922 316738 585978
rect 316806 585922 316862 585978
rect 343434 597156 343490 597212
rect 343558 597156 343614 597212
rect 343682 597156 343738 597212
rect 343806 597156 343862 597212
rect 343434 597032 343490 597088
rect 343558 597032 343614 597088
rect 343682 597032 343738 597088
rect 343806 597032 343862 597088
rect 343434 596908 343490 596964
rect 343558 596908 343614 596964
rect 343682 596908 343738 596964
rect 343806 596908 343862 596964
rect 343434 596784 343490 596840
rect 343558 596784 343614 596840
rect 343682 596784 343738 596840
rect 343806 596784 343862 596840
rect 343434 580294 343490 580350
rect 343558 580294 343614 580350
rect 343682 580294 343738 580350
rect 343806 580294 343862 580350
rect 343434 580170 343490 580226
rect 343558 580170 343614 580226
rect 343682 580170 343738 580226
rect 343806 580170 343862 580226
rect 343434 580046 343490 580102
rect 343558 580046 343614 580102
rect 343682 580046 343738 580102
rect 343806 580046 343862 580102
rect 343434 579922 343490 579978
rect 343558 579922 343614 579978
rect 343682 579922 343738 579978
rect 343806 579922 343862 579978
rect 316434 568294 316490 568350
rect 316558 568294 316614 568350
rect 316682 568294 316738 568350
rect 316806 568294 316862 568350
rect 316434 568170 316490 568226
rect 316558 568170 316614 568226
rect 316682 568170 316738 568226
rect 316806 568170 316862 568226
rect 316434 568046 316490 568102
rect 316558 568046 316614 568102
rect 316682 568046 316738 568102
rect 316806 568046 316862 568102
rect 316434 567922 316490 567978
rect 316558 567922 316614 567978
rect 316682 567922 316738 567978
rect 316806 567922 316862 567978
rect 330764 571228 330820 571258
rect 330764 571202 330820 571228
rect 333452 569582 333508 569638
rect 289324 566882 289380 566938
rect 272518 562294 272574 562350
rect 272642 562294 272698 562350
rect 272518 562170 272574 562226
rect 272642 562170 272698 562226
rect 272518 562046 272574 562102
rect 272642 562046 272698 562102
rect 272518 561922 272574 561978
rect 272642 561922 272698 561978
rect 303238 562294 303294 562350
rect 303362 562294 303418 562350
rect 303238 562170 303294 562226
rect 303362 562170 303418 562226
rect 303238 562046 303294 562102
rect 303362 562046 303418 562102
rect 303238 561922 303294 561978
rect 303362 561922 303418 561978
rect 254994 550294 255050 550350
rect 255118 550294 255174 550350
rect 255242 550294 255298 550350
rect 255366 550294 255422 550350
rect 254994 550170 255050 550226
rect 255118 550170 255174 550226
rect 255242 550170 255298 550226
rect 255366 550170 255422 550226
rect 254994 550046 255050 550102
rect 255118 550046 255174 550102
rect 255242 550046 255298 550102
rect 255366 550046 255422 550102
rect 254994 549922 255050 549978
rect 255118 549922 255174 549978
rect 255242 549922 255298 549978
rect 255366 549922 255422 549978
rect 254994 532294 255050 532350
rect 255118 532294 255174 532350
rect 255242 532294 255298 532350
rect 255366 532294 255422 532350
rect 254994 532170 255050 532226
rect 255118 532170 255174 532226
rect 255242 532170 255298 532226
rect 255366 532170 255422 532226
rect 254994 532046 255050 532102
rect 255118 532046 255174 532102
rect 255242 532046 255298 532102
rect 255366 532046 255422 532102
rect 254994 531922 255050 531978
rect 255118 531922 255174 531978
rect 255242 531922 255298 531978
rect 255366 531922 255422 531978
rect 251274 508294 251330 508350
rect 251398 508294 251454 508350
rect 251522 508294 251578 508350
rect 251646 508294 251702 508350
rect 251274 508170 251330 508226
rect 251398 508170 251454 508226
rect 251522 508170 251578 508226
rect 251646 508170 251702 508226
rect 251274 508046 251330 508102
rect 251398 508046 251454 508102
rect 251522 508046 251578 508102
rect 251646 508046 251702 508102
rect 251274 507922 251330 507978
rect 251398 507922 251454 507978
rect 251522 507922 251578 507978
rect 251646 507922 251702 507978
rect 251274 490294 251330 490350
rect 251398 490294 251454 490350
rect 251522 490294 251578 490350
rect 251646 490294 251702 490350
rect 251274 490170 251330 490226
rect 251398 490170 251454 490226
rect 251522 490170 251578 490226
rect 251646 490170 251702 490226
rect 251274 490046 251330 490102
rect 251398 490046 251454 490102
rect 251522 490046 251578 490102
rect 251646 490046 251702 490102
rect 251274 489922 251330 489978
rect 251398 489922 251454 489978
rect 251522 489922 251578 489978
rect 251646 489922 251702 489978
rect 247996 482282 248052 482338
rect 225878 478294 225934 478350
rect 226002 478294 226058 478350
rect 225878 478170 225934 478226
rect 226002 478170 226058 478226
rect 225878 478046 225934 478102
rect 226002 478046 226058 478102
rect 225878 477922 225934 477978
rect 226002 477922 226058 477978
rect 223356 474542 223412 474598
rect 223356 473642 223412 473698
rect 220554 472294 220610 472350
rect 220678 472294 220734 472350
rect 220802 472294 220858 472350
rect 220926 472294 220982 472350
rect 220554 472170 220610 472226
rect 220678 472170 220734 472226
rect 220802 472170 220858 472226
rect 220926 472170 220982 472226
rect 220554 472046 220610 472102
rect 220678 472046 220734 472102
rect 220802 472046 220858 472102
rect 220926 472046 220982 472102
rect 220554 471922 220610 471978
rect 220678 471922 220734 471978
rect 220802 471922 220858 471978
rect 220926 471922 220982 471978
rect 220554 454294 220610 454350
rect 220678 454294 220734 454350
rect 220802 454294 220858 454350
rect 220926 454294 220982 454350
rect 220554 454170 220610 454226
rect 220678 454170 220734 454226
rect 220802 454170 220858 454226
rect 220926 454170 220982 454226
rect 220554 454046 220610 454102
rect 220678 454046 220734 454102
rect 220802 454046 220858 454102
rect 220926 454046 220982 454102
rect 220554 453922 220610 453978
rect 220678 453922 220734 453978
rect 220802 453922 220858 453978
rect 220926 453922 220982 453978
rect 220554 436294 220610 436350
rect 220678 436294 220734 436350
rect 220802 436294 220858 436350
rect 220926 436294 220982 436350
rect 220554 436170 220610 436226
rect 220678 436170 220734 436226
rect 220802 436170 220858 436226
rect 220926 436170 220982 436226
rect 220554 436046 220610 436102
rect 220678 436046 220734 436102
rect 220802 436046 220858 436102
rect 220926 436046 220982 436102
rect 220554 435922 220610 435978
rect 220678 435922 220734 435978
rect 220802 435922 220858 435978
rect 220926 435922 220982 435978
rect 210518 418294 210574 418350
rect 210642 418294 210698 418350
rect 210518 418170 210574 418226
rect 210642 418170 210698 418226
rect 210518 418046 210574 418102
rect 210642 418046 210698 418102
rect 210518 417922 210574 417978
rect 210642 417922 210698 417978
rect 241238 472294 241294 472350
rect 241362 472294 241418 472350
rect 241238 472170 241294 472226
rect 241362 472170 241418 472226
rect 241238 472046 241294 472102
rect 241362 472046 241418 472102
rect 241238 471922 241294 471978
rect 241362 471922 241418 471978
rect 249452 473822 249508 473878
rect 254994 514294 255050 514350
rect 255118 514294 255174 514350
rect 255242 514294 255298 514350
rect 255366 514294 255422 514350
rect 254994 514170 255050 514226
rect 255118 514170 255174 514226
rect 255242 514170 255298 514226
rect 255366 514170 255422 514226
rect 254994 514046 255050 514102
rect 255118 514046 255174 514102
rect 255242 514046 255298 514102
rect 255366 514046 255422 514102
rect 254994 513922 255050 513978
rect 255118 513922 255174 513978
rect 255242 513922 255298 513978
rect 255366 513922 255422 513978
rect 254994 496294 255050 496350
rect 255118 496294 255174 496350
rect 255242 496294 255298 496350
rect 255366 496294 255422 496350
rect 254994 496170 255050 496226
rect 255118 496170 255174 496226
rect 255242 496170 255298 496226
rect 255366 496170 255422 496226
rect 254994 496046 255050 496102
rect 255118 496046 255174 496102
rect 255242 496046 255298 496102
rect 255366 496046 255422 496102
rect 254994 495922 255050 495978
rect 255118 495922 255174 495978
rect 255242 495922 255298 495978
rect 255366 495922 255422 495978
rect 254994 478294 255050 478350
rect 255118 478294 255174 478350
rect 255242 478294 255298 478350
rect 255366 478294 255422 478350
rect 254994 478170 255050 478226
rect 255118 478170 255174 478226
rect 255242 478170 255298 478226
rect 255366 478170 255422 478226
rect 254994 478046 255050 478102
rect 255118 478046 255174 478102
rect 255242 478046 255298 478102
rect 255366 478046 255422 478102
rect 254994 477922 255050 477978
rect 255118 477922 255174 477978
rect 255242 477922 255298 477978
rect 255366 477922 255422 477978
rect 251274 472294 251330 472350
rect 251398 472294 251454 472350
rect 251522 472294 251578 472350
rect 251646 472294 251702 472350
rect 251274 472170 251330 472226
rect 251398 472170 251454 472226
rect 251522 472170 251578 472226
rect 251646 472170 251702 472226
rect 251274 472046 251330 472102
rect 251398 472046 251454 472102
rect 251522 472046 251578 472102
rect 251646 472046 251702 472102
rect 251274 471922 251330 471978
rect 251398 471922 251454 471978
rect 251522 471922 251578 471978
rect 251646 471922 251702 471978
rect 249564 466082 249620 466138
rect 224274 460294 224330 460350
rect 224398 460294 224454 460350
rect 224522 460294 224578 460350
rect 224646 460294 224702 460350
rect 224274 460170 224330 460226
rect 224398 460170 224454 460226
rect 224522 460170 224578 460226
rect 224646 460170 224702 460226
rect 224274 460046 224330 460102
rect 224398 460046 224454 460102
rect 224522 460046 224578 460102
rect 224646 460046 224702 460102
rect 224274 459922 224330 459978
rect 224398 459922 224454 459978
rect 224522 459922 224578 459978
rect 224646 459922 224702 459978
rect 225878 460294 225934 460350
rect 226002 460294 226058 460350
rect 225878 460170 225934 460226
rect 226002 460170 226058 460226
rect 225878 460046 225934 460102
rect 226002 460046 226058 460102
rect 225878 459922 225934 459978
rect 226002 459922 226058 459978
rect 251274 454294 251330 454350
rect 251398 454294 251454 454350
rect 251522 454294 251578 454350
rect 251646 454294 251702 454350
rect 251274 454170 251330 454226
rect 251398 454170 251454 454226
rect 251522 454170 251578 454226
rect 251646 454170 251702 454226
rect 251274 454046 251330 454102
rect 251398 454046 251454 454102
rect 251522 454046 251578 454102
rect 251646 454046 251702 454102
rect 251274 453922 251330 453978
rect 251398 453922 251454 453978
rect 251522 453922 251578 453978
rect 251646 453922 251702 453978
rect 224274 442294 224330 442350
rect 224398 442294 224454 442350
rect 224522 442294 224578 442350
rect 224646 442294 224702 442350
rect 224274 442170 224330 442226
rect 224398 442170 224454 442226
rect 224522 442170 224578 442226
rect 224646 442170 224702 442226
rect 224274 442046 224330 442102
rect 224398 442046 224454 442102
rect 224522 442046 224578 442102
rect 224646 442046 224702 442102
rect 224274 441922 224330 441978
rect 224398 441922 224454 441978
rect 224522 441922 224578 441978
rect 224646 441922 224702 441978
rect 220554 418294 220610 418350
rect 220678 418294 220734 418350
rect 220802 418294 220858 418350
rect 220926 418294 220982 418350
rect 220554 418170 220610 418226
rect 220678 418170 220734 418226
rect 220802 418170 220858 418226
rect 220926 418170 220982 418226
rect 220554 418046 220610 418102
rect 220678 418046 220734 418102
rect 220802 418046 220858 418102
rect 220926 418046 220982 418102
rect 220554 417922 220610 417978
rect 220678 417922 220734 417978
rect 220802 417922 220858 417978
rect 220926 417922 220982 417978
rect 206668 414988 206724 415018
rect 206668 414962 206724 414988
rect 201628 412442 201684 412498
rect 204764 411722 204820 411778
rect 204988 407042 205044 407098
rect 204988 404162 205044 404218
rect 204988 402902 205044 402958
rect 210518 400294 210574 400350
rect 210642 400294 210698 400350
rect 210518 400170 210574 400226
rect 210642 400170 210698 400226
rect 210518 400046 210574 400102
rect 210642 400046 210698 400102
rect 210518 399922 210574 399978
rect 210642 399922 210698 399978
rect 220554 400294 220610 400350
rect 220678 400294 220734 400350
rect 220802 400294 220858 400350
rect 220926 400294 220982 400350
rect 220554 400170 220610 400226
rect 220678 400170 220734 400226
rect 220802 400170 220858 400226
rect 220926 400170 220982 400226
rect 220554 400046 220610 400102
rect 220678 400046 220734 400102
rect 220802 400046 220858 400102
rect 220926 400046 220982 400102
rect 220554 399922 220610 399978
rect 220678 399922 220734 399978
rect 220802 399922 220858 399978
rect 220926 399922 220982 399978
rect 220554 382294 220610 382350
rect 220678 382294 220734 382350
rect 220802 382294 220858 382350
rect 220926 382294 220982 382350
rect 220554 382170 220610 382226
rect 220678 382170 220734 382226
rect 220802 382170 220858 382226
rect 220926 382170 220982 382226
rect 220554 382046 220610 382102
rect 220678 382046 220734 382102
rect 220802 382046 220858 382102
rect 220926 382046 220982 382102
rect 220554 381922 220610 381978
rect 220678 381922 220734 381978
rect 220802 381922 220858 381978
rect 220926 381922 220982 381978
rect 220554 364294 220610 364350
rect 220678 364294 220734 364350
rect 220802 364294 220858 364350
rect 220926 364294 220982 364350
rect 220554 364170 220610 364226
rect 220678 364170 220734 364226
rect 220802 364170 220858 364226
rect 220926 364170 220982 364226
rect 220554 364046 220610 364102
rect 220678 364046 220734 364102
rect 220802 364046 220858 364102
rect 220926 364046 220982 364102
rect 220554 363922 220610 363978
rect 220678 363922 220734 363978
rect 220802 363922 220858 363978
rect 220926 363922 220982 363978
rect 201292 341162 201348 341218
rect 203084 348542 203140 348598
rect 205996 349442 206052 349498
rect 204876 324062 204932 324118
rect 210518 346294 210574 346350
rect 210642 346294 210698 346350
rect 210518 346170 210574 346226
rect 210642 346170 210698 346226
rect 210518 346046 210574 346102
rect 210642 346046 210698 346102
rect 210518 345922 210574 345978
rect 210642 345922 210698 345978
rect 220554 346294 220610 346350
rect 220678 346294 220734 346350
rect 220802 346294 220858 346350
rect 220926 346294 220982 346350
rect 220554 346170 220610 346226
rect 220678 346170 220734 346226
rect 220802 346170 220858 346226
rect 220926 346170 220982 346226
rect 220554 346046 220610 346102
rect 220678 346046 220734 346102
rect 220802 346046 220858 346102
rect 220926 346046 220982 346102
rect 220554 345922 220610 345978
rect 220678 345922 220734 345978
rect 220802 345922 220858 345978
rect 220926 345922 220982 345978
rect 210518 328294 210574 328350
rect 210642 328294 210698 328350
rect 210518 328170 210574 328226
rect 210642 328170 210698 328226
rect 210518 328046 210574 328102
rect 210642 328046 210698 328102
rect 210518 327922 210574 327978
rect 210642 327922 210698 327978
rect 220554 328294 220610 328350
rect 220678 328294 220734 328350
rect 220802 328294 220858 328350
rect 220926 328294 220982 328350
rect 220554 328170 220610 328226
rect 220678 328170 220734 328226
rect 220802 328170 220858 328226
rect 220926 328170 220982 328226
rect 220554 328046 220610 328102
rect 220678 328046 220734 328102
rect 220802 328046 220858 328102
rect 220926 328046 220982 328102
rect 220554 327922 220610 327978
rect 220678 327922 220734 327978
rect 220802 327922 220858 327978
rect 220926 327922 220982 327978
rect 206108 325502 206164 325558
rect 220554 310294 220610 310350
rect 220678 310294 220734 310350
rect 220802 310294 220858 310350
rect 220926 310294 220982 310350
rect 220554 310170 220610 310226
rect 220678 310170 220734 310226
rect 220802 310170 220858 310226
rect 220926 310170 220982 310226
rect 220554 310046 220610 310102
rect 220678 310046 220734 310102
rect 220802 310046 220858 310102
rect 220926 310046 220982 310102
rect 220554 309922 220610 309978
rect 220678 309922 220734 309978
rect 220802 309922 220858 309978
rect 220926 309922 220982 309978
rect 201628 271322 201684 271378
rect 220554 292294 220610 292350
rect 220678 292294 220734 292350
rect 220802 292294 220858 292350
rect 220926 292294 220982 292350
rect 220554 292170 220610 292226
rect 220678 292170 220734 292226
rect 220802 292170 220858 292226
rect 220926 292170 220982 292226
rect 220554 292046 220610 292102
rect 220678 292046 220734 292102
rect 220802 292046 220858 292102
rect 220926 292046 220982 292102
rect 220554 291922 220610 291978
rect 220678 291922 220734 291978
rect 220802 291922 220858 291978
rect 220926 291922 220982 291978
rect 210518 274294 210574 274350
rect 210642 274294 210698 274350
rect 210518 274170 210574 274226
rect 210642 274170 210698 274226
rect 210518 274046 210574 274102
rect 210642 274046 210698 274102
rect 210518 273922 210574 273978
rect 210642 273922 210698 273978
rect 220554 274294 220610 274350
rect 220678 274294 220734 274350
rect 220802 274294 220858 274350
rect 220926 274294 220982 274350
rect 220554 274170 220610 274226
rect 220678 274170 220734 274226
rect 220802 274170 220858 274226
rect 220926 274170 220982 274226
rect 220554 274046 220610 274102
rect 220678 274046 220734 274102
rect 220802 274046 220858 274102
rect 220926 274046 220982 274102
rect 220554 273922 220610 273978
rect 220678 273922 220734 273978
rect 220802 273922 220858 273978
rect 220926 273922 220982 273978
rect 206444 267182 206500 267238
rect 206332 266462 206388 266518
rect 206444 261604 206500 261658
rect 206444 261602 206500 261604
rect 210518 256294 210574 256350
rect 210642 256294 210698 256350
rect 210518 256170 210574 256226
rect 210642 256170 210698 256226
rect 210518 256046 210574 256102
rect 210642 256046 210698 256102
rect 210518 255922 210574 255978
rect 210642 255922 210698 255978
rect 220554 256294 220610 256350
rect 220678 256294 220734 256350
rect 220802 256294 220858 256350
rect 220926 256294 220982 256350
rect 220554 256170 220610 256226
rect 220678 256170 220734 256226
rect 220802 256170 220858 256226
rect 220926 256170 220982 256226
rect 220554 256046 220610 256102
rect 220678 256046 220734 256102
rect 220802 256046 220858 256102
rect 220926 256046 220982 256102
rect 220554 255922 220610 255978
rect 220678 255922 220734 255978
rect 220802 255922 220858 255978
rect 220926 255922 220982 255978
rect 220554 238294 220610 238350
rect 220678 238294 220734 238350
rect 220802 238294 220858 238350
rect 220926 238294 220982 238350
rect 220554 238170 220610 238226
rect 220678 238170 220734 238226
rect 220802 238170 220858 238226
rect 220926 238170 220982 238226
rect 220554 238046 220610 238102
rect 220678 238046 220734 238102
rect 220802 238046 220858 238102
rect 220926 238046 220982 238102
rect 220554 237922 220610 237978
rect 220678 237922 220734 237978
rect 220802 237922 220858 237978
rect 220926 237922 220982 237978
rect 202972 205802 203028 205858
rect 201628 198962 201684 199018
rect 220554 220294 220610 220350
rect 220678 220294 220734 220350
rect 220802 220294 220858 220350
rect 220926 220294 220982 220350
rect 220554 220170 220610 220226
rect 220678 220170 220734 220226
rect 220802 220170 220858 220226
rect 220926 220170 220982 220226
rect 220554 220046 220610 220102
rect 220678 220046 220734 220102
rect 220802 220046 220858 220102
rect 220926 220046 220982 220102
rect 220554 219922 220610 219978
rect 220678 219922 220734 219978
rect 220802 219922 220858 219978
rect 220926 219922 220982 219978
rect 210518 202294 210574 202350
rect 210642 202294 210698 202350
rect 210518 202170 210574 202226
rect 210642 202170 210698 202226
rect 210518 202046 210574 202102
rect 210642 202046 210698 202102
rect 210518 201922 210574 201978
rect 210642 201922 210698 201978
rect 220554 202294 220610 202350
rect 220678 202294 220734 202350
rect 220802 202294 220858 202350
rect 220926 202294 220982 202350
rect 220554 202170 220610 202226
rect 220678 202170 220734 202226
rect 220802 202170 220858 202226
rect 220926 202170 220982 202226
rect 220554 202046 220610 202102
rect 220678 202046 220734 202102
rect 220802 202046 220858 202102
rect 220926 202046 220982 202102
rect 220554 201922 220610 201978
rect 220678 201922 220734 201978
rect 220802 201922 220858 201978
rect 220926 201922 220982 201978
rect 205660 198242 205716 198298
rect 204988 195002 205044 195058
rect 210518 184294 210574 184350
rect 210642 184294 210698 184350
rect 210518 184170 210574 184226
rect 210642 184170 210698 184226
rect 210518 184046 210574 184102
rect 210642 184046 210698 184102
rect 210518 183922 210574 183978
rect 210642 183922 210698 183978
rect 220554 184294 220610 184350
rect 220678 184294 220734 184350
rect 220802 184294 220858 184350
rect 220926 184294 220982 184350
rect 220554 184170 220610 184226
rect 220678 184170 220734 184226
rect 220802 184170 220858 184226
rect 220926 184170 220982 184226
rect 220554 184046 220610 184102
rect 220678 184046 220734 184102
rect 220802 184046 220858 184102
rect 220926 184046 220982 184102
rect 220554 183922 220610 183978
rect 220678 183922 220734 183978
rect 220802 183922 220858 183978
rect 220926 183922 220982 183978
rect 201628 128402 201684 128458
rect 220554 166294 220610 166350
rect 220678 166294 220734 166350
rect 220802 166294 220858 166350
rect 220926 166294 220982 166350
rect 220554 166170 220610 166226
rect 220678 166170 220734 166226
rect 220802 166170 220858 166226
rect 220926 166170 220982 166226
rect 220554 166046 220610 166102
rect 220678 166046 220734 166102
rect 220802 166046 220858 166102
rect 220926 166046 220982 166102
rect 220554 165922 220610 165978
rect 220678 165922 220734 165978
rect 220802 165922 220858 165978
rect 220926 165922 220982 165978
rect 220554 148294 220610 148350
rect 220678 148294 220734 148350
rect 220802 148294 220858 148350
rect 220926 148294 220982 148350
rect 220554 148170 220610 148226
rect 220678 148170 220734 148226
rect 220802 148170 220858 148226
rect 220926 148170 220982 148226
rect 220554 148046 220610 148102
rect 220678 148046 220734 148102
rect 220802 148046 220858 148102
rect 220926 148046 220982 148102
rect 220554 147922 220610 147978
rect 220678 147922 220734 147978
rect 220802 147922 220858 147978
rect 220926 147922 220982 147978
rect 210518 130294 210574 130350
rect 210642 130294 210698 130350
rect 210518 130170 210574 130226
rect 210642 130170 210698 130226
rect 210518 130046 210574 130102
rect 210642 130046 210698 130102
rect 210518 129922 210574 129978
rect 210642 129922 210698 129978
rect 220554 130294 220610 130350
rect 220678 130294 220734 130350
rect 220802 130294 220858 130350
rect 220926 130294 220982 130350
rect 220554 130170 220610 130226
rect 220678 130170 220734 130226
rect 220802 130170 220858 130226
rect 220926 130170 220982 130226
rect 220554 130046 220610 130102
rect 220678 130046 220734 130102
rect 220802 130046 220858 130102
rect 220926 130046 220982 130102
rect 220554 129922 220610 129978
rect 220678 129922 220734 129978
rect 220802 129922 220858 129978
rect 220926 129922 220982 129978
rect 210518 112294 210574 112350
rect 210642 112294 210698 112350
rect 210518 112170 210574 112226
rect 210642 112170 210698 112226
rect 210518 112046 210574 112102
rect 210642 112046 210698 112102
rect 210518 111922 210574 111978
rect 210642 111922 210698 111978
rect 220554 112294 220610 112350
rect 220678 112294 220734 112350
rect 220802 112294 220858 112350
rect 220926 112294 220982 112350
rect 220554 112170 220610 112226
rect 220678 112170 220734 112226
rect 220802 112170 220858 112226
rect 220926 112170 220982 112226
rect 220554 112046 220610 112102
rect 220678 112046 220734 112102
rect 220802 112046 220858 112102
rect 220926 112046 220982 112102
rect 220554 111922 220610 111978
rect 220678 111922 220734 111978
rect 220802 111922 220858 111978
rect 220926 111922 220982 111978
rect 220554 94294 220610 94350
rect 220678 94294 220734 94350
rect 220802 94294 220858 94350
rect 220926 94294 220982 94350
rect 220554 94170 220610 94226
rect 220678 94170 220734 94226
rect 220802 94170 220858 94226
rect 220926 94170 220982 94226
rect 220554 94046 220610 94102
rect 220678 94046 220734 94102
rect 220802 94046 220858 94102
rect 220926 94046 220982 94102
rect 220554 93922 220610 93978
rect 220678 93922 220734 93978
rect 220802 93922 220858 93978
rect 220926 93922 220982 93978
rect 203196 56222 203252 56278
rect 220554 76294 220610 76350
rect 220678 76294 220734 76350
rect 220802 76294 220858 76350
rect 220926 76294 220982 76350
rect 220554 76170 220610 76226
rect 220678 76170 220734 76226
rect 220802 76170 220858 76226
rect 220926 76170 220982 76226
rect 220554 76046 220610 76102
rect 220678 76046 220734 76102
rect 220802 76046 220858 76102
rect 220926 76046 220982 76102
rect 220554 75922 220610 75978
rect 220678 75922 220734 75978
rect 220802 75922 220858 75978
rect 220926 75922 220982 75978
rect 210518 58294 210574 58350
rect 210642 58294 210698 58350
rect 210518 58170 210574 58226
rect 210642 58170 210698 58226
rect 210518 58046 210574 58102
rect 210642 58046 210698 58102
rect 210518 57922 210574 57978
rect 210642 57922 210698 57978
rect 220554 58294 220610 58350
rect 220678 58294 220734 58350
rect 220802 58294 220858 58350
rect 220926 58294 220982 58350
rect 220554 58170 220610 58226
rect 220678 58170 220734 58226
rect 220802 58170 220858 58226
rect 220926 58170 220982 58226
rect 220554 58046 220610 58102
rect 220678 58046 220734 58102
rect 220802 58046 220858 58102
rect 220926 58046 220982 58102
rect 220554 57922 220610 57978
rect 220678 57922 220734 57978
rect 220802 57922 220858 57978
rect 220926 57922 220982 57978
rect 206108 56042 206164 56098
rect 210518 40294 210574 40350
rect 210642 40294 210698 40350
rect 210518 40170 210574 40226
rect 210642 40170 210698 40226
rect 210518 40046 210574 40102
rect 210642 40046 210698 40102
rect 210518 39922 210574 39978
rect 210642 39922 210698 39978
rect 220554 40294 220610 40350
rect 220678 40294 220734 40350
rect 220802 40294 220858 40350
rect 220926 40294 220982 40350
rect 220554 40170 220610 40226
rect 220678 40170 220734 40226
rect 220802 40170 220858 40226
rect 220926 40170 220982 40226
rect 220554 40046 220610 40102
rect 220678 40046 220734 40102
rect 220802 40046 220858 40102
rect 220926 40046 220982 40102
rect 220554 39922 220610 39978
rect 220678 39922 220734 39978
rect 220802 39922 220858 39978
rect 220926 39922 220982 39978
rect 220554 22294 220610 22350
rect 220678 22294 220734 22350
rect 220802 22294 220858 22350
rect 220926 22294 220982 22350
rect 220554 22170 220610 22226
rect 220678 22170 220734 22226
rect 220802 22170 220858 22226
rect 220926 22170 220982 22226
rect 220554 22046 220610 22102
rect 220678 22046 220734 22102
rect 220802 22046 220858 22102
rect 220926 22046 220982 22102
rect 220554 21922 220610 21978
rect 220678 21922 220734 21978
rect 220802 21922 220858 21978
rect 220926 21922 220982 21978
rect 193554 -1176 193610 -1120
rect 193678 -1176 193734 -1120
rect 193802 -1176 193858 -1120
rect 193926 -1176 193982 -1120
rect 193554 -1300 193610 -1244
rect 193678 -1300 193734 -1244
rect 193802 -1300 193858 -1244
rect 193926 -1300 193982 -1244
rect 193554 -1424 193610 -1368
rect 193678 -1424 193734 -1368
rect 193802 -1424 193858 -1368
rect 193926 -1424 193982 -1368
rect 193554 -1548 193610 -1492
rect 193678 -1548 193734 -1492
rect 193802 -1548 193858 -1492
rect 193926 -1548 193982 -1492
rect 220554 4294 220610 4350
rect 220678 4294 220734 4350
rect 220802 4294 220858 4350
rect 220926 4294 220982 4350
rect 220554 4170 220610 4226
rect 220678 4170 220734 4226
rect 220802 4170 220858 4226
rect 220926 4170 220982 4226
rect 220554 4046 220610 4102
rect 220678 4046 220734 4102
rect 220802 4046 220858 4102
rect 220926 4046 220982 4102
rect 220554 3922 220610 3978
rect 220678 3922 220734 3978
rect 220802 3922 220858 3978
rect 220926 3922 220982 3978
rect 220554 -216 220610 -160
rect 220678 -216 220734 -160
rect 220802 -216 220858 -160
rect 220926 -216 220982 -160
rect 220554 -340 220610 -284
rect 220678 -340 220734 -284
rect 220802 -340 220858 -284
rect 220926 -340 220982 -284
rect 220554 -464 220610 -408
rect 220678 -464 220734 -408
rect 220802 -464 220858 -408
rect 220926 -464 220982 -408
rect 220554 -588 220610 -532
rect 220678 -588 220734 -532
rect 220802 -588 220858 -532
rect 220926 -588 220982 -532
rect 224274 424294 224330 424350
rect 224398 424294 224454 424350
rect 224522 424294 224578 424350
rect 224646 424294 224702 424350
rect 224274 424170 224330 424226
rect 224398 424170 224454 424226
rect 224522 424170 224578 424226
rect 224646 424170 224702 424226
rect 224274 424046 224330 424102
rect 224398 424046 224454 424102
rect 224522 424046 224578 424102
rect 224646 424046 224702 424102
rect 224274 423922 224330 423978
rect 224398 423922 224454 423978
rect 224522 423922 224578 423978
rect 224646 423922 224702 423978
rect 287878 550294 287934 550350
rect 288002 550294 288058 550350
rect 287878 550170 287934 550226
rect 288002 550170 288058 550226
rect 287878 550046 287934 550102
rect 288002 550046 288058 550102
rect 287878 549922 287934 549978
rect 288002 549922 288058 549978
rect 318598 550294 318654 550350
rect 318722 550294 318778 550350
rect 318598 550170 318654 550226
rect 318722 550170 318778 550226
rect 318598 550046 318654 550102
rect 318722 550046 318778 550102
rect 318598 549922 318654 549978
rect 318722 549922 318778 549978
rect 263788 533402 263844 533458
rect 254994 460294 255050 460350
rect 255118 460294 255174 460350
rect 255242 460294 255298 460350
rect 255366 460294 255422 460350
rect 254994 460170 255050 460226
rect 255118 460170 255174 460226
rect 255242 460170 255298 460226
rect 255366 460170 255422 460226
rect 254994 460046 255050 460102
rect 255118 460046 255174 460102
rect 255242 460046 255298 460102
rect 255366 460046 255422 460102
rect 254994 459922 255050 459978
rect 255118 459922 255174 459978
rect 255242 459922 255298 459978
rect 255366 459922 255422 459978
rect 251274 436294 251330 436350
rect 251398 436294 251454 436350
rect 251522 436294 251578 436350
rect 251646 436294 251702 436350
rect 251274 436170 251330 436226
rect 251398 436170 251454 436226
rect 251522 436170 251578 436226
rect 251646 436170 251702 436226
rect 251274 436046 251330 436102
rect 251398 436046 251454 436102
rect 251522 436046 251578 436102
rect 251646 436046 251702 436102
rect 251274 435922 251330 435978
rect 251398 435922 251454 435978
rect 251522 435922 251578 435978
rect 251646 435922 251702 435978
rect 241238 418294 241294 418350
rect 241362 418294 241418 418350
rect 241238 418170 241294 418226
rect 241362 418170 241418 418226
rect 241238 418046 241294 418102
rect 241362 418046 241418 418102
rect 241238 417922 241294 417978
rect 241362 417922 241418 417978
rect 254994 442294 255050 442350
rect 255118 442294 255174 442350
rect 255242 442294 255298 442350
rect 255366 442294 255422 442350
rect 254994 442170 255050 442226
rect 255118 442170 255174 442226
rect 255242 442170 255298 442226
rect 255366 442170 255422 442226
rect 254994 442046 255050 442102
rect 255118 442046 255174 442102
rect 255242 442046 255298 442102
rect 255366 442046 255422 442102
rect 254994 441922 255050 441978
rect 255118 441922 255174 441978
rect 255242 441922 255298 441978
rect 255366 441922 255422 441978
rect 251274 418294 251330 418350
rect 251398 418294 251454 418350
rect 251522 418294 251578 418350
rect 251646 418294 251702 418350
rect 251274 418170 251330 418226
rect 251398 418170 251454 418226
rect 251522 418170 251578 418226
rect 251646 418170 251702 418226
rect 251274 418046 251330 418102
rect 251398 418046 251454 418102
rect 251522 418046 251578 418102
rect 251646 418046 251702 418102
rect 251274 417922 251330 417978
rect 251398 417922 251454 417978
rect 251522 417922 251578 417978
rect 251646 417922 251702 417978
rect 249452 409022 249508 409078
rect 224274 406294 224330 406350
rect 224398 406294 224454 406350
rect 224522 406294 224578 406350
rect 224646 406294 224702 406350
rect 224274 406170 224330 406226
rect 224398 406170 224454 406226
rect 224522 406170 224578 406226
rect 224646 406170 224702 406226
rect 224274 406046 224330 406102
rect 224398 406046 224454 406102
rect 224522 406046 224578 406102
rect 224646 406046 224702 406102
rect 224274 405922 224330 405978
rect 224398 405922 224454 405978
rect 224522 405922 224578 405978
rect 224646 405922 224702 405978
rect 225878 406294 225934 406350
rect 226002 406294 226058 406350
rect 225878 406170 225934 406226
rect 226002 406170 226058 406226
rect 225878 406046 225934 406102
rect 226002 406046 226058 406102
rect 225878 405922 225934 405978
rect 226002 405922 226058 405978
rect 241238 400294 241294 400350
rect 241362 400294 241418 400350
rect 241238 400170 241294 400226
rect 241362 400170 241418 400226
rect 241238 400046 241294 400102
rect 241362 400046 241418 400102
rect 241238 399922 241294 399978
rect 241362 399922 241418 399978
rect 254994 424294 255050 424350
rect 255118 424294 255174 424350
rect 255242 424294 255298 424350
rect 255366 424294 255422 424350
rect 254994 424170 255050 424226
rect 255118 424170 255174 424226
rect 255242 424170 255298 424226
rect 255366 424170 255422 424226
rect 254994 424046 255050 424102
rect 255118 424046 255174 424102
rect 255242 424046 255298 424102
rect 255366 424046 255422 424102
rect 254994 423922 255050 423978
rect 255118 423922 255174 423978
rect 255242 423922 255298 423978
rect 255366 423922 255422 423978
rect 252812 409922 252868 409978
rect 272518 544294 272574 544350
rect 272642 544294 272698 544350
rect 272518 544170 272574 544226
rect 272642 544170 272698 544226
rect 272518 544046 272574 544102
rect 272642 544046 272698 544102
rect 272518 543922 272574 543978
rect 272642 543922 272698 543978
rect 303238 544294 303294 544350
rect 303362 544294 303418 544350
rect 303238 544170 303294 544226
rect 303362 544170 303418 544226
rect 303238 544046 303294 544102
rect 303362 544046 303418 544102
rect 303238 543922 303294 543978
rect 303362 543922 303418 543978
rect 287878 532294 287934 532350
rect 288002 532294 288058 532350
rect 287878 532170 287934 532226
rect 288002 532170 288058 532226
rect 287878 532046 287934 532102
rect 288002 532046 288058 532102
rect 287878 531922 287934 531978
rect 288002 531922 288058 531978
rect 318598 532294 318654 532350
rect 318722 532294 318778 532350
rect 318598 532170 318654 532226
rect 318722 532170 318778 532226
rect 318598 532046 318654 532102
rect 318722 532046 318778 532102
rect 318598 531922 318654 531978
rect 318722 531922 318778 531978
rect 272518 526294 272574 526350
rect 272642 526294 272698 526350
rect 272518 526170 272574 526226
rect 272642 526170 272698 526226
rect 272518 526046 272574 526102
rect 272642 526046 272698 526102
rect 272518 525922 272574 525978
rect 272642 525922 272698 525978
rect 303238 526294 303294 526350
rect 303362 526294 303418 526350
rect 303238 526170 303294 526226
rect 303362 526170 303418 526226
rect 303238 526046 303294 526102
rect 303362 526046 303418 526102
rect 303238 525922 303294 525978
rect 303362 525922 303418 525978
rect 287878 514294 287934 514350
rect 288002 514294 288058 514350
rect 287878 514170 287934 514226
rect 288002 514170 288058 514226
rect 287878 514046 287934 514102
rect 288002 514046 288058 514102
rect 287878 513922 287934 513978
rect 288002 513922 288058 513978
rect 318598 514294 318654 514350
rect 318722 514294 318778 514350
rect 318598 514170 318654 514226
rect 318722 514170 318778 514226
rect 318598 514046 318654 514102
rect 318722 514046 318778 514102
rect 318598 513922 318654 513978
rect 318722 513922 318778 513978
rect 272518 508294 272574 508350
rect 272642 508294 272698 508350
rect 272518 508170 272574 508226
rect 272642 508170 272698 508226
rect 272518 508046 272574 508102
rect 272642 508046 272698 508102
rect 272518 507922 272574 507978
rect 272642 507922 272698 507978
rect 303238 508294 303294 508350
rect 303362 508294 303418 508350
rect 303238 508170 303294 508226
rect 303362 508170 303418 508226
rect 303238 508046 303294 508102
rect 303362 508046 303418 508102
rect 303238 507922 303294 507978
rect 303362 507922 303418 507978
rect 287878 496294 287934 496350
rect 288002 496294 288058 496350
rect 287878 496170 287934 496226
rect 288002 496170 288058 496226
rect 287878 496046 287934 496102
rect 288002 496046 288058 496102
rect 287878 495922 287934 495978
rect 288002 495922 288058 495978
rect 318598 496294 318654 496350
rect 318722 496294 318778 496350
rect 318598 496170 318654 496226
rect 318722 496170 318778 496226
rect 318598 496046 318654 496102
rect 318722 496046 318778 496102
rect 318598 495922 318654 495978
rect 318722 495922 318778 495978
rect 272518 490294 272574 490350
rect 272642 490294 272698 490350
rect 272518 490170 272574 490226
rect 272642 490170 272698 490226
rect 272518 490046 272574 490102
rect 272642 490046 272698 490102
rect 272518 489922 272574 489978
rect 272642 489922 272698 489978
rect 303238 490294 303294 490350
rect 303362 490294 303418 490350
rect 303238 490170 303294 490226
rect 303362 490170 303418 490226
rect 303238 490046 303294 490102
rect 303362 490046 303418 490102
rect 303238 489922 303294 489978
rect 303362 489922 303418 489978
rect 287878 478294 287934 478350
rect 288002 478294 288058 478350
rect 287878 478170 287934 478226
rect 288002 478170 288058 478226
rect 287878 478046 287934 478102
rect 288002 478046 288058 478102
rect 287878 477922 287934 477978
rect 288002 477922 288058 477978
rect 318598 478294 318654 478350
rect 318722 478294 318778 478350
rect 318598 478170 318654 478226
rect 318722 478170 318778 478226
rect 318598 478046 318654 478102
rect 318722 478046 318778 478102
rect 318598 477922 318654 477978
rect 318722 477922 318778 477978
rect 263788 473642 263844 473698
rect 264124 469502 264180 469558
rect 264012 467882 264068 467938
rect 263788 465182 263844 465238
rect 263788 463562 263844 463618
rect 264684 474542 264740 474598
rect 272518 472294 272574 472350
rect 272642 472294 272698 472350
rect 272518 472170 272574 472226
rect 272642 472170 272698 472226
rect 272518 472046 272574 472102
rect 272642 472046 272698 472102
rect 272518 471922 272574 471978
rect 272642 471922 272698 471978
rect 303238 472294 303294 472350
rect 303362 472294 303418 472350
rect 303238 472170 303294 472226
rect 303362 472170 303418 472226
rect 303238 472046 303294 472102
rect 303362 472046 303418 472102
rect 303238 471922 303294 471978
rect 303362 471922 303418 471978
rect 287878 460294 287934 460350
rect 288002 460294 288058 460350
rect 287878 460170 287934 460226
rect 288002 460170 288058 460226
rect 287878 460046 287934 460102
rect 288002 460046 288058 460102
rect 287878 459922 287934 459978
rect 288002 459922 288058 459978
rect 318598 460294 318654 460350
rect 318722 460294 318778 460350
rect 318598 460170 318654 460226
rect 318722 460170 318778 460226
rect 318598 460046 318654 460102
rect 318722 460046 318778 460102
rect 318598 459922 318654 459978
rect 318722 459922 318778 459978
rect 272518 454294 272574 454350
rect 272642 454294 272698 454350
rect 272518 454170 272574 454226
rect 272642 454170 272698 454226
rect 272518 454046 272574 454102
rect 272642 454046 272698 454102
rect 272518 453922 272574 453978
rect 272642 453922 272698 453978
rect 303238 454294 303294 454350
rect 303362 454294 303418 454350
rect 303238 454170 303294 454226
rect 303362 454170 303418 454226
rect 303238 454046 303294 454102
rect 303362 454046 303418 454102
rect 303238 453922 303294 453978
rect 303362 453922 303418 453978
rect 287878 442294 287934 442350
rect 288002 442294 288058 442350
rect 287878 442170 287934 442226
rect 288002 442170 288058 442226
rect 287878 442046 287934 442102
rect 288002 442046 288058 442102
rect 287878 441922 287934 441978
rect 288002 441922 288058 441978
rect 318598 442294 318654 442350
rect 318722 442294 318778 442350
rect 318598 442170 318654 442226
rect 318722 442170 318778 442226
rect 318598 442046 318654 442102
rect 318722 442046 318778 442102
rect 318598 441922 318654 441978
rect 318722 441922 318778 441978
rect 272518 436294 272574 436350
rect 272642 436294 272698 436350
rect 272518 436170 272574 436226
rect 272642 436170 272698 436226
rect 272518 436046 272574 436102
rect 272642 436046 272698 436102
rect 272518 435922 272574 435978
rect 272642 435922 272698 435978
rect 303238 436294 303294 436350
rect 303362 436294 303418 436350
rect 303238 436170 303294 436226
rect 303362 436170 303418 436226
rect 303238 436046 303294 436102
rect 303362 436046 303418 436102
rect 303238 435922 303294 435978
rect 303362 435922 303418 435978
rect 287878 424294 287934 424350
rect 288002 424294 288058 424350
rect 287878 424170 287934 424226
rect 288002 424170 288058 424226
rect 287878 424046 287934 424102
rect 288002 424046 288058 424102
rect 287878 423922 287934 423978
rect 288002 423922 288058 423978
rect 318598 424294 318654 424350
rect 318722 424294 318778 424350
rect 318598 424170 318654 424226
rect 318722 424170 318778 424226
rect 318598 424046 318654 424102
rect 318722 424046 318778 424102
rect 318598 423922 318654 423978
rect 318722 423922 318778 423978
rect 272518 418294 272574 418350
rect 272642 418294 272698 418350
rect 272518 418170 272574 418226
rect 272642 418170 272698 418226
rect 272518 418046 272574 418102
rect 272642 418046 272698 418102
rect 272518 417922 272574 417978
rect 272642 417922 272698 417978
rect 303238 418294 303294 418350
rect 303362 418294 303418 418350
rect 303238 418170 303294 418226
rect 303362 418170 303418 418226
rect 303238 418046 303294 418102
rect 303362 418046 303418 418102
rect 303238 417922 303294 417978
rect 303362 417922 303418 417978
rect 260316 414962 260372 415018
rect 254994 406294 255050 406350
rect 255118 406294 255174 406350
rect 255242 406294 255298 406350
rect 255366 406294 255422 406350
rect 254994 406170 255050 406226
rect 255118 406170 255174 406226
rect 255242 406170 255298 406226
rect 255366 406170 255422 406226
rect 251274 400294 251330 400350
rect 251398 400294 251454 400350
rect 251522 400294 251578 400350
rect 251646 400294 251702 400350
rect 251274 400170 251330 400226
rect 251398 400170 251454 400226
rect 251522 400170 251578 400226
rect 251646 400170 251702 400226
rect 251274 400046 251330 400102
rect 251398 400046 251454 400102
rect 251522 400046 251578 400102
rect 251646 400046 251702 400102
rect 251274 399922 251330 399978
rect 251398 399922 251454 399978
rect 251522 399922 251578 399978
rect 251646 399922 251702 399978
rect 224274 388294 224330 388350
rect 224398 388294 224454 388350
rect 224522 388294 224578 388350
rect 224646 388294 224702 388350
rect 225836 388333 225892 388389
rect 225940 388333 225996 388389
rect 226044 388333 226100 388389
rect 224274 388170 224330 388226
rect 224398 388170 224454 388226
rect 224522 388170 224578 388226
rect 224646 388170 224702 388226
rect 224274 388046 224330 388102
rect 224398 388046 224454 388102
rect 224522 388046 224578 388102
rect 224646 388046 224702 388102
rect 224274 387922 224330 387978
rect 224398 387922 224454 387978
rect 224522 387922 224578 387978
rect 224646 387922 224702 387978
rect 224274 370294 224330 370350
rect 224398 370294 224454 370350
rect 224522 370294 224578 370350
rect 224646 370294 224702 370350
rect 224274 370170 224330 370226
rect 224398 370170 224454 370226
rect 224522 370170 224578 370226
rect 224646 370170 224702 370226
rect 224274 370046 224330 370102
rect 224398 370046 224454 370102
rect 224522 370046 224578 370102
rect 224646 370046 224702 370102
rect 224274 369922 224330 369978
rect 224398 369922 224454 369978
rect 224522 369922 224578 369978
rect 224646 369922 224702 369978
rect 254994 406046 255050 406102
rect 255118 406046 255174 406102
rect 255242 406046 255298 406102
rect 255366 406046 255422 406102
rect 254994 405922 255050 405978
rect 255118 405922 255174 405978
rect 255242 405922 255298 405978
rect 255366 405922 255422 405978
rect 251274 382294 251330 382350
rect 251398 382294 251454 382350
rect 251522 382294 251578 382350
rect 251646 382294 251702 382350
rect 251274 382170 251330 382226
rect 251398 382170 251454 382226
rect 251522 382170 251578 382226
rect 251646 382170 251702 382226
rect 251274 382046 251330 382102
rect 251398 382046 251454 382102
rect 251522 382046 251578 382102
rect 251646 382046 251702 382102
rect 251274 381922 251330 381978
rect 251398 381922 251454 381978
rect 251522 381922 251578 381978
rect 251646 381922 251702 381978
rect 251274 364294 251330 364350
rect 251398 364294 251454 364350
rect 251522 364294 251578 364350
rect 251646 364294 251702 364350
rect 251274 364170 251330 364226
rect 251398 364170 251454 364226
rect 251522 364170 251578 364226
rect 251646 364170 251702 364226
rect 251274 364046 251330 364102
rect 251398 364046 251454 364102
rect 251522 364046 251578 364102
rect 251646 364046 251702 364102
rect 251274 363922 251330 363978
rect 251398 363922 251454 363978
rect 251522 363922 251578 363978
rect 251646 363922 251702 363978
rect 224274 352294 224330 352350
rect 224398 352294 224454 352350
rect 224522 352294 224578 352350
rect 224646 352294 224702 352350
rect 224274 352170 224330 352226
rect 224398 352170 224454 352226
rect 224522 352170 224578 352226
rect 224646 352170 224702 352226
rect 224274 352046 224330 352102
rect 224398 352046 224454 352102
rect 224522 352046 224578 352102
rect 224646 352046 224702 352102
rect 224274 351922 224330 351978
rect 224398 351922 224454 351978
rect 224522 351922 224578 351978
rect 224646 351922 224702 351978
rect 225878 352294 225934 352350
rect 226002 352294 226058 352350
rect 225878 352170 225934 352226
rect 226002 352170 226058 352226
rect 225878 352046 225934 352102
rect 226002 352046 226058 352102
rect 225878 351922 225934 351978
rect 226002 351922 226058 351978
rect 241238 346294 241294 346350
rect 241362 346294 241418 346350
rect 241238 346170 241294 346226
rect 241362 346170 241418 346226
rect 241238 346046 241294 346102
rect 241362 346046 241418 346102
rect 241238 345922 241294 345978
rect 241362 345922 241418 345978
rect 251274 346294 251330 346350
rect 251398 346294 251454 346350
rect 251522 346294 251578 346350
rect 251646 346294 251702 346350
rect 251274 346170 251330 346226
rect 251398 346170 251454 346226
rect 251522 346170 251578 346226
rect 251646 346170 251702 346226
rect 251274 346046 251330 346102
rect 251398 346046 251454 346102
rect 251522 346046 251578 346102
rect 251646 346046 251702 346102
rect 251274 345922 251330 345978
rect 251398 345922 251454 345978
rect 251522 345922 251578 345978
rect 251646 345922 251702 345978
rect 224274 334294 224330 334350
rect 224398 334294 224454 334350
rect 224522 334294 224578 334350
rect 224646 334294 224702 334350
rect 224274 334170 224330 334226
rect 224398 334170 224454 334226
rect 224522 334170 224578 334226
rect 224646 334170 224702 334226
rect 224274 334046 224330 334102
rect 224398 334046 224454 334102
rect 224522 334046 224578 334102
rect 224646 334046 224702 334102
rect 224274 333922 224330 333978
rect 224398 333922 224454 333978
rect 224522 333922 224578 333978
rect 224646 333922 224702 333978
rect 225878 334294 225934 334350
rect 226002 334294 226058 334350
rect 225878 334170 225934 334226
rect 226002 334170 226058 334226
rect 225878 334046 225934 334102
rect 226002 334046 226058 334102
rect 225878 333922 225934 333978
rect 226002 333922 226058 333978
rect 241238 328294 241294 328350
rect 241362 328294 241418 328350
rect 241238 328170 241294 328226
rect 241362 328170 241418 328226
rect 241238 328046 241294 328102
rect 241362 328046 241418 328102
rect 241238 327922 241294 327978
rect 241362 327922 241418 327978
rect 254994 388294 255050 388350
rect 255118 388294 255174 388350
rect 255242 388294 255298 388350
rect 255366 388294 255422 388350
rect 254994 388170 255050 388226
rect 255118 388170 255174 388226
rect 255242 388170 255298 388226
rect 255366 388170 255422 388226
rect 254994 388046 255050 388102
rect 255118 388046 255174 388102
rect 255242 388046 255298 388102
rect 255366 388046 255422 388102
rect 254994 387922 255050 387978
rect 255118 387922 255174 387978
rect 255242 387922 255298 387978
rect 255366 387922 255422 387978
rect 262220 406682 262276 406738
rect 262108 404702 262164 404758
rect 260316 404522 260372 404578
rect 263788 411722 263844 411778
rect 263452 408302 263508 408358
rect 263788 406862 263844 406918
rect 263900 407042 263956 407098
rect 287878 406294 287934 406350
rect 288002 406294 288058 406350
rect 287878 406170 287934 406226
rect 288002 406170 288058 406226
rect 287878 406046 287934 406102
rect 288002 406046 288058 406102
rect 287878 405922 287934 405978
rect 288002 405922 288058 405978
rect 318598 406294 318654 406350
rect 318722 406294 318778 406350
rect 318598 406170 318654 406226
rect 318722 406170 318778 406226
rect 318598 406046 318654 406102
rect 318722 406046 318778 406102
rect 318598 405922 318654 405978
rect 318722 405922 318778 405978
rect 263788 403982 263844 404038
rect 263788 403082 263844 403138
rect 263900 402902 263956 402958
rect 272518 400294 272574 400350
rect 272642 400294 272698 400350
rect 272518 400170 272574 400226
rect 272642 400170 272698 400226
rect 272518 400046 272574 400102
rect 272642 400046 272698 400102
rect 272518 399922 272574 399978
rect 272642 399922 272698 399978
rect 303238 400294 303294 400350
rect 303362 400294 303418 400350
rect 303238 400170 303294 400226
rect 303362 400170 303418 400226
rect 303238 400046 303294 400102
rect 303362 400046 303418 400102
rect 303238 399922 303294 399978
rect 303362 399922 303418 399978
rect 262108 399482 262164 399538
rect 263788 399662 263844 399718
rect 263788 398042 263844 398098
rect 263788 396422 263844 396478
rect 263900 396242 263956 396298
rect 263788 393002 263844 393058
rect 263788 391382 263844 391438
rect 287878 388294 287934 388350
rect 288002 388294 288058 388350
rect 287878 388170 287934 388226
rect 288002 388170 288058 388226
rect 287878 388046 287934 388102
rect 288002 388046 288058 388102
rect 287878 387922 287934 387978
rect 288002 387922 288058 387978
rect 318598 388294 318654 388350
rect 318722 388294 318778 388350
rect 318598 388170 318654 388226
rect 318722 388170 318778 388226
rect 318598 388046 318654 388102
rect 318722 388046 318778 388102
rect 318598 387922 318654 387978
rect 318722 387922 318778 387978
rect 272518 382294 272574 382350
rect 272642 382294 272698 382350
rect 272518 382170 272574 382226
rect 272642 382170 272698 382226
rect 272518 382046 272574 382102
rect 272642 382046 272698 382102
rect 272518 381922 272574 381978
rect 272642 381922 272698 381978
rect 303238 382294 303294 382350
rect 303362 382294 303418 382350
rect 303238 382170 303294 382226
rect 303362 382170 303418 382226
rect 303238 382046 303294 382102
rect 303362 382046 303418 382102
rect 303238 381922 303294 381978
rect 303362 381922 303418 381978
rect 254994 370294 255050 370350
rect 255118 370294 255174 370350
rect 255242 370294 255298 370350
rect 255366 370294 255422 370350
rect 254994 370170 255050 370226
rect 255118 370170 255174 370226
rect 255242 370170 255298 370226
rect 255366 370170 255422 370226
rect 254994 370046 255050 370102
rect 255118 370046 255174 370102
rect 255242 370046 255298 370102
rect 255366 370046 255422 370102
rect 254994 369922 255050 369978
rect 255118 369922 255174 369978
rect 255242 369922 255298 369978
rect 255366 369922 255422 369978
rect 287878 370294 287934 370350
rect 288002 370294 288058 370350
rect 287878 370170 287934 370226
rect 288002 370170 288058 370226
rect 287878 370046 287934 370102
rect 288002 370046 288058 370102
rect 287878 369922 287934 369978
rect 288002 369922 288058 369978
rect 318598 370294 318654 370350
rect 318722 370294 318778 370350
rect 318598 370170 318654 370226
rect 318722 370170 318778 370226
rect 318598 370046 318654 370102
rect 318722 370046 318778 370102
rect 318598 369922 318654 369978
rect 318722 369922 318778 369978
rect 272518 364294 272574 364350
rect 272642 364294 272698 364350
rect 272518 364170 272574 364226
rect 272642 364170 272698 364226
rect 272518 364046 272574 364102
rect 272642 364046 272698 364102
rect 272518 363922 272574 363978
rect 272642 363922 272698 363978
rect 303238 364294 303294 364350
rect 303362 364294 303418 364350
rect 303238 364170 303294 364226
rect 303362 364170 303418 364226
rect 303238 364046 303294 364102
rect 303362 364046 303418 364102
rect 303238 363922 303294 363978
rect 303362 363922 303418 363978
rect 254994 352294 255050 352350
rect 255118 352294 255174 352350
rect 255242 352294 255298 352350
rect 255366 352294 255422 352350
rect 254994 352170 255050 352226
rect 255118 352170 255174 352226
rect 255242 352170 255298 352226
rect 255366 352170 255422 352226
rect 254994 352046 255050 352102
rect 255118 352046 255174 352102
rect 255242 352046 255298 352102
rect 255366 352046 255422 352102
rect 254994 351922 255050 351978
rect 255118 351922 255174 351978
rect 255242 351922 255298 351978
rect 255366 351922 255422 351978
rect 263788 349442 263844 349498
rect 263340 348542 263396 348598
rect 263788 347822 263844 347878
rect 263788 344582 263844 344638
rect 263900 344402 263956 344458
rect 262108 343502 262164 343558
rect 263788 342962 263844 343018
rect 263788 341702 263844 341758
rect 263900 341522 263956 341578
rect 263788 341342 263844 341398
rect 263788 340442 263844 340498
rect 260092 338462 260148 338518
rect 260316 340262 260372 340318
rect 264684 342782 264740 342838
rect 254994 334294 255050 334350
rect 255118 334294 255174 334350
rect 255242 334294 255298 334350
rect 255366 334294 255422 334350
rect 254994 334170 255050 334226
rect 255118 334170 255174 334226
rect 255242 334170 255298 334226
rect 255366 334170 255422 334226
rect 254994 334046 255050 334102
rect 255118 334046 255174 334102
rect 255242 334046 255298 334102
rect 255366 334046 255422 334102
rect 254994 333922 255050 333978
rect 255118 333922 255174 333978
rect 255242 333922 255298 333978
rect 255366 333922 255422 333978
rect 251274 328294 251330 328350
rect 251398 328294 251454 328350
rect 251522 328294 251578 328350
rect 251646 328294 251702 328350
rect 251274 328170 251330 328226
rect 251398 328170 251454 328226
rect 251522 328170 251578 328226
rect 251646 328170 251702 328226
rect 251274 328046 251330 328102
rect 251398 328046 251454 328102
rect 251522 328046 251578 328102
rect 251646 328046 251702 328102
rect 251274 327922 251330 327978
rect 251398 327922 251454 327978
rect 251522 327922 251578 327978
rect 251646 327922 251702 327978
rect 224274 316294 224330 316350
rect 224398 316294 224454 316350
rect 224522 316294 224578 316350
rect 224646 316294 224702 316350
rect 224274 316170 224330 316226
rect 224398 316170 224454 316226
rect 224522 316170 224578 316226
rect 224646 316170 224702 316226
rect 224274 316046 224330 316102
rect 224398 316046 224454 316102
rect 224522 316046 224578 316102
rect 224646 316046 224702 316102
rect 224274 315922 224330 315978
rect 224398 315922 224454 315978
rect 224522 315922 224578 315978
rect 224646 315922 224702 315978
rect 224274 298294 224330 298350
rect 224398 298294 224454 298350
rect 224522 298294 224578 298350
rect 224646 298294 224702 298350
rect 224274 298170 224330 298226
rect 224398 298170 224454 298226
rect 224522 298170 224578 298226
rect 224646 298170 224702 298226
rect 224274 298046 224330 298102
rect 224398 298046 224454 298102
rect 224522 298046 224578 298102
rect 224646 298046 224702 298102
rect 224274 297922 224330 297978
rect 224398 297922 224454 297978
rect 224522 297922 224578 297978
rect 224646 297922 224702 297978
rect 251274 310294 251330 310350
rect 251398 310294 251454 310350
rect 251522 310294 251578 310350
rect 251646 310294 251702 310350
rect 251274 310170 251330 310226
rect 251398 310170 251454 310226
rect 251522 310170 251578 310226
rect 251646 310170 251702 310226
rect 251274 310046 251330 310102
rect 251398 310046 251454 310102
rect 251522 310046 251578 310102
rect 251646 310046 251702 310102
rect 251274 309922 251330 309978
rect 251398 309922 251454 309978
rect 251522 309922 251578 309978
rect 251646 309922 251702 309978
rect 263788 331442 263844 331498
rect 263900 331082 263956 331138
rect 263788 330902 263844 330958
rect 264012 330722 264068 330778
rect 263788 330596 263844 330598
rect 263788 330542 263844 330596
rect 263788 327482 263844 327538
rect 263900 327302 263956 327358
rect 287878 352294 287934 352350
rect 288002 352294 288058 352350
rect 287878 352170 287934 352226
rect 288002 352170 288058 352226
rect 287878 352046 287934 352102
rect 288002 352046 288058 352102
rect 287878 351922 287934 351978
rect 288002 351922 288058 351978
rect 318598 352294 318654 352350
rect 318722 352294 318778 352350
rect 318598 352170 318654 352226
rect 318722 352170 318778 352226
rect 318598 352046 318654 352102
rect 318722 352046 318778 352102
rect 318598 351922 318654 351978
rect 318722 351922 318778 351978
rect 272518 346294 272574 346350
rect 272642 346294 272698 346350
rect 272518 346170 272574 346226
rect 272642 346170 272698 346226
rect 272518 346046 272574 346102
rect 272642 346046 272698 346102
rect 272518 345922 272574 345978
rect 272642 345922 272698 345978
rect 303238 346294 303294 346350
rect 303362 346294 303418 346350
rect 303238 346170 303294 346226
rect 303362 346170 303418 346226
rect 303238 346046 303294 346102
rect 303362 346046 303418 346102
rect 303238 345922 303294 345978
rect 303362 345922 303418 345978
rect 287878 334294 287934 334350
rect 288002 334294 288058 334350
rect 287878 334170 287934 334226
rect 288002 334170 288058 334226
rect 287878 334046 287934 334102
rect 288002 334046 288058 334102
rect 287878 333922 287934 333978
rect 288002 333922 288058 333978
rect 318598 334294 318654 334350
rect 318722 334294 318778 334350
rect 318598 334170 318654 334226
rect 318722 334170 318778 334226
rect 318598 334046 318654 334102
rect 318722 334046 318778 334102
rect 318598 333922 318654 333978
rect 318722 333922 318778 333978
rect 272518 328294 272574 328350
rect 272642 328294 272698 328350
rect 272518 328170 272574 328226
rect 272642 328170 272698 328226
rect 272518 328046 272574 328102
rect 272642 328046 272698 328102
rect 272518 327922 272574 327978
rect 272642 327922 272698 327978
rect 303238 328294 303294 328350
rect 303362 328294 303418 328350
rect 303238 328170 303294 328226
rect 303362 328170 303418 328226
rect 303238 328046 303294 328102
rect 303362 328046 303418 328102
rect 303238 327922 303294 327978
rect 303362 327922 303418 327978
rect 264908 325862 264964 325918
rect 264572 325682 264628 325738
rect 263788 325556 263844 325558
rect 263788 325502 263844 325556
rect 263788 324062 263844 324118
rect 254994 316294 255050 316350
rect 255118 316294 255174 316350
rect 255242 316294 255298 316350
rect 255366 316294 255422 316350
rect 254994 316170 255050 316226
rect 255118 316170 255174 316226
rect 255242 316170 255298 316226
rect 255366 316170 255422 316226
rect 254994 316046 255050 316102
rect 255118 316046 255174 316102
rect 255242 316046 255298 316102
rect 255366 316046 255422 316102
rect 254994 315922 255050 315978
rect 255118 315922 255174 315978
rect 255242 315922 255298 315978
rect 255366 315922 255422 315978
rect 287878 316294 287934 316350
rect 288002 316294 288058 316350
rect 287878 316170 287934 316226
rect 288002 316170 288058 316226
rect 287878 316046 287934 316102
rect 288002 316046 288058 316102
rect 287878 315922 287934 315978
rect 288002 315922 288058 315978
rect 318598 316294 318654 316350
rect 318722 316294 318778 316350
rect 318598 316170 318654 316226
rect 318722 316170 318778 316226
rect 318598 316046 318654 316102
rect 318722 316046 318778 316102
rect 318598 315922 318654 315978
rect 318722 315922 318778 315978
rect 272518 310294 272574 310350
rect 272642 310294 272698 310350
rect 272518 310170 272574 310226
rect 272642 310170 272698 310226
rect 272518 310046 272574 310102
rect 272642 310046 272698 310102
rect 272518 309922 272574 309978
rect 272642 309922 272698 309978
rect 303238 310294 303294 310350
rect 303362 310294 303418 310350
rect 303238 310170 303294 310226
rect 303362 310170 303418 310226
rect 303238 310046 303294 310102
rect 303362 310046 303418 310102
rect 303238 309922 303294 309978
rect 303362 309922 303418 309978
rect 254994 298294 255050 298350
rect 255118 298294 255174 298350
rect 255242 298294 255298 298350
rect 255366 298294 255422 298350
rect 254994 298170 255050 298226
rect 255118 298170 255174 298226
rect 255242 298170 255298 298226
rect 255366 298170 255422 298226
rect 254994 298046 255050 298102
rect 255118 298046 255174 298102
rect 255242 298046 255298 298102
rect 255366 298046 255422 298102
rect 254994 297922 255050 297978
rect 255118 297922 255174 297978
rect 255242 297922 255298 297978
rect 255366 297922 255422 297978
rect 251274 292294 251330 292350
rect 251398 292294 251454 292350
rect 251522 292294 251578 292350
rect 251646 292294 251702 292350
rect 251274 292170 251330 292226
rect 251398 292170 251454 292226
rect 251522 292170 251578 292226
rect 251646 292170 251702 292226
rect 251274 292046 251330 292102
rect 251398 292046 251454 292102
rect 251522 292046 251578 292102
rect 251646 292046 251702 292102
rect 251274 291922 251330 291978
rect 251398 291922 251454 291978
rect 251522 291922 251578 291978
rect 251646 291922 251702 291978
rect 224274 280294 224330 280350
rect 224398 280294 224454 280350
rect 224522 280294 224578 280350
rect 224646 280294 224702 280350
rect 224274 280170 224330 280226
rect 224398 280170 224454 280226
rect 224522 280170 224578 280226
rect 224646 280170 224702 280226
rect 224274 280046 224330 280102
rect 224398 280046 224454 280102
rect 224522 280046 224578 280102
rect 224646 280046 224702 280102
rect 224274 279922 224330 279978
rect 224398 279922 224454 279978
rect 224522 279922 224578 279978
rect 224646 279922 224702 279978
rect 225878 280294 225934 280350
rect 226002 280294 226058 280350
rect 225878 280170 225934 280226
rect 226002 280170 226058 280226
rect 225878 280046 225934 280102
rect 226002 280046 226058 280102
rect 225878 279922 225934 279978
rect 226002 279922 226058 279978
rect 241238 274294 241294 274350
rect 241362 274294 241418 274350
rect 241238 274170 241294 274226
rect 241362 274170 241418 274226
rect 241238 274046 241294 274102
rect 241362 274046 241418 274102
rect 241238 273922 241294 273978
rect 241362 273922 241418 273978
rect 249452 268622 249508 268678
rect 251274 274294 251330 274350
rect 251398 274294 251454 274350
rect 251522 274294 251578 274350
rect 251646 274294 251702 274350
rect 251274 274170 251330 274226
rect 251398 274170 251454 274226
rect 251522 274170 251578 274226
rect 251646 274170 251702 274226
rect 251274 274046 251330 274102
rect 251398 274046 251454 274102
rect 251522 274046 251578 274102
rect 251646 274046 251702 274102
rect 251274 273922 251330 273978
rect 251398 273922 251454 273978
rect 251522 273922 251578 273978
rect 251646 273922 251702 273978
rect 224274 262294 224330 262350
rect 224398 262294 224454 262350
rect 224522 262294 224578 262350
rect 224646 262294 224702 262350
rect 224274 262170 224330 262226
rect 224398 262170 224454 262226
rect 224522 262170 224578 262226
rect 224646 262170 224702 262226
rect 224274 262046 224330 262102
rect 224398 262046 224454 262102
rect 224522 262046 224578 262102
rect 224646 262046 224702 262102
rect 224274 261922 224330 261978
rect 224398 261922 224454 261978
rect 224522 261922 224578 261978
rect 224646 261922 224702 261978
rect 225878 262294 225934 262350
rect 226002 262294 226058 262350
rect 225878 262170 225934 262226
rect 226002 262170 226058 262226
rect 225878 262046 225934 262102
rect 226002 262046 226058 262102
rect 225878 261922 225934 261978
rect 226002 261922 226058 261978
rect 241238 256294 241294 256350
rect 241362 256294 241418 256350
rect 241238 256170 241294 256226
rect 241362 256170 241418 256226
rect 241238 256046 241294 256102
rect 241362 256046 241418 256102
rect 241238 255922 241294 255978
rect 241362 255922 241418 255978
rect 254994 280294 255050 280350
rect 255118 280294 255174 280350
rect 255242 280294 255298 280350
rect 255366 280294 255422 280350
rect 254994 280170 255050 280226
rect 255118 280170 255174 280226
rect 255242 280170 255298 280226
rect 255366 280170 255422 280226
rect 254994 280046 255050 280102
rect 255118 280046 255174 280102
rect 255242 280046 255298 280102
rect 255366 280046 255422 280102
rect 254994 279922 255050 279978
rect 255118 279922 255174 279978
rect 255242 279922 255298 279978
rect 255366 279922 255422 279978
rect 287878 298294 287934 298350
rect 288002 298294 288058 298350
rect 287878 298170 287934 298226
rect 288002 298170 288058 298226
rect 287878 298046 287934 298102
rect 288002 298046 288058 298102
rect 287878 297922 287934 297978
rect 288002 297922 288058 297978
rect 318598 298294 318654 298350
rect 318722 298294 318778 298350
rect 318598 298170 318654 298226
rect 318722 298170 318778 298226
rect 318598 298046 318654 298102
rect 318722 298046 318778 298102
rect 318598 297922 318654 297978
rect 318722 297922 318778 297978
rect 272518 292294 272574 292350
rect 272642 292294 272698 292350
rect 272518 292170 272574 292226
rect 272642 292170 272698 292226
rect 272518 292046 272574 292102
rect 272642 292046 272698 292102
rect 272518 291922 272574 291978
rect 272642 291922 272698 291978
rect 303238 292294 303294 292350
rect 303362 292294 303418 292350
rect 303238 292170 303294 292226
rect 303362 292170 303418 292226
rect 303238 292046 303294 292102
rect 303362 292046 303418 292102
rect 303238 291922 303294 291978
rect 303362 291922 303418 291978
rect 287878 280294 287934 280350
rect 288002 280294 288058 280350
rect 287878 280170 287934 280226
rect 288002 280170 288058 280226
rect 287878 280046 287934 280102
rect 288002 280046 288058 280102
rect 287878 279922 287934 279978
rect 288002 279922 288058 279978
rect 318598 280294 318654 280350
rect 318722 280294 318778 280350
rect 318598 280170 318654 280226
rect 318722 280170 318778 280226
rect 318598 280046 318654 280102
rect 318722 280046 318778 280102
rect 318598 279922 318654 279978
rect 318722 279922 318778 279978
rect 263788 278162 263844 278218
rect 263340 277982 263396 278038
rect 262108 276362 262164 276418
rect 263788 275642 263844 275698
rect 272518 274294 272574 274350
rect 272642 274294 272698 274350
rect 272518 274170 272574 274226
rect 272642 274170 272698 274226
rect 272518 274046 272574 274102
rect 272642 274046 272698 274102
rect 272518 273922 272574 273978
rect 272642 273922 272698 273978
rect 303238 274294 303294 274350
rect 303362 274294 303418 274350
rect 303238 274170 303294 274226
rect 303362 274170 303418 274226
rect 303238 274046 303294 274102
rect 303362 274046 303418 274102
rect 303238 273922 303294 273978
rect 303362 273922 303418 273978
rect 262220 272942 262276 272998
rect 263788 271502 263844 271558
rect 263900 270782 263956 270838
rect 262108 270242 262164 270298
rect 263788 268802 263844 268858
rect 263788 268442 263844 268498
rect 254994 262294 255050 262350
rect 255118 262294 255174 262350
rect 255242 262294 255298 262350
rect 255366 262294 255422 262350
rect 254994 262170 255050 262226
rect 255118 262170 255174 262226
rect 255242 262170 255298 262226
rect 255366 262170 255422 262226
rect 254994 262046 255050 262102
rect 255118 262046 255174 262102
rect 255242 262046 255298 262102
rect 255366 262046 255422 262102
rect 254994 261922 255050 261978
rect 255118 261922 255174 261978
rect 255242 261922 255298 261978
rect 255366 261922 255422 261978
rect 251274 256294 251330 256350
rect 251398 256294 251454 256350
rect 251522 256294 251578 256350
rect 251646 256294 251702 256350
rect 251274 256170 251330 256226
rect 251398 256170 251454 256226
rect 251522 256170 251578 256226
rect 251646 256170 251702 256226
rect 251274 256046 251330 256102
rect 251398 256046 251454 256102
rect 251522 256046 251578 256102
rect 251646 256046 251702 256102
rect 251274 255922 251330 255978
rect 251398 255922 251454 255978
rect 251522 255922 251578 255978
rect 251646 255922 251702 255978
rect 224274 244294 224330 244350
rect 224398 244294 224454 244350
rect 224522 244294 224578 244350
rect 224646 244294 224702 244350
rect 224274 244170 224330 244226
rect 224398 244170 224454 244226
rect 224522 244170 224578 244226
rect 224646 244170 224702 244226
rect 224274 244046 224330 244102
rect 224398 244046 224454 244102
rect 224522 244046 224578 244102
rect 224646 244046 224702 244102
rect 224274 243922 224330 243978
rect 224398 243922 224454 243978
rect 224522 243922 224578 243978
rect 224646 243922 224702 243978
rect 251274 238294 251330 238350
rect 251398 238294 251454 238350
rect 251522 238294 251578 238350
rect 251646 238294 251702 238350
rect 251274 238170 251330 238226
rect 251398 238170 251454 238226
rect 251522 238170 251578 238226
rect 251646 238170 251702 238226
rect 251274 238046 251330 238102
rect 251398 238046 251454 238102
rect 251522 238046 251578 238102
rect 251646 238046 251702 238102
rect 251274 237922 251330 237978
rect 251398 237922 251454 237978
rect 251522 237922 251578 237978
rect 251646 237922 251702 237978
rect 224274 226294 224330 226350
rect 224398 226294 224454 226350
rect 224522 226294 224578 226350
rect 224646 226294 224702 226350
rect 224274 226170 224330 226226
rect 224398 226170 224454 226226
rect 224522 226170 224578 226226
rect 224646 226170 224702 226226
rect 224274 226046 224330 226102
rect 224398 226046 224454 226102
rect 224522 226046 224578 226102
rect 224646 226046 224702 226102
rect 224274 225922 224330 225978
rect 224398 225922 224454 225978
rect 224522 225922 224578 225978
rect 224646 225922 224702 225978
rect 251274 220294 251330 220350
rect 251398 220294 251454 220350
rect 251522 220294 251578 220350
rect 251646 220294 251702 220350
rect 251274 220170 251330 220226
rect 251398 220170 251454 220226
rect 251522 220170 251578 220226
rect 251646 220170 251702 220226
rect 251274 220046 251330 220102
rect 251398 220046 251454 220102
rect 251522 220046 251578 220102
rect 251646 220046 251702 220102
rect 251274 219922 251330 219978
rect 251398 219922 251454 219978
rect 251522 219922 251578 219978
rect 251646 219922 251702 219978
rect 224274 208294 224330 208350
rect 224398 208294 224454 208350
rect 224522 208294 224578 208350
rect 224646 208294 224702 208350
rect 224274 208170 224330 208226
rect 224398 208170 224454 208226
rect 224522 208170 224578 208226
rect 224646 208170 224702 208226
rect 224274 208046 224330 208102
rect 224398 208046 224454 208102
rect 224522 208046 224578 208102
rect 224646 208046 224702 208102
rect 224274 207922 224330 207978
rect 224398 207922 224454 207978
rect 224522 207922 224578 207978
rect 224646 207922 224702 207978
rect 225878 208294 225934 208350
rect 226002 208294 226058 208350
rect 225878 208170 225934 208226
rect 226002 208170 226058 208226
rect 225878 208046 225934 208102
rect 226002 208046 226058 208102
rect 225878 207922 225934 207978
rect 226002 207922 226058 207978
rect 241238 202294 241294 202350
rect 241362 202294 241418 202350
rect 241238 202170 241294 202226
rect 241362 202170 241418 202226
rect 241238 202046 241294 202102
rect 241362 202046 241418 202102
rect 241238 201922 241294 201978
rect 241362 201922 241418 201978
rect 259980 264662 260036 264718
rect 260316 261602 260372 261658
rect 263788 267002 263844 267058
rect 263788 266462 263844 266518
rect 262556 264842 262612 264898
rect 263788 260342 263844 260398
rect 263900 260162 263956 260218
rect 263788 258542 263844 258598
rect 263900 258362 263956 258418
rect 287878 262294 287934 262350
rect 288002 262294 288058 262350
rect 287878 262170 287934 262226
rect 288002 262170 288058 262226
rect 287878 262046 287934 262102
rect 288002 262046 288058 262102
rect 287878 261922 287934 261978
rect 288002 261922 288058 261978
rect 318598 262294 318654 262350
rect 318722 262294 318778 262350
rect 318598 262170 318654 262226
rect 318722 262170 318778 262226
rect 318598 262046 318654 262102
rect 318722 262046 318778 262102
rect 318598 261922 318654 261978
rect 318722 261922 318778 261978
rect 272518 256294 272574 256350
rect 272642 256294 272698 256350
rect 272518 256170 272574 256226
rect 272642 256170 272698 256226
rect 272518 256046 272574 256102
rect 272642 256046 272698 256102
rect 272518 255922 272574 255978
rect 272642 255922 272698 255978
rect 303238 256294 303294 256350
rect 303362 256294 303418 256350
rect 303238 256170 303294 256226
rect 303362 256170 303418 256226
rect 303238 256046 303294 256102
rect 303362 256046 303418 256102
rect 303238 255922 303294 255978
rect 303362 255922 303418 255978
rect 263788 255302 263844 255358
rect 260316 254402 260372 254458
rect 263788 253502 263844 253558
rect 263900 253322 263956 253378
rect 263788 251882 263844 251938
rect 263788 250262 263844 250318
rect 254994 244294 255050 244350
rect 255118 244294 255174 244350
rect 255242 244294 255298 244350
rect 255366 244294 255422 244350
rect 254994 244170 255050 244226
rect 255118 244170 255174 244226
rect 255242 244170 255298 244226
rect 255366 244170 255422 244226
rect 254994 244046 255050 244102
rect 255118 244046 255174 244102
rect 255242 244046 255298 244102
rect 255366 244046 255422 244102
rect 254994 243922 255050 243978
rect 255118 243922 255174 243978
rect 255242 243922 255298 243978
rect 255366 243922 255422 243978
rect 287878 244294 287934 244350
rect 288002 244294 288058 244350
rect 287878 244170 287934 244226
rect 288002 244170 288058 244226
rect 287878 244046 287934 244102
rect 288002 244046 288058 244102
rect 287878 243922 287934 243978
rect 288002 243922 288058 243978
rect 318598 244294 318654 244350
rect 318722 244294 318778 244350
rect 318598 244170 318654 244226
rect 318722 244170 318778 244226
rect 318598 244046 318654 244102
rect 318722 244046 318778 244102
rect 318598 243922 318654 243978
rect 318722 243922 318778 243978
rect 254994 226294 255050 226350
rect 255118 226294 255174 226350
rect 255242 226294 255298 226350
rect 255366 226294 255422 226350
rect 254994 226170 255050 226226
rect 255118 226170 255174 226226
rect 255242 226170 255298 226226
rect 255366 226170 255422 226226
rect 254994 226046 255050 226102
rect 255118 226046 255174 226102
rect 255242 226046 255298 226102
rect 255366 226046 255422 226102
rect 254994 225922 255050 225978
rect 255118 225922 255174 225978
rect 255242 225922 255298 225978
rect 255366 225922 255422 225978
rect 251274 202294 251330 202350
rect 251398 202294 251454 202350
rect 251522 202294 251578 202350
rect 251646 202294 251702 202350
rect 251274 202170 251330 202226
rect 251398 202170 251454 202226
rect 251522 202170 251578 202226
rect 251646 202170 251702 202226
rect 251274 202046 251330 202102
rect 251398 202046 251454 202102
rect 251522 202046 251578 202102
rect 251646 202046 251702 202102
rect 251274 201922 251330 201978
rect 251398 201922 251454 201978
rect 251522 201922 251578 201978
rect 251646 201922 251702 201978
rect 248556 196442 248612 196498
rect 248556 194102 248612 194158
rect 224274 190294 224330 190350
rect 224398 190294 224454 190350
rect 224522 190294 224578 190350
rect 224646 190294 224702 190350
rect 224274 190170 224330 190226
rect 224398 190170 224454 190226
rect 224522 190170 224578 190226
rect 224646 190170 224702 190226
rect 224274 190046 224330 190102
rect 224398 190046 224454 190102
rect 224522 190046 224578 190102
rect 224646 190046 224702 190102
rect 224274 189922 224330 189978
rect 224398 189922 224454 189978
rect 224522 189922 224578 189978
rect 224646 189922 224702 189978
rect 225878 190294 225934 190350
rect 226002 190294 226058 190350
rect 225878 190170 225934 190226
rect 226002 190170 226058 190226
rect 225878 190046 225934 190102
rect 226002 190046 226058 190102
rect 225878 189922 225934 189978
rect 226002 189922 226058 189978
rect 241238 184294 241294 184350
rect 241362 184294 241418 184350
rect 241238 184170 241294 184226
rect 241362 184170 241418 184226
rect 241238 184046 241294 184102
rect 241362 184046 241418 184102
rect 241238 183922 241294 183978
rect 241362 183922 241418 183978
rect 254994 208294 255050 208350
rect 255118 208294 255174 208350
rect 255242 208294 255298 208350
rect 255366 208294 255422 208350
rect 254994 208170 255050 208226
rect 255118 208170 255174 208226
rect 255242 208170 255298 208226
rect 255366 208170 255422 208226
rect 254994 208046 255050 208102
rect 255118 208046 255174 208102
rect 255242 208046 255298 208102
rect 255366 208046 255422 208102
rect 254994 207922 255050 207978
rect 255118 207922 255174 207978
rect 255242 207922 255298 207978
rect 255366 207922 255422 207978
rect 254994 190294 255050 190350
rect 255118 190294 255174 190350
rect 255242 190294 255298 190350
rect 255366 190294 255422 190350
rect 254994 190170 255050 190226
rect 255118 190170 255174 190226
rect 255242 190170 255298 190226
rect 255366 190170 255422 190226
rect 254994 190046 255050 190102
rect 255118 190046 255174 190102
rect 255242 190046 255298 190102
rect 255366 190046 255422 190102
rect 254994 189922 255050 189978
rect 255118 189922 255174 189978
rect 255242 189922 255298 189978
rect 255366 189922 255422 189978
rect 251274 184294 251330 184350
rect 251398 184294 251454 184350
rect 251522 184294 251578 184350
rect 251646 184294 251702 184350
rect 251274 184170 251330 184226
rect 251398 184170 251454 184226
rect 251522 184170 251578 184226
rect 251646 184170 251702 184226
rect 251274 184046 251330 184102
rect 251398 184046 251454 184102
rect 251522 184046 251578 184102
rect 251646 184046 251702 184102
rect 251274 183922 251330 183978
rect 251398 183922 251454 183978
rect 251522 183922 251578 183978
rect 251646 183922 251702 183978
rect 224274 172294 224330 172350
rect 224398 172294 224454 172350
rect 224522 172294 224578 172350
rect 224646 172294 224702 172350
rect 224274 172170 224330 172226
rect 224398 172170 224454 172226
rect 224522 172170 224578 172226
rect 224646 172170 224702 172226
rect 224274 172046 224330 172102
rect 224398 172046 224454 172102
rect 224522 172046 224578 172102
rect 224646 172046 224702 172102
rect 224274 171922 224330 171978
rect 224398 171922 224454 171978
rect 224522 171922 224578 171978
rect 224646 171922 224702 171978
rect 224274 154294 224330 154350
rect 224398 154294 224454 154350
rect 224522 154294 224578 154350
rect 224646 154294 224702 154350
rect 224274 154170 224330 154226
rect 224398 154170 224454 154226
rect 224522 154170 224578 154226
rect 224646 154170 224702 154226
rect 224274 154046 224330 154102
rect 224398 154046 224454 154102
rect 224522 154046 224578 154102
rect 224646 154046 224702 154102
rect 224274 153922 224330 153978
rect 224398 153922 224454 153978
rect 224522 153922 224578 153978
rect 224646 153922 224702 153978
rect 251274 166294 251330 166350
rect 251398 166294 251454 166350
rect 251522 166294 251578 166350
rect 251646 166294 251702 166350
rect 251274 166170 251330 166226
rect 251398 166170 251454 166226
rect 251522 166170 251578 166226
rect 251646 166170 251702 166226
rect 251274 166046 251330 166102
rect 251398 166046 251454 166102
rect 251522 166046 251578 166102
rect 251646 166046 251702 166102
rect 251274 165922 251330 165978
rect 251398 165922 251454 165978
rect 251522 165922 251578 165978
rect 251646 165922 251702 165978
rect 251274 148294 251330 148350
rect 251398 148294 251454 148350
rect 251522 148294 251578 148350
rect 251646 148294 251702 148350
rect 251274 148170 251330 148226
rect 251398 148170 251454 148226
rect 251522 148170 251578 148226
rect 251646 148170 251702 148226
rect 251274 148046 251330 148102
rect 251398 148046 251454 148102
rect 251522 148046 251578 148102
rect 251646 148046 251702 148102
rect 251274 147922 251330 147978
rect 251398 147922 251454 147978
rect 251522 147922 251578 147978
rect 251646 147922 251702 147978
rect 224274 136294 224330 136350
rect 224398 136294 224454 136350
rect 224522 136294 224578 136350
rect 224646 136294 224702 136350
rect 224274 136170 224330 136226
rect 224398 136170 224454 136226
rect 224522 136170 224578 136226
rect 224646 136170 224702 136226
rect 224274 136046 224330 136102
rect 224398 136046 224454 136102
rect 224522 136046 224578 136102
rect 224646 136046 224702 136102
rect 224274 135922 224330 135978
rect 224398 135922 224454 135978
rect 224522 135922 224578 135978
rect 224646 135922 224702 135978
rect 225878 136294 225934 136350
rect 226002 136294 226058 136350
rect 225878 136170 225934 136226
rect 226002 136170 226058 136226
rect 225878 136046 225934 136102
rect 226002 136046 226058 136102
rect 225878 135922 225934 135978
rect 226002 135922 226058 135978
rect 241238 130294 241294 130350
rect 241362 130294 241418 130350
rect 241238 130170 241294 130226
rect 241362 130170 241418 130226
rect 241238 130046 241294 130102
rect 241362 130046 241418 130102
rect 241238 129922 241294 129978
rect 241362 129922 241418 129978
rect 251274 130294 251330 130350
rect 251398 130294 251454 130350
rect 251522 130294 251578 130350
rect 251646 130294 251702 130350
rect 251274 130170 251330 130226
rect 251398 130170 251454 130226
rect 251522 130170 251578 130226
rect 251646 130170 251702 130226
rect 251274 130046 251330 130102
rect 251398 130046 251454 130102
rect 251522 130046 251578 130102
rect 251646 130046 251702 130102
rect 251274 129922 251330 129978
rect 251398 129922 251454 129978
rect 251522 129922 251578 129978
rect 251646 129922 251702 129978
rect 224274 118294 224330 118350
rect 224398 118294 224454 118350
rect 224522 118294 224578 118350
rect 224646 118294 224702 118350
rect 224274 118170 224330 118226
rect 224398 118170 224454 118226
rect 224522 118170 224578 118226
rect 224646 118170 224702 118226
rect 224274 118046 224330 118102
rect 224398 118046 224454 118102
rect 224522 118046 224578 118102
rect 224646 118046 224702 118102
rect 224274 117922 224330 117978
rect 224398 117922 224454 117978
rect 224522 117922 224578 117978
rect 224646 117922 224702 117978
rect 225878 118294 225934 118350
rect 226002 118294 226058 118350
rect 225878 118170 225934 118226
rect 226002 118170 226058 118226
rect 225878 118046 225934 118102
rect 226002 118046 226058 118102
rect 225878 117922 225934 117978
rect 226002 117922 226058 117978
rect 241238 112294 241294 112350
rect 241362 112294 241418 112350
rect 241238 112170 241294 112226
rect 241362 112170 241418 112226
rect 241238 112046 241294 112102
rect 241362 112046 241418 112102
rect 241238 111922 241294 111978
rect 241362 111922 241418 111978
rect 272518 238294 272574 238350
rect 272642 238294 272698 238350
rect 272518 238170 272574 238226
rect 272642 238170 272698 238226
rect 272518 238046 272574 238102
rect 272642 238046 272698 238102
rect 272518 237922 272574 237978
rect 272642 237922 272698 237978
rect 303238 238294 303294 238350
rect 303362 238294 303418 238350
rect 303238 238170 303294 238226
rect 303362 238170 303418 238226
rect 303238 238046 303294 238102
rect 303362 238046 303418 238102
rect 303238 237922 303294 237978
rect 303362 237922 303418 237978
rect 262108 205802 262164 205858
rect 287878 226294 287934 226350
rect 288002 226294 288058 226350
rect 287878 226170 287934 226226
rect 288002 226170 288058 226226
rect 287878 226046 287934 226102
rect 288002 226046 288058 226102
rect 287878 225922 287934 225978
rect 288002 225922 288058 225978
rect 318598 226294 318654 226350
rect 318722 226294 318778 226350
rect 318598 226170 318654 226226
rect 318722 226170 318778 226226
rect 318598 226046 318654 226102
rect 318722 226046 318778 226102
rect 318598 225922 318654 225978
rect 318722 225922 318778 225978
rect 272518 220294 272574 220350
rect 272642 220294 272698 220350
rect 272518 220170 272574 220226
rect 272642 220170 272698 220226
rect 272518 220046 272574 220102
rect 272642 220046 272698 220102
rect 272518 219922 272574 219978
rect 272642 219922 272698 219978
rect 303238 220294 303294 220350
rect 303362 220294 303418 220350
rect 303238 220170 303294 220226
rect 303362 220170 303418 220226
rect 303238 220046 303294 220102
rect 303362 220046 303418 220102
rect 303238 219922 303294 219978
rect 303362 219922 303418 219978
rect 287878 208294 287934 208350
rect 288002 208294 288058 208350
rect 287878 208170 287934 208226
rect 288002 208170 288058 208226
rect 287878 208046 287934 208102
rect 288002 208046 288058 208102
rect 287878 207922 287934 207978
rect 288002 207922 288058 207978
rect 318598 208294 318654 208350
rect 318722 208294 318778 208350
rect 318598 208170 318654 208226
rect 318722 208170 318778 208226
rect 318598 208046 318654 208102
rect 318722 208046 318778 208102
rect 318598 207922 318654 207978
rect 318722 207922 318778 207978
rect 263788 198242 263844 198298
rect 263788 196802 263844 196858
rect 263900 196622 263956 196678
rect 263788 195002 263844 195058
rect 262108 193202 262164 193258
rect 263788 192122 263844 192178
rect 263788 189602 263844 189658
rect 263900 189422 263956 189478
rect 263900 187442 263956 187498
rect 258636 186362 258692 186418
rect 258412 186182 258468 186238
rect 263788 186002 263844 186058
rect 272518 202294 272574 202350
rect 272642 202294 272698 202350
rect 272518 202170 272574 202226
rect 272642 202170 272698 202226
rect 272518 202046 272574 202102
rect 272642 202046 272698 202102
rect 272518 201922 272574 201978
rect 272642 201922 272698 201978
rect 303238 202294 303294 202350
rect 303362 202294 303418 202350
rect 303238 202170 303294 202226
rect 303362 202170 303418 202226
rect 303238 202046 303294 202102
rect 303362 202046 303418 202102
rect 303238 201922 303294 201978
rect 303362 201922 303418 201978
rect 287878 190294 287934 190350
rect 288002 190294 288058 190350
rect 287878 190170 287934 190226
rect 288002 190170 288058 190226
rect 287878 190046 287934 190102
rect 288002 190046 288058 190102
rect 287878 189922 287934 189978
rect 288002 189922 288058 189978
rect 318598 190294 318654 190350
rect 318722 190294 318778 190350
rect 318598 190170 318654 190226
rect 318722 190170 318778 190226
rect 318598 190046 318654 190102
rect 318722 190046 318778 190102
rect 318598 189922 318654 189978
rect 318722 189922 318778 189978
rect 264012 187262 264068 187318
rect 272518 184294 272574 184350
rect 272642 184294 272698 184350
rect 272518 184170 272574 184226
rect 272642 184170 272698 184226
rect 272518 184046 272574 184102
rect 272642 184046 272698 184102
rect 272518 183922 272574 183978
rect 272642 183922 272698 183978
rect 303238 184294 303294 184350
rect 303362 184294 303418 184350
rect 303238 184170 303294 184226
rect 303362 184170 303418 184226
rect 303238 184046 303294 184102
rect 303362 184046 303418 184102
rect 303238 183922 303294 183978
rect 303362 183922 303418 183978
rect 254994 172294 255050 172350
rect 255118 172294 255174 172350
rect 255242 172294 255298 172350
rect 255366 172294 255422 172350
rect 254994 172170 255050 172226
rect 255118 172170 255174 172226
rect 255242 172170 255298 172226
rect 255366 172170 255422 172226
rect 254994 172046 255050 172102
rect 255118 172046 255174 172102
rect 255242 172046 255298 172102
rect 255366 172046 255422 172102
rect 254994 171922 255050 171978
rect 255118 171922 255174 171978
rect 255242 171922 255298 171978
rect 255366 171922 255422 171978
rect 254994 154294 255050 154350
rect 255118 154294 255174 154350
rect 255242 154294 255298 154350
rect 255366 154294 255422 154350
rect 254994 154170 255050 154226
rect 255118 154170 255174 154226
rect 255242 154170 255298 154226
rect 255366 154170 255422 154226
rect 254994 154046 255050 154102
rect 255118 154046 255174 154102
rect 255242 154046 255298 154102
rect 255366 154046 255422 154102
rect 254994 153922 255050 153978
rect 255118 153922 255174 153978
rect 255242 153922 255298 153978
rect 255366 153922 255422 153978
rect 254994 136294 255050 136350
rect 255118 136294 255174 136350
rect 255242 136294 255298 136350
rect 255366 136294 255422 136350
rect 254994 136170 255050 136226
rect 255118 136170 255174 136226
rect 255242 136170 255298 136226
rect 255366 136170 255422 136226
rect 254994 136046 255050 136102
rect 255118 136046 255174 136102
rect 255242 136046 255298 136102
rect 255366 136046 255422 136102
rect 254994 135922 255050 135978
rect 255118 135922 255174 135978
rect 255242 135922 255298 135978
rect 255366 135922 255422 135978
rect 251274 112294 251330 112350
rect 251398 112294 251454 112350
rect 251522 112294 251578 112350
rect 251646 112294 251702 112350
rect 251274 112170 251330 112226
rect 251398 112170 251454 112226
rect 251522 112170 251578 112226
rect 251646 112170 251702 112226
rect 251274 112046 251330 112102
rect 251398 112046 251454 112102
rect 251522 112046 251578 112102
rect 251646 112046 251702 112102
rect 251274 111922 251330 111978
rect 251398 111922 251454 111978
rect 251522 111922 251578 111978
rect 251646 111922 251702 111978
rect 224274 100294 224330 100350
rect 224398 100294 224454 100350
rect 224522 100294 224578 100350
rect 224646 100294 224702 100350
rect 224274 100170 224330 100226
rect 224398 100170 224454 100226
rect 224522 100170 224578 100226
rect 224646 100170 224702 100226
rect 224274 100046 224330 100102
rect 224398 100046 224454 100102
rect 224522 100046 224578 100102
rect 224646 100046 224702 100102
rect 224274 99922 224330 99978
rect 224398 99922 224454 99978
rect 224522 99922 224578 99978
rect 224646 99922 224702 99978
rect 224274 82294 224330 82350
rect 224398 82294 224454 82350
rect 224522 82294 224578 82350
rect 224646 82294 224702 82350
rect 224274 82170 224330 82226
rect 224398 82170 224454 82226
rect 224522 82170 224578 82226
rect 224646 82170 224702 82226
rect 224274 82046 224330 82102
rect 224398 82046 224454 82102
rect 224522 82046 224578 82102
rect 224646 82046 224702 82102
rect 224274 81922 224330 81978
rect 224398 81922 224454 81978
rect 224522 81922 224578 81978
rect 224646 81922 224702 81978
rect 251274 94294 251330 94350
rect 251398 94294 251454 94350
rect 251522 94294 251578 94350
rect 251646 94294 251702 94350
rect 251274 94170 251330 94226
rect 251398 94170 251454 94226
rect 251522 94170 251578 94226
rect 251646 94170 251702 94226
rect 251274 94046 251330 94102
rect 251398 94046 251454 94102
rect 251522 94046 251578 94102
rect 251646 94046 251702 94102
rect 251274 93922 251330 93978
rect 251398 93922 251454 93978
rect 251522 93922 251578 93978
rect 251646 93922 251702 93978
rect 251274 76294 251330 76350
rect 251398 76294 251454 76350
rect 251522 76294 251578 76350
rect 251646 76294 251702 76350
rect 251274 76170 251330 76226
rect 251398 76170 251454 76226
rect 251522 76170 251578 76226
rect 251646 76170 251702 76226
rect 251274 76046 251330 76102
rect 251398 76046 251454 76102
rect 251522 76046 251578 76102
rect 251646 76046 251702 76102
rect 251274 75922 251330 75978
rect 251398 75922 251454 75978
rect 251522 75922 251578 75978
rect 251646 75922 251702 75978
rect 224274 64294 224330 64350
rect 224398 64294 224454 64350
rect 224522 64294 224578 64350
rect 224646 64294 224702 64350
rect 224274 64170 224330 64226
rect 224398 64170 224454 64226
rect 224522 64170 224578 64226
rect 224646 64170 224702 64226
rect 224274 64046 224330 64102
rect 224398 64046 224454 64102
rect 224522 64046 224578 64102
rect 224646 64046 224702 64102
rect 224274 63922 224330 63978
rect 224398 63922 224454 63978
rect 224522 63922 224578 63978
rect 224646 63922 224702 63978
rect 225878 64294 225934 64350
rect 226002 64294 226058 64350
rect 225878 64170 225934 64226
rect 226002 64170 226058 64226
rect 225878 64046 225934 64102
rect 226002 64046 226058 64102
rect 225878 63922 225934 63978
rect 226002 63922 226058 63978
rect 241238 58294 241294 58350
rect 241362 58294 241418 58350
rect 241238 58170 241294 58226
rect 241362 58170 241418 58226
rect 241238 58046 241294 58102
rect 241362 58046 241418 58102
rect 241238 57922 241294 57978
rect 241362 57922 241418 57978
rect 251274 58294 251330 58350
rect 251398 58294 251454 58350
rect 251522 58294 251578 58350
rect 251646 58294 251702 58350
rect 251274 58170 251330 58226
rect 251398 58170 251454 58226
rect 251522 58170 251578 58226
rect 251646 58170 251702 58226
rect 251274 58046 251330 58102
rect 251398 58046 251454 58102
rect 251522 58046 251578 58102
rect 251646 58046 251702 58102
rect 251274 57922 251330 57978
rect 251398 57922 251454 57978
rect 251522 57922 251578 57978
rect 251646 57922 251702 57978
rect 224274 46294 224330 46350
rect 224398 46294 224454 46350
rect 224522 46294 224578 46350
rect 224646 46294 224702 46350
rect 224274 46170 224330 46226
rect 224398 46170 224454 46226
rect 224522 46170 224578 46226
rect 224646 46170 224702 46226
rect 224274 46046 224330 46102
rect 224398 46046 224454 46102
rect 224522 46046 224578 46102
rect 224646 46046 224702 46102
rect 224274 45922 224330 45978
rect 224398 45922 224454 45978
rect 224522 45922 224578 45978
rect 224646 45922 224702 45978
rect 225878 46294 225934 46350
rect 226002 46294 226058 46350
rect 225878 46170 225934 46226
rect 226002 46170 226058 46226
rect 225878 46046 225934 46102
rect 226002 46046 226058 46102
rect 225878 45922 225934 45978
rect 226002 45922 226058 45978
rect 241238 40294 241294 40350
rect 241362 40294 241418 40350
rect 241238 40170 241294 40226
rect 241362 40170 241418 40226
rect 241238 40046 241294 40102
rect 241362 40046 241418 40102
rect 241238 39922 241294 39978
rect 241362 39922 241418 39978
rect 254994 118294 255050 118350
rect 255118 118294 255174 118350
rect 255242 118294 255298 118350
rect 255366 118294 255422 118350
rect 254994 118170 255050 118226
rect 255118 118170 255174 118226
rect 255242 118170 255298 118226
rect 255366 118170 255422 118226
rect 254994 118046 255050 118102
rect 255118 118046 255174 118102
rect 255242 118046 255298 118102
rect 255366 118046 255422 118102
rect 254994 117922 255050 117978
rect 255118 117922 255174 117978
rect 255242 117922 255298 117978
rect 255366 117922 255422 117978
rect 254994 100294 255050 100350
rect 255118 100294 255174 100350
rect 255242 100294 255298 100350
rect 255366 100294 255422 100350
rect 254994 100170 255050 100226
rect 255118 100170 255174 100226
rect 255242 100170 255298 100226
rect 255366 100170 255422 100226
rect 254994 100046 255050 100102
rect 255118 100046 255174 100102
rect 255242 100046 255298 100102
rect 255366 100046 255422 100102
rect 254994 99922 255050 99978
rect 255118 99922 255174 99978
rect 255242 99922 255298 99978
rect 255366 99922 255422 99978
rect 254994 82294 255050 82350
rect 255118 82294 255174 82350
rect 255242 82294 255298 82350
rect 255366 82294 255422 82350
rect 254994 82170 255050 82226
rect 255118 82170 255174 82226
rect 255242 82170 255298 82226
rect 255366 82170 255422 82226
rect 254994 82046 255050 82102
rect 255118 82046 255174 82102
rect 255242 82046 255298 82102
rect 255366 82046 255422 82102
rect 254994 81922 255050 81978
rect 255118 81922 255174 81978
rect 255242 81922 255298 81978
rect 255366 81922 255422 81978
rect 254994 64294 255050 64350
rect 255118 64294 255174 64350
rect 255242 64294 255298 64350
rect 255366 64294 255422 64350
rect 254994 64170 255050 64226
rect 255118 64170 255174 64226
rect 255242 64170 255298 64226
rect 255366 64170 255422 64226
rect 254994 64046 255050 64102
rect 255118 64046 255174 64102
rect 255242 64046 255298 64102
rect 255366 64046 255422 64102
rect 254994 63922 255050 63978
rect 255118 63922 255174 63978
rect 255242 63922 255298 63978
rect 255366 63922 255422 63978
rect 259980 117422 260036 117478
rect 263788 137762 263844 137818
rect 263788 132902 263844 132958
rect 263900 132722 263956 132778
rect 263900 131282 263956 131338
rect 263788 128582 263844 128638
rect 287878 172294 287934 172350
rect 288002 172294 288058 172350
rect 287878 172170 287934 172226
rect 288002 172170 288058 172226
rect 287878 172046 287934 172102
rect 288002 172046 288058 172102
rect 287878 171922 287934 171978
rect 288002 171922 288058 171978
rect 318598 172294 318654 172350
rect 318722 172294 318778 172350
rect 318598 172170 318654 172226
rect 318722 172170 318778 172226
rect 318598 172046 318654 172102
rect 318722 172046 318778 172102
rect 318598 171922 318654 171978
rect 318722 171922 318778 171978
rect 272518 166294 272574 166350
rect 272642 166294 272698 166350
rect 272518 166170 272574 166226
rect 272642 166170 272698 166226
rect 272518 166046 272574 166102
rect 272642 166046 272698 166102
rect 272518 165922 272574 165978
rect 272642 165922 272698 165978
rect 303238 166294 303294 166350
rect 303362 166294 303418 166350
rect 303238 166170 303294 166226
rect 303362 166170 303418 166226
rect 303238 166046 303294 166102
rect 303362 166046 303418 166102
rect 303238 165922 303294 165978
rect 303362 165922 303418 165978
rect 287878 154294 287934 154350
rect 288002 154294 288058 154350
rect 287878 154170 287934 154226
rect 288002 154170 288058 154226
rect 287878 154046 287934 154102
rect 288002 154046 288058 154102
rect 287878 153922 287934 153978
rect 288002 153922 288058 153978
rect 318598 154294 318654 154350
rect 318722 154294 318778 154350
rect 318598 154170 318654 154226
rect 318722 154170 318778 154226
rect 318598 154046 318654 154102
rect 318722 154046 318778 154102
rect 318598 153922 318654 153978
rect 318722 153922 318778 153978
rect 272518 148294 272574 148350
rect 272642 148294 272698 148350
rect 272518 148170 272574 148226
rect 272642 148170 272698 148226
rect 272518 148046 272574 148102
rect 272642 148046 272698 148102
rect 272518 147922 272574 147978
rect 272642 147922 272698 147978
rect 303238 148294 303294 148350
rect 303362 148294 303418 148350
rect 303238 148170 303294 148226
rect 303362 148170 303418 148226
rect 303238 148046 303294 148102
rect 303362 148046 303418 148102
rect 303238 147922 303294 147978
rect 303362 147922 303418 147978
rect 287878 136294 287934 136350
rect 288002 136294 288058 136350
rect 287878 136170 287934 136226
rect 288002 136170 288058 136226
rect 287878 136046 287934 136102
rect 288002 136046 288058 136102
rect 287878 135922 287934 135978
rect 288002 135922 288058 135978
rect 318598 136294 318654 136350
rect 318722 136294 318778 136350
rect 318598 136170 318654 136226
rect 318722 136170 318778 136226
rect 318598 136046 318654 136102
rect 318722 136046 318778 136102
rect 318598 135922 318654 135978
rect 318722 135922 318778 135978
rect 264796 131102 264852 131158
rect 263900 127862 263956 127918
rect 263788 126062 263844 126118
rect 263900 125162 263956 125218
rect 264012 121742 264068 121798
rect 272518 130294 272574 130350
rect 272642 130294 272698 130350
rect 272518 130170 272574 130226
rect 272642 130170 272698 130226
rect 272518 130046 272574 130102
rect 272642 130046 272698 130102
rect 272518 129922 272574 129978
rect 272642 129922 272698 129978
rect 303238 130294 303294 130350
rect 303362 130294 303418 130350
rect 303238 130170 303294 130226
rect 303362 130170 303418 130226
rect 303238 130046 303294 130102
rect 303362 130046 303418 130102
rect 303238 129922 303294 129978
rect 303362 129922 303418 129978
rect 287878 118294 287934 118350
rect 288002 118294 288058 118350
rect 287878 118170 287934 118226
rect 288002 118170 288058 118226
rect 287878 118046 287934 118102
rect 288002 118046 288058 118102
rect 287878 117922 287934 117978
rect 288002 117922 288058 117978
rect 318598 118294 318654 118350
rect 318722 118294 318778 118350
rect 318598 118170 318654 118226
rect 318722 118170 318778 118226
rect 318598 118046 318654 118102
rect 318722 118046 318778 118102
rect 318598 117922 318654 117978
rect 318722 117922 318778 117978
rect 272518 112294 272574 112350
rect 272642 112294 272698 112350
rect 272518 112170 272574 112226
rect 272642 112170 272698 112226
rect 272518 112046 272574 112102
rect 272642 112046 272698 112102
rect 272518 111922 272574 111978
rect 272642 111922 272698 111978
rect 303238 112294 303294 112350
rect 303362 112294 303418 112350
rect 303238 112170 303294 112226
rect 303362 112170 303418 112226
rect 303238 112046 303294 112102
rect 303362 112046 303418 112102
rect 303238 111922 303294 111978
rect 303362 111922 303418 111978
rect 287878 100294 287934 100350
rect 288002 100294 288058 100350
rect 287878 100170 287934 100226
rect 288002 100170 288058 100226
rect 287878 100046 287934 100102
rect 288002 100046 288058 100102
rect 287878 99922 287934 99978
rect 288002 99922 288058 99978
rect 318598 100294 318654 100350
rect 318722 100294 318778 100350
rect 318598 100170 318654 100226
rect 318722 100170 318778 100226
rect 318598 100046 318654 100102
rect 318722 100046 318778 100102
rect 318598 99922 318654 99978
rect 318722 99922 318778 99978
rect 272518 94294 272574 94350
rect 272642 94294 272698 94350
rect 272518 94170 272574 94226
rect 272642 94170 272698 94226
rect 272518 94046 272574 94102
rect 272642 94046 272698 94102
rect 272518 93922 272574 93978
rect 272642 93922 272698 93978
rect 303238 94294 303294 94350
rect 303362 94294 303418 94350
rect 303238 94170 303294 94226
rect 303362 94170 303418 94226
rect 303238 94046 303294 94102
rect 303362 94046 303418 94102
rect 303238 93922 303294 93978
rect 303362 93922 303418 93978
rect 287878 82294 287934 82350
rect 288002 82294 288058 82350
rect 287878 82170 287934 82226
rect 288002 82170 288058 82226
rect 287878 82046 287934 82102
rect 288002 82046 288058 82102
rect 287878 81922 287934 81978
rect 288002 81922 288058 81978
rect 318598 82294 318654 82350
rect 318722 82294 318778 82350
rect 318598 82170 318654 82226
rect 318722 82170 318778 82226
rect 318598 82046 318654 82102
rect 318722 82046 318778 82102
rect 318598 81922 318654 81978
rect 318722 81922 318778 81978
rect 272518 76294 272574 76350
rect 272642 76294 272698 76350
rect 272518 76170 272574 76226
rect 272642 76170 272698 76226
rect 272518 76046 272574 76102
rect 272642 76046 272698 76102
rect 272518 75922 272574 75978
rect 272642 75922 272698 75978
rect 303238 76294 303294 76350
rect 303362 76294 303418 76350
rect 303238 76170 303294 76226
rect 303362 76170 303418 76226
rect 303238 76046 303294 76102
rect 303362 76046 303418 76102
rect 303238 75922 303294 75978
rect 303362 75922 303418 75978
rect 343434 562294 343490 562350
rect 343558 562294 343614 562350
rect 343682 562294 343738 562350
rect 343806 562294 343862 562350
rect 343434 562170 343490 562226
rect 343558 562170 343614 562226
rect 343682 562170 343738 562226
rect 343806 562170 343862 562226
rect 343434 562046 343490 562102
rect 343558 562046 343614 562102
rect 343682 562046 343738 562102
rect 343806 562046 343862 562102
rect 343434 561922 343490 561978
rect 343558 561922 343614 561978
rect 343682 561922 343738 561978
rect 343806 561922 343862 561978
rect 334460 473642 334516 473698
rect 334460 470596 334516 470638
rect 334460 470582 334516 470596
rect 334460 470402 334516 470458
rect 334460 469502 334516 469558
rect 334460 466082 334516 466138
rect 334460 465182 334516 465238
rect 334460 462842 334516 462898
rect 339388 480482 339444 480538
rect 347154 598116 347210 598172
rect 347278 598116 347334 598172
rect 347402 598116 347458 598172
rect 347526 598116 347582 598172
rect 347154 597992 347210 598048
rect 347278 597992 347334 598048
rect 347402 597992 347458 598048
rect 347526 597992 347582 598048
rect 347154 597868 347210 597924
rect 347278 597868 347334 597924
rect 347402 597868 347458 597924
rect 347526 597868 347582 597924
rect 347154 597744 347210 597800
rect 347278 597744 347334 597800
rect 347402 597744 347458 597800
rect 347526 597744 347582 597800
rect 347154 586294 347210 586350
rect 347278 586294 347334 586350
rect 347402 586294 347458 586350
rect 347526 586294 347582 586350
rect 347154 586170 347210 586226
rect 347278 586170 347334 586226
rect 347402 586170 347458 586226
rect 347526 586170 347582 586226
rect 347154 586046 347210 586102
rect 347278 586046 347334 586102
rect 347402 586046 347458 586102
rect 347526 586046 347582 586102
rect 347154 585922 347210 585978
rect 347278 585922 347334 585978
rect 347402 585922 347458 585978
rect 347526 585922 347582 585978
rect 347154 568294 347210 568350
rect 347278 568294 347334 568350
rect 347402 568294 347458 568350
rect 347526 568294 347582 568350
rect 347154 568170 347210 568226
rect 347278 568170 347334 568226
rect 347402 568170 347458 568226
rect 347526 568170 347582 568226
rect 347154 568046 347210 568102
rect 347278 568046 347334 568102
rect 347402 568046 347458 568102
rect 347526 568046 347582 568102
rect 347154 567922 347210 567978
rect 347278 567922 347334 567978
rect 347402 567922 347458 567978
rect 347526 567922 347582 567978
rect 343434 544294 343490 544350
rect 343558 544294 343614 544350
rect 343682 544294 343738 544350
rect 343806 544294 343862 544350
rect 343434 544170 343490 544226
rect 343558 544170 343614 544226
rect 343682 544170 343738 544226
rect 343806 544170 343862 544226
rect 343434 544046 343490 544102
rect 343558 544046 343614 544102
rect 343682 544046 343738 544102
rect 343806 544046 343862 544102
rect 343434 543922 343490 543978
rect 343558 543922 343614 543978
rect 343682 543922 343738 543978
rect 343806 543922 343862 543978
rect 343434 526294 343490 526350
rect 343558 526294 343614 526350
rect 343682 526294 343738 526350
rect 343806 526294 343862 526350
rect 343434 526170 343490 526226
rect 343558 526170 343614 526226
rect 343682 526170 343738 526226
rect 343806 526170 343862 526226
rect 343434 526046 343490 526102
rect 343558 526046 343614 526102
rect 343682 526046 343738 526102
rect 343806 526046 343862 526102
rect 343434 525922 343490 525978
rect 343558 525922 343614 525978
rect 343682 525922 343738 525978
rect 343806 525922 343862 525978
rect 343434 508294 343490 508350
rect 343558 508294 343614 508350
rect 343682 508294 343738 508350
rect 343806 508294 343862 508350
rect 343434 508170 343490 508226
rect 343558 508170 343614 508226
rect 343682 508170 343738 508226
rect 343806 508170 343862 508226
rect 343434 508046 343490 508102
rect 343558 508046 343614 508102
rect 343682 508046 343738 508102
rect 343806 508046 343862 508102
rect 343434 507922 343490 507978
rect 343558 507922 343614 507978
rect 343682 507922 343738 507978
rect 343806 507922 343862 507978
rect 343434 490294 343490 490350
rect 343558 490294 343614 490350
rect 343682 490294 343738 490350
rect 343806 490294 343862 490350
rect 343434 490170 343490 490226
rect 343558 490170 343614 490226
rect 343682 490170 343738 490226
rect 343806 490170 343862 490226
rect 343434 490046 343490 490102
rect 343558 490046 343614 490102
rect 343682 490046 343738 490102
rect 343806 490046 343862 490102
rect 343434 489922 343490 489978
rect 343558 489922 343614 489978
rect 343682 489922 343738 489978
rect 343806 489922 343862 489978
rect 374154 597156 374210 597212
rect 374278 597156 374334 597212
rect 374402 597156 374458 597212
rect 374526 597156 374582 597212
rect 374154 597032 374210 597088
rect 374278 597032 374334 597088
rect 374402 597032 374458 597088
rect 374526 597032 374582 597088
rect 374154 596908 374210 596964
rect 374278 596908 374334 596964
rect 374402 596908 374458 596964
rect 374526 596908 374582 596964
rect 374154 596784 374210 596840
rect 374278 596784 374334 596840
rect 374402 596784 374458 596840
rect 374526 596784 374582 596840
rect 374154 580294 374210 580350
rect 374278 580294 374334 580350
rect 374402 580294 374458 580350
rect 374526 580294 374582 580350
rect 374154 580170 374210 580226
rect 374278 580170 374334 580226
rect 374402 580170 374458 580226
rect 374526 580170 374582 580226
rect 374154 580046 374210 580102
rect 374278 580046 374334 580102
rect 374402 580046 374458 580102
rect 374526 580046 374582 580102
rect 374154 579922 374210 579978
rect 374278 579922 374334 579978
rect 374402 579922 374458 579978
rect 374526 579922 374582 579978
rect 356518 562294 356574 562350
rect 356642 562294 356698 562350
rect 356518 562170 356574 562226
rect 356642 562170 356698 562226
rect 356518 562046 356574 562102
rect 356642 562046 356698 562102
rect 356518 561922 356574 561978
rect 356642 561922 356698 561978
rect 374154 562294 374210 562350
rect 374278 562294 374334 562350
rect 374402 562294 374458 562350
rect 374526 562294 374582 562350
rect 374154 562170 374210 562226
rect 374278 562170 374334 562226
rect 374402 562170 374458 562226
rect 374526 562170 374582 562226
rect 374154 562046 374210 562102
rect 374278 562046 374334 562102
rect 374402 562046 374458 562102
rect 374526 562046 374582 562102
rect 374154 561922 374210 561978
rect 374278 561922 374334 561978
rect 374402 561922 374458 561978
rect 374526 561922 374582 561978
rect 352716 555212 352772 555238
rect 352716 555182 352772 555212
rect 347154 550294 347210 550350
rect 347278 550294 347334 550350
rect 347402 550294 347458 550350
rect 347526 550294 347582 550350
rect 347154 550170 347210 550226
rect 347278 550170 347334 550226
rect 347402 550170 347458 550226
rect 347526 550170 347582 550226
rect 347154 550046 347210 550102
rect 347278 550046 347334 550102
rect 347402 550046 347458 550102
rect 347526 550046 347582 550102
rect 347154 549922 347210 549978
rect 347278 549922 347334 549978
rect 347402 549922 347458 549978
rect 347526 549922 347582 549978
rect 347154 532294 347210 532350
rect 347278 532294 347334 532350
rect 347402 532294 347458 532350
rect 347526 532294 347582 532350
rect 347154 532170 347210 532226
rect 347278 532170 347334 532226
rect 347402 532170 347458 532226
rect 347526 532170 347582 532226
rect 347154 532046 347210 532102
rect 347278 532046 347334 532102
rect 347402 532046 347458 532102
rect 347526 532046 347582 532102
rect 347154 531922 347210 531978
rect 347278 531922 347334 531978
rect 347402 531922 347458 531978
rect 347526 531922 347582 531978
rect 347154 514294 347210 514350
rect 347278 514294 347334 514350
rect 347402 514294 347458 514350
rect 347526 514294 347582 514350
rect 347154 514170 347210 514226
rect 347278 514170 347334 514226
rect 347402 514170 347458 514226
rect 347526 514170 347582 514226
rect 347154 514046 347210 514102
rect 347278 514046 347334 514102
rect 347402 514046 347458 514102
rect 347526 514046 347582 514102
rect 347154 513922 347210 513978
rect 347278 513922 347334 513978
rect 347402 513922 347458 513978
rect 347526 513922 347582 513978
rect 347154 496294 347210 496350
rect 347278 496294 347334 496350
rect 347402 496294 347458 496350
rect 347526 496294 347582 496350
rect 347154 496170 347210 496226
rect 347278 496170 347334 496226
rect 347402 496170 347458 496226
rect 347526 496170 347582 496226
rect 347154 496046 347210 496102
rect 347278 496046 347334 496102
rect 347402 496046 347458 496102
rect 347526 496046 347582 496102
rect 347154 495922 347210 495978
rect 347278 495922 347334 495978
rect 347402 495922 347458 495978
rect 347526 495922 347582 495978
rect 371878 550294 371934 550350
rect 372002 550294 372058 550350
rect 371878 550170 371934 550226
rect 372002 550170 372058 550226
rect 371878 550046 371934 550102
rect 372002 550046 372058 550102
rect 371878 549922 371934 549978
rect 372002 549922 372058 549978
rect 356518 544294 356574 544350
rect 356642 544294 356698 544350
rect 356518 544170 356574 544226
rect 356642 544170 356698 544226
rect 356518 544046 356574 544102
rect 356642 544046 356698 544102
rect 356518 543922 356574 543978
rect 356642 543922 356698 543978
rect 374154 544294 374210 544350
rect 374278 544294 374334 544350
rect 374402 544294 374458 544350
rect 374526 544294 374582 544350
rect 374154 544170 374210 544226
rect 374278 544170 374334 544226
rect 374402 544170 374458 544226
rect 374526 544170 374582 544226
rect 374154 544046 374210 544102
rect 374278 544046 374334 544102
rect 374402 544046 374458 544102
rect 374526 544046 374582 544102
rect 374154 543922 374210 543978
rect 374278 543922 374334 543978
rect 374402 543922 374458 543978
rect 374526 543922 374582 543978
rect 371878 532294 371934 532350
rect 372002 532294 372058 532350
rect 371878 532170 371934 532226
rect 372002 532170 372058 532226
rect 371878 532046 371934 532102
rect 372002 532046 372058 532102
rect 371878 531922 371934 531978
rect 372002 531922 372058 531978
rect 374154 526294 374210 526350
rect 374278 526294 374334 526350
rect 374402 526294 374458 526350
rect 374526 526294 374582 526350
rect 374154 526170 374210 526226
rect 374278 526170 374334 526226
rect 374402 526170 374458 526226
rect 374526 526170 374582 526226
rect 374154 526046 374210 526102
rect 374278 526046 374334 526102
rect 374402 526046 374458 526102
rect 374526 526046 374582 526102
rect 374154 525922 374210 525978
rect 374278 525922 374334 525978
rect 374402 525922 374458 525978
rect 374526 525922 374582 525978
rect 347154 478294 347210 478350
rect 347278 478294 347334 478350
rect 347402 478294 347458 478350
rect 347526 478294 347582 478350
rect 347154 478170 347210 478226
rect 347278 478170 347334 478226
rect 347402 478170 347458 478226
rect 347526 478170 347582 478226
rect 347154 478046 347210 478102
rect 347278 478046 347334 478102
rect 347402 478046 347458 478102
rect 347526 478046 347582 478102
rect 347154 477922 347210 477978
rect 347278 477922 347334 477978
rect 347402 477922 347458 477978
rect 347526 477922 347582 477978
rect 343434 472294 343490 472350
rect 343558 472294 343614 472350
rect 343682 472294 343738 472350
rect 343806 472294 343862 472350
rect 343434 472170 343490 472226
rect 343558 472170 343614 472226
rect 343682 472170 343738 472226
rect 343806 472170 343862 472226
rect 343434 472046 343490 472102
rect 343558 472046 343614 472102
rect 343682 472046 343738 472102
rect 343806 472046 343862 472102
rect 343434 471922 343490 471978
rect 343558 471922 343614 471978
rect 343682 471922 343738 471978
rect 343806 471922 343862 471978
rect 343434 454294 343490 454350
rect 343558 454294 343614 454350
rect 343682 454294 343738 454350
rect 343806 454294 343862 454350
rect 343434 454170 343490 454226
rect 343558 454170 343614 454226
rect 343682 454170 343738 454226
rect 343806 454170 343862 454226
rect 343434 454046 343490 454102
rect 343558 454046 343614 454102
rect 343682 454046 343738 454102
rect 343806 454046 343862 454102
rect 343434 453922 343490 453978
rect 343558 453922 343614 453978
rect 343682 453922 343738 453978
rect 343806 453922 343862 453978
rect 347154 460294 347210 460350
rect 347278 460294 347334 460350
rect 347402 460294 347458 460350
rect 347526 460294 347582 460350
rect 347154 460170 347210 460226
rect 347278 460170 347334 460226
rect 347402 460170 347458 460226
rect 347526 460170 347582 460226
rect 347154 460046 347210 460102
rect 347278 460046 347334 460102
rect 347402 460046 347458 460102
rect 347526 460046 347582 460102
rect 347154 459922 347210 459978
rect 347278 459922 347334 459978
rect 347402 459922 347458 459978
rect 347526 459922 347582 459978
rect 343434 436294 343490 436350
rect 343558 436294 343614 436350
rect 343682 436294 343738 436350
rect 343806 436294 343862 436350
rect 343434 436170 343490 436226
rect 343558 436170 343614 436226
rect 343682 436170 343738 436226
rect 343806 436170 343862 436226
rect 343434 436046 343490 436102
rect 343558 436046 343614 436102
rect 343682 436046 343738 436102
rect 343806 436046 343862 436102
rect 343434 435922 343490 435978
rect 343558 435922 343614 435978
rect 343682 435922 343738 435978
rect 343806 435922 343862 435978
rect 343434 418294 343490 418350
rect 343558 418294 343614 418350
rect 343682 418294 343738 418350
rect 343806 418294 343862 418350
rect 343434 418170 343490 418226
rect 343558 418170 343614 418226
rect 343682 418170 343738 418226
rect 343806 418170 343862 418226
rect 343434 418046 343490 418102
rect 343558 418046 343614 418102
rect 343682 418046 343738 418102
rect 343806 418046 343862 418102
rect 343434 417922 343490 417978
rect 343558 417922 343614 417978
rect 343682 417922 343738 417978
rect 343806 417922 343862 417978
rect 334460 414962 334516 415018
rect 334460 413702 334516 413758
rect 334460 413522 334516 413578
rect 334348 411722 334404 411778
rect 334460 411902 334516 411958
rect 334460 410642 334516 410698
rect 334460 409562 334516 409618
rect 334460 408122 334516 408178
rect 334460 407402 334516 407458
rect 336252 406682 336308 406738
rect 336028 404702 336084 404758
rect 334460 403262 334516 403318
rect 334460 403082 334516 403138
rect 334460 399662 334516 399718
rect 334460 398042 334516 398098
rect 334460 397862 334516 397918
rect 334460 396422 334516 396478
rect 334348 396242 334404 396298
rect 334460 394622 334516 394678
rect 334460 394442 334516 394498
rect 334460 393002 334516 393058
rect 334460 391562 334516 391618
rect 347154 442294 347210 442350
rect 347278 442294 347334 442350
rect 347402 442294 347458 442350
rect 347526 442294 347582 442350
rect 347154 442170 347210 442226
rect 347278 442170 347334 442226
rect 347402 442170 347458 442226
rect 347526 442170 347582 442226
rect 347154 442046 347210 442102
rect 347278 442046 347334 442102
rect 347402 442046 347458 442102
rect 347526 442046 347582 442102
rect 347154 441922 347210 441978
rect 347278 441922 347334 441978
rect 347402 441922 347458 441978
rect 347526 441922 347582 441978
rect 347154 424294 347210 424350
rect 347278 424294 347334 424350
rect 347402 424294 347458 424350
rect 347526 424294 347582 424350
rect 347154 424170 347210 424226
rect 347278 424170 347334 424226
rect 347402 424170 347458 424226
rect 347526 424170 347582 424226
rect 347154 424046 347210 424102
rect 347278 424046 347334 424102
rect 347402 424046 347458 424102
rect 347526 424046 347582 424102
rect 347154 423922 347210 423978
rect 347278 423922 347334 423978
rect 347402 423922 347458 423978
rect 347526 423922 347582 423978
rect 374154 508294 374210 508350
rect 374278 508294 374334 508350
rect 374402 508294 374458 508350
rect 374526 508294 374582 508350
rect 374154 508170 374210 508226
rect 374278 508170 374334 508226
rect 374402 508170 374458 508226
rect 374526 508170 374582 508226
rect 374154 508046 374210 508102
rect 374278 508046 374334 508102
rect 374402 508046 374458 508102
rect 374526 508046 374582 508102
rect 374154 507922 374210 507978
rect 374278 507922 374334 507978
rect 374402 507922 374458 507978
rect 374526 507922 374582 507978
rect 356518 490294 356574 490350
rect 356642 490294 356698 490350
rect 356518 490170 356574 490226
rect 356642 490170 356698 490226
rect 356518 490046 356574 490102
rect 356642 490046 356698 490102
rect 356518 489922 356574 489978
rect 356642 489922 356698 489978
rect 374154 490294 374210 490350
rect 374278 490294 374334 490350
rect 374402 490294 374458 490350
rect 374526 490294 374582 490350
rect 374154 490170 374210 490226
rect 374278 490170 374334 490226
rect 374402 490170 374458 490226
rect 374526 490170 374582 490226
rect 374154 490046 374210 490102
rect 374278 490046 374334 490102
rect 374402 490046 374458 490102
rect 374526 490046 374582 490102
rect 374154 489922 374210 489978
rect 374278 489922 374334 489978
rect 374402 489922 374458 489978
rect 374526 489922 374582 489978
rect 352716 483002 352772 483058
rect 371878 478294 371934 478350
rect 372002 478294 372058 478350
rect 371878 478170 371934 478226
rect 372002 478170 372058 478226
rect 371878 478046 371934 478102
rect 372002 478046 372058 478102
rect 371878 477922 371934 477978
rect 372002 477922 372058 477978
rect 356518 472294 356574 472350
rect 356642 472294 356698 472350
rect 356518 472170 356574 472226
rect 356642 472170 356698 472226
rect 356518 472046 356574 472102
rect 356642 472046 356698 472102
rect 356518 471922 356574 471978
rect 356642 471922 356698 471978
rect 374154 472294 374210 472350
rect 374278 472294 374334 472350
rect 374402 472294 374458 472350
rect 374526 472294 374582 472350
rect 374154 472170 374210 472226
rect 374278 472170 374334 472226
rect 374402 472170 374458 472226
rect 374526 472170 374582 472226
rect 374154 472046 374210 472102
rect 374278 472046 374334 472102
rect 374402 472046 374458 472102
rect 374526 472046 374582 472102
rect 374154 471922 374210 471978
rect 374278 471922 374334 471978
rect 374402 471922 374458 471978
rect 374526 471922 374582 471978
rect 351036 468602 351092 468658
rect 371878 460294 371934 460350
rect 372002 460294 372058 460350
rect 371878 460170 371934 460226
rect 372002 460170 372058 460226
rect 371878 460046 371934 460102
rect 372002 460046 372058 460102
rect 371878 459922 371934 459978
rect 372002 459922 372058 459978
rect 374154 454294 374210 454350
rect 374278 454294 374334 454350
rect 374402 454294 374458 454350
rect 374526 454294 374582 454350
rect 374154 454170 374210 454226
rect 374278 454170 374334 454226
rect 374402 454170 374458 454226
rect 374526 454170 374582 454226
rect 374154 454046 374210 454102
rect 374278 454046 374334 454102
rect 374402 454046 374458 454102
rect 374526 454046 374582 454102
rect 374154 453922 374210 453978
rect 374278 453922 374334 453978
rect 374402 453922 374458 453978
rect 374526 453922 374582 453978
rect 347154 406294 347210 406350
rect 347278 406294 347334 406350
rect 347402 406294 347458 406350
rect 347526 406294 347582 406350
rect 347154 406170 347210 406226
rect 347278 406170 347334 406226
rect 347402 406170 347458 406226
rect 347526 406170 347582 406226
rect 347154 406046 347210 406102
rect 347278 406046 347334 406102
rect 347402 406046 347458 406102
rect 347526 406046 347582 406102
rect 347154 405922 347210 405978
rect 347278 405922 347334 405978
rect 347402 405922 347458 405978
rect 347526 405922 347582 405978
rect 343434 400294 343490 400350
rect 343558 400294 343614 400350
rect 343682 400294 343738 400350
rect 343806 400294 343862 400350
rect 343434 400170 343490 400226
rect 343558 400170 343614 400226
rect 343682 400170 343738 400226
rect 343806 400170 343862 400226
rect 343434 400046 343490 400102
rect 343558 400046 343614 400102
rect 343682 400046 343738 400102
rect 343806 400046 343862 400102
rect 343434 399922 343490 399978
rect 343558 399922 343614 399978
rect 343682 399922 343738 399978
rect 343806 399922 343862 399978
rect 343434 382294 343490 382350
rect 343558 382294 343614 382350
rect 343682 382294 343738 382350
rect 343806 382294 343862 382350
rect 343434 382170 343490 382226
rect 343558 382170 343614 382226
rect 343682 382170 343738 382226
rect 343806 382170 343862 382226
rect 343434 382046 343490 382102
rect 343558 382046 343614 382102
rect 343682 382046 343738 382102
rect 343806 382046 343862 382102
rect 343434 381922 343490 381978
rect 343558 381922 343614 381978
rect 343682 381922 343738 381978
rect 343806 381922 343862 381978
rect 343434 364294 343490 364350
rect 343558 364294 343614 364350
rect 343682 364294 343738 364350
rect 343806 364294 343862 364350
rect 343434 364170 343490 364226
rect 343558 364170 343614 364226
rect 343682 364170 343738 364226
rect 343806 364170 343862 364226
rect 343434 364046 343490 364102
rect 343558 364046 343614 364102
rect 343682 364046 343738 364102
rect 343806 364046 343862 364102
rect 343434 363922 343490 363978
rect 343558 363922 343614 363978
rect 343682 363922 343738 363978
rect 343806 363922 343862 363978
rect 334460 349442 334516 349498
rect 350252 420002 350308 420058
rect 374154 436294 374210 436350
rect 374278 436294 374334 436350
rect 374402 436294 374458 436350
rect 374526 436294 374582 436350
rect 374154 436170 374210 436226
rect 374278 436170 374334 436226
rect 374402 436170 374458 436226
rect 374526 436170 374582 436226
rect 374154 436046 374210 436102
rect 374278 436046 374334 436102
rect 374402 436046 374458 436102
rect 374526 436046 374582 436102
rect 374154 435922 374210 435978
rect 374278 435922 374334 435978
rect 374402 435922 374458 435978
rect 374526 435922 374582 435978
rect 356518 418294 356574 418350
rect 356642 418294 356698 418350
rect 356518 418170 356574 418226
rect 356642 418170 356698 418226
rect 356518 418046 356574 418102
rect 356642 418046 356698 418102
rect 356518 417922 356574 417978
rect 356642 417922 356698 417978
rect 374154 418294 374210 418350
rect 374278 418294 374334 418350
rect 374402 418294 374458 418350
rect 374526 418294 374582 418350
rect 374154 418170 374210 418226
rect 374278 418170 374334 418226
rect 374402 418170 374458 418226
rect 374526 418170 374582 418226
rect 374154 418046 374210 418102
rect 374278 418046 374334 418102
rect 374402 418046 374458 418102
rect 374526 418046 374582 418102
rect 374154 417922 374210 417978
rect 374278 417922 374334 417978
rect 374402 417922 374458 417978
rect 374526 417922 374582 417978
rect 352716 411542 352772 411598
rect 351036 409742 351092 409798
rect 371878 406294 371934 406350
rect 372002 406294 372058 406350
rect 371878 406170 371934 406226
rect 372002 406170 372058 406226
rect 371878 406046 371934 406102
rect 372002 406046 372058 406102
rect 371878 405922 371934 405978
rect 372002 405922 372058 405978
rect 377874 598116 377930 598172
rect 377998 598116 378054 598172
rect 378122 598116 378178 598172
rect 378246 598116 378302 598172
rect 377874 597992 377930 598048
rect 377998 597992 378054 598048
rect 378122 597992 378178 598048
rect 378246 597992 378302 598048
rect 377874 597868 377930 597924
rect 377998 597868 378054 597924
rect 378122 597868 378178 597924
rect 378246 597868 378302 597924
rect 377874 597744 377930 597800
rect 377998 597744 378054 597800
rect 378122 597744 378178 597800
rect 378246 597744 378302 597800
rect 377874 586294 377930 586350
rect 377998 586294 378054 586350
rect 378122 586294 378178 586350
rect 378246 586294 378302 586350
rect 377874 586170 377930 586226
rect 377998 586170 378054 586226
rect 378122 586170 378178 586226
rect 378246 586170 378302 586226
rect 377874 586046 377930 586102
rect 377998 586046 378054 586102
rect 378122 586046 378178 586102
rect 378246 586046 378302 586102
rect 377874 585922 377930 585978
rect 377998 585922 378054 585978
rect 378122 585922 378178 585978
rect 378246 585922 378302 585978
rect 377874 568294 377930 568350
rect 377998 568294 378054 568350
rect 378122 568294 378178 568350
rect 378246 568294 378302 568350
rect 377874 568170 377930 568226
rect 377998 568170 378054 568226
rect 378122 568170 378178 568226
rect 378246 568170 378302 568226
rect 377874 568046 377930 568102
rect 377998 568046 378054 568102
rect 378122 568046 378178 568102
rect 378246 568046 378302 568102
rect 377874 567922 377930 567978
rect 377998 567922 378054 567978
rect 378122 567922 378178 567978
rect 378246 567922 378302 567978
rect 404874 597156 404930 597212
rect 404998 597156 405054 597212
rect 405122 597156 405178 597212
rect 405246 597156 405302 597212
rect 404874 597032 404930 597088
rect 404998 597032 405054 597088
rect 405122 597032 405178 597088
rect 405246 597032 405302 597088
rect 404874 596908 404930 596964
rect 404998 596908 405054 596964
rect 405122 596908 405178 596964
rect 405246 596908 405302 596964
rect 404874 596784 404930 596840
rect 404998 596784 405054 596840
rect 405122 596784 405178 596840
rect 405246 596784 405302 596840
rect 404874 580294 404930 580350
rect 404998 580294 405054 580350
rect 405122 580294 405178 580350
rect 405246 580294 405302 580350
rect 404874 580170 404930 580226
rect 404998 580170 405054 580226
rect 405122 580170 405178 580226
rect 405246 580170 405302 580226
rect 404874 580046 404930 580102
rect 404998 580046 405054 580102
rect 405122 580046 405178 580102
rect 405246 580046 405302 580102
rect 404874 579922 404930 579978
rect 404998 579922 405054 579978
rect 405122 579922 405178 579978
rect 405246 579922 405302 579978
rect 387238 562294 387294 562350
rect 387362 562294 387418 562350
rect 387238 562170 387294 562226
rect 387362 562170 387418 562226
rect 387238 562046 387294 562102
rect 387362 562046 387418 562102
rect 387238 561922 387294 561978
rect 387362 561922 387418 561978
rect 404874 562294 404930 562350
rect 404998 562294 405054 562350
rect 405122 562294 405178 562350
rect 405246 562294 405302 562350
rect 404874 562170 404930 562226
rect 404998 562170 405054 562226
rect 405122 562170 405178 562226
rect 405246 562170 405302 562226
rect 404874 562046 404930 562102
rect 404998 562046 405054 562102
rect 405122 562046 405178 562102
rect 405246 562046 405302 562102
rect 404874 561922 404930 561978
rect 404998 561922 405054 561978
rect 405122 561922 405178 561978
rect 405246 561922 405302 561978
rect 377874 550294 377930 550350
rect 377998 550294 378054 550350
rect 378122 550294 378178 550350
rect 378246 550294 378302 550350
rect 377874 550170 377930 550226
rect 377998 550170 378054 550226
rect 378122 550170 378178 550226
rect 378246 550170 378302 550226
rect 377874 550046 377930 550102
rect 377998 550046 378054 550102
rect 378122 550046 378178 550102
rect 378246 550046 378302 550102
rect 377874 549922 377930 549978
rect 377998 549922 378054 549978
rect 378122 549922 378178 549978
rect 378246 549922 378302 549978
rect 387238 544294 387294 544350
rect 387362 544294 387418 544350
rect 387238 544170 387294 544226
rect 387362 544170 387418 544226
rect 387238 544046 387294 544102
rect 387362 544046 387418 544102
rect 387238 543922 387294 543978
rect 387362 543922 387418 543978
rect 377874 532294 377930 532350
rect 377998 532294 378054 532350
rect 378122 532294 378178 532350
rect 378246 532294 378302 532350
rect 377874 532170 377930 532226
rect 377998 532170 378054 532226
rect 378122 532170 378178 532226
rect 378246 532170 378302 532226
rect 377874 532046 377930 532102
rect 377998 532046 378054 532102
rect 378122 532046 378178 532102
rect 378246 532046 378302 532102
rect 377874 531922 377930 531978
rect 377998 531922 378054 531978
rect 378122 531922 378178 531978
rect 378246 531922 378302 531978
rect 377874 514294 377930 514350
rect 377998 514294 378054 514350
rect 378122 514294 378178 514350
rect 378246 514294 378302 514350
rect 377874 514170 377930 514226
rect 377998 514170 378054 514226
rect 378122 514170 378178 514226
rect 378246 514170 378302 514226
rect 377874 514046 377930 514102
rect 377998 514046 378054 514102
rect 378122 514046 378178 514102
rect 378246 514046 378302 514102
rect 377874 513922 377930 513978
rect 377998 513922 378054 513978
rect 378122 513922 378178 513978
rect 378246 513922 378302 513978
rect 377874 496294 377930 496350
rect 377998 496294 378054 496350
rect 378122 496294 378178 496350
rect 378246 496294 378302 496350
rect 377874 496170 377930 496226
rect 377998 496170 378054 496226
rect 378122 496170 378178 496226
rect 378246 496170 378302 496226
rect 377874 496046 377930 496102
rect 377998 496046 378054 496102
rect 378122 496046 378178 496102
rect 378246 496046 378302 496102
rect 377874 495922 377930 495978
rect 377998 495922 378054 495978
rect 378122 495922 378178 495978
rect 378246 495922 378302 495978
rect 404874 544294 404930 544350
rect 404998 544294 405054 544350
rect 405122 544294 405178 544350
rect 405246 544294 405302 544350
rect 404874 544170 404930 544226
rect 404998 544170 405054 544226
rect 405122 544170 405178 544226
rect 405246 544170 405302 544226
rect 404874 544046 404930 544102
rect 404998 544046 405054 544102
rect 405122 544046 405178 544102
rect 405246 544046 405302 544102
rect 404874 543922 404930 543978
rect 404998 543922 405054 543978
rect 405122 543922 405178 543978
rect 405246 543922 405302 543978
rect 404874 526294 404930 526350
rect 404998 526294 405054 526350
rect 405122 526294 405178 526350
rect 405246 526294 405302 526350
rect 404874 526170 404930 526226
rect 404998 526170 405054 526226
rect 405122 526170 405178 526226
rect 405246 526170 405302 526226
rect 404874 526046 404930 526102
rect 404998 526046 405054 526102
rect 405122 526046 405178 526102
rect 405246 526046 405302 526102
rect 404874 525922 404930 525978
rect 404998 525922 405054 525978
rect 405122 525922 405178 525978
rect 405246 525922 405302 525978
rect 404874 508294 404930 508350
rect 404998 508294 405054 508350
rect 405122 508294 405178 508350
rect 405246 508294 405302 508350
rect 404874 508170 404930 508226
rect 404998 508170 405054 508226
rect 405122 508170 405178 508226
rect 405246 508170 405302 508226
rect 404874 508046 404930 508102
rect 404998 508046 405054 508102
rect 405122 508046 405178 508102
rect 405246 508046 405302 508102
rect 404874 507922 404930 507978
rect 404998 507922 405054 507978
rect 405122 507922 405178 507978
rect 405246 507922 405302 507978
rect 387238 490294 387294 490350
rect 387362 490294 387418 490350
rect 387238 490170 387294 490226
rect 387362 490170 387418 490226
rect 387238 490046 387294 490102
rect 387362 490046 387418 490102
rect 387238 489922 387294 489978
rect 387362 489922 387418 489978
rect 404874 490294 404930 490350
rect 404998 490294 405054 490350
rect 405122 490294 405178 490350
rect 405246 490294 405302 490350
rect 404874 490170 404930 490226
rect 404998 490170 405054 490226
rect 405122 490170 405178 490226
rect 405246 490170 405302 490226
rect 404874 490046 404930 490102
rect 404998 490046 405054 490102
rect 405122 490046 405178 490102
rect 405246 490046 405302 490102
rect 404874 489922 404930 489978
rect 404998 489922 405054 489978
rect 405122 489922 405178 489978
rect 405246 489922 405302 489978
rect 377874 478294 377930 478350
rect 377998 478294 378054 478350
rect 378122 478294 378178 478350
rect 378246 478294 378302 478350
rect 377874 478170 377930 478226
rect 377998 478170 378054 478226
rect 378122 478170 378178 478226
rect 378246 478170 378302 478226
rect 377874 478046 377930 478102
rect 377998 478046 378054 478102
rect 378122 478046 378178 478102
rect 378246 478046 378302 478102
rect 377874 477922 377930 477978
rect 377998 477922 378054 477978
rect 378122 477922 378178 477978
rect 378246 477922 378302 477978
rect 387238 472294 387294 472350
rect 387362 472294 387418 472350
rect 387238 472170 387294 472226
rect 387362 472170 387418 472226
rect 387238 472046 387294 472102
rect 387362 472046 387418 472102
rect 387238 471922 387294 471978
rect 387362 471922 387418 471978
rect 377874 460294 377930 460350
rect 377998 460294 378054 460350
rect 378122 460294 378178 460350
rect 378246 460294 378302 460350
rect 377874 460170 377930 460226
rect 377998 460170 378054 460226
rect 378122 460170 378178 460226
rect 378246 460170 378302 460226
rect 377874 460046 377930 460102
rect 377998 460046 378054 460102
rect 378122 460046 378178 460102
rect 378246 460046 378302 460102
rect 377874 459922 377930 459978
rect 377998 459922 378054 459978
rect 378122 459922 378178 459978
rect 378246 459922 378302 459978
rect 377874 442294 377930 442350
rect 377998 442294 378054 442350
rect 378122 442294 378178 442350
rect 378246 442294 378302 442350
rect 377874 442170 377930 442226
rect 377998 442170 378054 442226
rect 378122 442170 378178 442226
rect 378246 442170 378302 442226
rect 377874 442046 377930 442102
rect 377998 442046 378054 442102
rect 378122 442046 378178 442102
rect 378246 442046 378302 442102
rect 377874 441922 377930 441978
rect 377998 441922 378054 441978
rect 378122 441922 378178 441978
rect 378246 441922 378302 441978
rect 404874 472294 404930 472350
rect 404998 472294 405054 472350
rect 405122 472294 405178 472350
rect 405246 472294 405302 472350
rect 404874 472170 404930 472226
rect 404998 472170 405054 472226
rect 405122 472170 405178 472226
rect 405246 472170 405302 472226
rect 404874 472046 404930 472102
rect 404998 472046 405054 472102
rect 405122 472046 405178 472102
rect 405246 472046 405302 472102
rect 404874 471922 404930 471978
rect 404998 471922 405054 471978
rect 405122 471922 405178 471978
rect 405246 471922 405302 471978
rect 404874 454294 404930 454350
rect 404998 454294 405054 454350
rect 405122 454294 405178 454350
rect 405246 454294 405302 454350
rect 404874 454170 404930 454226
rect 404998 454170 405054 454226
rect 405122 454170 405178 454226
rect 405246 454170 405302 454226
rect 404874 454046 404930 454102
rect 404998 454046 405054 454102
rect 405122 454046 405178 454102
rect 405246 454046 405302 454102
rect 404874 453922 404930 453978
rect 404998 453922 405054 453978
rect 405122 453922 405178 453978
rect 405246 453922 405302 453978
rect 404874 436294 404930 436350
rect 404998 436294 405054 436350
rect 405122 436294 405178 436350
rect 405246 436294 405302 436350
rect 404874 436170 404930 436226
rect 404998 436170 405054 436226
rect 405122 436170 405178 436226
rect 405246 436170 405302 436226
rect 404874 436046 404930 436102
rect 404998 436046 405054 436102
rect 405122 436046 405178 436102
rect 405246 436046 405302 436102
rect 404874 435922 404930 435978
rect 404998 435922 405054 435978
rect 405122 435922 405178 435978
rect 405246 435922 405302 435978
rect 377874 424294 377930 424350
rect 377998 424294 378054 424350
rect 378122 424294 378178 424350
rect 378246 424294 378302 424350
rect 377874 424170 377930 424226
rect 377998 424170 378054 424226
rect 378122 424170 378178 424226
rect 378246 424170 378302 424226
rect 377874 424046 377930 424102
rect 377998 424046 378054 424102
rect 378122 424046 378178 424102
rect 378246 424046 378302 424102
rect 377874 423922 377930 423978
rect 377998 423922 378054 423978
rect 378122 423922 378178 423978
rect 378246 423922 378302 423978
rect 387238 418294 387294 418350
rect 387362 418294 387418 418350
rect 387238 418170 387294 418226
rect 387362 418170 387418 418226
rect 387238 418046 387294 418102
rect 387362 418046 387418 418102
rect 387238 417922 387294 417978
rect 387362 417922 387418 417978
rect 377874 406294 377930 406350
rect 377998 406294 378054 406350
rect 378122 406294 378178 406350
rect 378246 406294 378302 406350
rect 377874 406170 377930 406226
rect 377998 406170 378054 406226
rect 378122 406170 378178 406226
rect 378246 406170 378302 406226
rect 377874 406046 377930 406102
rect 377998 406046 378054 406102
rect 378122 406046 378178 406102
rect 378246 406046 378302 406102
rect 377874 405922 377930 405978
rect 377998 405922 378054 405978
rect 378122 405922 378178 405978
rect 378246 405922 378302 405978
rect 351036 402362 351092 402418
rect 356518 400294 356574 400350
rect 356642 400294 356698 400350
rect 356518 400170 356574 400226
rect 356642 400170 356698 400226
rect 356518 400046 356574 400102
rect 356642 400046 356698 400102
rect 356518 399922 356574 399978
rect 356642 399922 356698 399978
rect 350364 391382 350420 391438
rect 347154 388294 347210 388350
rect 347278 388294 347334 388350
rect 347402 388294 347458 388350
rect 347526 388294 347582 388350
rect 371836 388333 371892 388389
rect 371940 388333 371996 388389
rect 372044 388333 372100 388389
rect 347154 388170 347210 388226
rect 347278 388170 347334 388226
rect 347402 388170 347458 388226
rect 347526 388170 347582 388226
rect 347154 388046 347210 388102
rect 347278 388046 347334 388102
rect 347402 388046 347458 388102
rect 347526 388046 347582 388102
rect 347154 387922 347210 387978
rect 347278 387922 347334 387978
rect 347402 387922 347458 387978
rect 347526 387922 347582 387978
rect 374154 382294 374210 382350
rect 374278 382294 374334 382350
rect 374402 382294 374458 382350
rect 374526 382294 374582 382350
rect 374154 382170 374210 382226
rect 374278 382170 374334 382226
rect 374402 382170 374458 382226
rect 374526 382170 374582 382226
rect 374154 382046 374210 382102
rect 374278 382046 374334 382102
rect 374402 382046 374458 382102
rect 374526 382046 374582 382102
rect 374154 381922 374210 381978
rect 374278 381922 374334 381978
rect 374402 381922 374458 381978
rect 374526 381922 374582 381978
rect 347154 370294 347210 370350
rect 347278 370294 347334 370350
rect 347402 370294 347458 370350
rect 347526 370294 347582 370350
rect 347154 370170 347210 370226
rect 347278 370170 347334 370226
rect 347402 370170 347458 370226
rect 347526 370170 347582 370226
rect 347154 370046 347210 370102
rect 347278 370046 347334 370102
rect 347402 370046 347458 370102
rect 347526 370046 347582 370102
rect 347154 369922 347210 369978
rect 347278 369922 347334 369978
rect 347402 369922 347458 369978
rect 347526 369922 347582 369978
rect 343434 346294 343490 346350
rect 343558 346294 343614 346350
rect 343682 346294 343738 346350
rect 343806 346294 343862 346350
rect 343434 346170 343490 346226
rect 343558 346170 343614 346226
rect 343682 346170 343738 346226
rect 343806 346170 343862 346226
rect 343434 346046 343490 346102
rect 343558 346046 343614 346102
rect 343682 346046 343738 346102
rect 343806 346046 343862 346102
rect 343434 345922 343490 345978
rect 343558 345922 343614 345978
rect 343682 345922 343738 345978
rect 343806 345922 343862 345978
rect 334460 344402 334516 344458
rect 334348 343502 334404 343558
rect 334460 344222 334516 344278
rect 334348 341342 334404 341398
rect 334460 341522 334516 341578
rect 334460 339722 334516 339778
rect 334460 339362 334516 339418
rect 338604 338642 338660 338698
rect 334348 337922 334404 337978
rect 334460 337742 334516 337798
rect 334460 337562 334516 337618
rect 334348 336122 334404 336178
rect 334460 336302 334516 336358
rect 334460 335942 334516 335998
rect 334460 334682 334516 334738
rect 334460 333602 334516 333658
rect 334460 332522 334516 332578
rect 337708 330902 337764 330958
rect 334460 330722 334516 330778
rect 334460 329282 334516 329338
rect 334460 327482 334516 327538
rect 334460 327302 334516 327358
rect 334460 325862 334516 325918
rect 334460 324062 334516 324118
rect 334348 323882 334404 323938
rect 334460 322442 334516 322498
rect 334460 320822 334516 320878
rect 334460 319022 334516 319078
rect 374154 364294 374210 364350
rect 374278 364294 374334 364350
rect 374402 364294 374458 364350
rect 374526 364294 374582 364350
rect 374154 364170 374210 364226
rect 374278 364170 374334 364226
rect 374402 364170 374458 364226
rect 374526 364170 374582 364226
rect 374154 364046 374210 364102
rect 374278 364046 374334 364102
rect 374402 364046 374458 364102
rect 374526 364046 374582 364102
rect 374154 363922 374210 363978
rect 374278 363922 374334 363978
rect 374402 363922 374458 363978
rect 374526 363922 374582 363978
rect 347154 352294 347210 352350
rect 347278 352294 347334 352350
rect 347402 352294 347458 352350
rect 347526 352294 347582 352350
rect 347154 352170 347210 352226
rect 347278 352170 347334 352226
rect 347402 352170 347458 352226
rect 347526 352170 347582 352226
rect 347154 352046 347210 352102
rect 347278 352046 347334 352102
rect 347402 352046 347458 352102
rect 347526 352046 347582 352102
rect 347154 351922 347210 351978
rect 347278 351922 347334 351978
rect 347402 351922 347458 351978
rect 347526 351922 347582 351978
rect 344428 331982 344484 332038
rect 343434 328294 343490 328350
rect 343558 328294 343614 328350
rect 343682 328294 343738 328350
rect 343806 328294 343862 328350
rect 343434 328170 343490 328226
rect 343558 328170 343614 328226
rect 343682 328170 343738 328226
rect 343806 328170 343862 328226
rect 343434 328046 343490 328102
rect 343558 328046 343614 328102
rect 343682 328046 343738 328102
rect 343806 328046 343862 328102
rect 343434 327922 343490 327978
rect 343558 327922 343614 327978
rect 343682 327922 343738 327978
rect 343806 327922 343862 327978
rect 343434 310294 343490 310350
rect 343558 310294 343614 310350
rect 343682 310294 343738 310350
rect 343806 310294 343862 310350
rect 343434 310170 343490 310226
rect 343558 310170 343614 310226
rect 343682 310170 343738 310226
rect 343806 310170 343862 310226
rect 343434 310046 343490 310102
rect 343558 310046 343614 310102
rect 343682 310046 343738 310102
rect 343806 310046 343862 310102
rect 343434 309922 343490 309978
rect 343558 309922 343614 309978
rect 343682 309922 343738 309978
rect 343806 309922 343862 309978
rect 371878 352294 371934 352350
rect 372002 352294 372058 352350
rect 371878 352170 371934 352226
rect 372002 352170 372058 352226
rect 371878 352046 371934 352102
rect 372002 352046 372058 352102
rect 371878 351922 371934 351978
rect 372002 351922 372058 351978
rect 347154 334294 347210 334350
rect 347278 334294 347334 334350
rect 347402 334294 347458 334350
rect 347526 334294 347582 334350
rect 347154 334170 347210 334226
rect 347278 334170 347334 334226
rect 347402 334170 347458 334226
rect 347526 334170 347582 334226
rect 347154 334046 347210 334102
rect 347278 334046 347334 334102
rect 347402 334046 347458 334102
rect 347526 334046 347582 334102
rect 347154 333922 347210 333978
rect 347278 333922 347334 333978
rect 347402 333922 347458 333978
rect 347526 333922 347582 333978
rect 350252 348722 350308 348778
rect 356518 346294 356574 346350
rect 356642 346294 356698 346350
rect 356518 346170 356574 346226
rect 356642 346170 356698 346226
rect 356518 346046 356574 346102
rect 356642 346046 356698 346102
rect 356518 345922 356574 345978
rect 356642 345922 356698 345978
rect 374154 346294 374210 346350
rect 374278 346294 374334 346350
rect 374402 346294 374458 346350
rect 374526 346294 374582 346350
rect 374154 346170 374210 346226
rect 374278 346170 374334 346226
rect 374402 346170 374458 346226
rect 374526 346170 374582 346226
rect 374154 346046 374210 346102
rect 374278 346046 374334 346102
rect 374402 346046 374458 346102
rect 374526 346046 374582 346102
rect 374154 345922 374210 345978
rect 374278 345922 374334 345978
rect 374402 345922 374458 345978
rect 374526 345922 374582 345978
rect 352716 341162 352772 341218
rect 351148 339542 351204 339598
rect 371878 334294 371934 334350
rect 372002 334294 372058 334350
rect 371878 334170 371934 334226
rect 372002 334170 372058 334226
rect 371878 334046 371934 334102
rect 372002 334046 372058 334102
rect 371878 333922 371934 333978
rect 372002 333922 372058 333978
rect 356518 328294 356574 328350
rect 356642 328294 356698 328350
rect 356518 328170 356574 328226
rect 356642 328170 356698 328226
rect 356518 328046 356574 328102
rect 356642 328046 356698 328102
rect 356518 327922 356574 327978
rect 356642 327922 356698 327978
rect 374154 328294 374210 328350
rect 374278 328294 374334 328350
rect 374402 328294 374458 328350
rect 374526 328294 374582 328350
rect 374154 328170 374210 328226
rect 374278 328170 374334 328226
rect 374402 328170 374458 328226
rect 374526 328170 374582 328226
rect 374154 328046 374210 328102
rect 374278 328046 374334 328102
rect 374402 328046 374458 328102
rect 374526 328046 374582 328102
rect 374154 327922 374210 327978
rect 374278 327922 374334 327978
rect 374402 327922 374458 327978
rect 374526 327922 374582 327978
rect 347154 316294 347210 316350
rect 347278 316294 347334 316350
rect 347402 316294 347458 316350
rect 347526 316294 347582 316350
rect 347154 316170 347210 316226
rect 347278 316170 347334 316226
rect 347402 316170 347458 316226
rect 347526 316170 347582 316226
rect 347154 316046 347210 316102
rect 347278 316046 347334 316102
rect 347402 316046 347458 316102
rect 347526 316046 347582 316102
rect 347154 315922 347210 315978
rect 347278 315922 347334 315978
rect 347402 315922 347458 315978
rect 347526 315922 347582 315978
rect 343434 292294 343490 292350
rect 343558 292294 343614 292350
rect 343682 292294 343738 292350
rect 343806 292294 343862 292350
rect 343434 292170 343490 292226
rect 343558 292170 343614 292226
rect 343682 292170 343738 292226
rect 343806 292170 343862 292226
rect 343434 292046 343490 292102
rect 343558 292046 343614 292102
rect 343682 292046 343738 292102
rect 343806 292046 343862 292102
rect 343434 291922 343490 291978
rect 343558 291922 343614 291978
rect 343682 291922 343738 291978
rect 343806 291922 343862 291978
rect 334348 277982 334404 278038
rect 334460 277262 334516 277318
rect 334460 275642 334516 275698
rect 334460 272942 334516 272998
rect 334348 272222 334404 272278
rect 334460 271502 334516 271558
rect 334572 269702 334628 269758
rect 334460 268802 334516 268858
rect 334348 267362 334404 267418
rect 334460 267902 334516 267958
rect 334460 266462 334516 266518
rect 334572 266282 334628 266338
rect 334460 265382 334516 265438
rect 334460 263762 334516 263818
rect 334460 263582 334516 263638
rect 334460 260702 334516 260758
rect 334460 260540 334516 260578
rect 334460 260522 334516 260540
rect 334460 260342 334516 260398
rect 334460 258916 334516 258958
rect 334460 258902 334516 258916
rect 334460 258542 334516 258598
rect 334460 258182 334516 258238
rect 343434 274294 343490 274350
rect 343558 274294 343614 274350
rect 343682 274294 343738 274350
rect 343806 274294 343862 274350
rect 343434 274170 343490 274226
rect 343558 274170 343614 274226
rect 343682 274170 343738 274226
rect 343806 274170 343862 274226
rect 343434 274046 343490 274102
rect 343558 274046 343614 274102
rect 343682 274046 343738 274102
rect 343806 274046 343862 274102
rect 343434 273922 343490 273978
rect 343558 273922 343614 273978
rect 343682 273922 343738 273978
rect 343806 273922 343862 273978
rect 336924 267002 336980 267058
rect 334684 255302 334740 255358
rect 334460 255122 334516 255178
rect 334348 254942 334404 254998
rect 334460 253502 334516 253558
rect 334460 251882 334516 251938
rect 334348 251702 334404 251758
rect 334460 250082 334516 250138
rect 334460 248462 334516 248518
rect 351932 313982 351988 314038
rect 347154 298294 347210 298350
rect 347278 298294 347334 298350
rect 347402 298294 347458 298350
rect 347526 298294 347582 298350
rect 347154 298170 347210 298226
rect 347278 298170 347334 298226
rect 347402 298170 347458 298226
rect 347526 298170 347582 298226
rect 347154 298046 347210 298102
rect 347278 298046 347334 298102
rect 347402 298046 347458 298102
rect 347526 298046 347582 298102
rect 347154 297922 347210 297978
rect 347278 297922 347334 297978
rect 347402 297922 347458 297978
rect 347526 297922 347582 297978
rect 374154 310294 374210 310350
rect 374278 310294 374334 310350
rect 374402 310294 374458 310350
rect 374526 310294 374582 310350
rect 374154 310170 374210 310226
rect 374278 310170 374334 310226
rect 374402 310170 374458 310226
rect 374526 310170 374582 310226
rect 374154 310046 374210 310102
rect 374278 310046 374334 310102
rect 374402 310046 374458 310102
rect 374526 310046 374582 310102
rect 374154 309922 374210 309978
rect 374278 309922 374334 309978
rect 374402 309922 374458 309978
rect 374526 309922 374582 309978
rect 374154 292294 374210 292350
rect 374278 292294 374334 292350
rect 374402 292294 374458 292350
rect 374526 292294 374582 292350
rect 374154 292170 374210 292226
rect 374278 292170 374334 292226
rect 374402 292170 374458 292226
rect 374526 292170 374582 292226
rect 374154 292046 374210 292102
rect 374278 292046 374334 292102
rect 374402 292046 374458 292102
rect 374526 292046 374582 292102
rect 374154 291922 374210 291978
rect 374278 291922 374334 291978
rect 374402 291922 374458 291978
rect 374526 291922 374582 291978
rect 347154 280294 347210 280350
rect 347278 280294 347334 280350
rect 347402 280294 347458 280350
rect 347526 280294 347582 280350
rect 347154 280170 347210 280226
rect 347278 280170 347334 280226
rect 347402 280170 347458 280226
rect 347526 280170 347582 280226
rect 347154 280046 347210 280102
rect 347278 280046 347334 280102
rect 347402 280046 347458 280102
rect 347526 280046 347582 280102
rect 347154 279922 347210 279978
rect 347278 279922 347334 279978
rect 347402 279922 347458 279978
rect 347526 279922 347582 279978
rect 343434 256294 343490 256350
rect 343558 256294 343614 256350
rect 343682 256294 343738 256350
rect 343806 256294 343862 256350
rect 343434 256170 343490 256226
rect 343558 256170 343614 256226
rect 343682 256170 343738 256226
rect 343806 256170 343862 256226
rect 343434 256046 343490 256102
rect 343558 256046 343614 256102
rect 343682 256046 343738 256102
rect 343806 256046 343862 256102
rect 343434 255922 343490 255978
rect 343558 255922 343614 255978
rect 343682 255922 343738 255978
rect 343806 255922 343862 255978
rect 371878 280294 371934 280350
rect 372002 280294 372058 280350
rect 371878 280170 371934 280226
rect 372002 280170 372058 280226
rect 371878 280046 371934 280102
rect 372002 280046 372058 280102
rect 371878 279922 371934 279978
rect 372002 279922 372058 279978
rect 356518 274294 356574 274350
rect 356642 274294 356698 274350
rect 356518 274170 356574 274226
rect 356642 274170 356698 274226
rect 356518 274046 356574 274102
rect 356642 274046 356698 274102
rect 356518 273922 356574 273978
rect 356642 273922 356698 273978
rect 374154 274294 374210 274350
rect 374278 274294 374334 274350
rect 374402 274294 374458 274350
rect 374526 274294 374582 274350
rect 374154 274170 374210 274226
rect 374278 274170 374334 274226
rect 374402 274170 374458 274226
rect 374526 274170 374582 274226
rect 374154 274046 374210 274102
rect 374278 274046 374334 274102
rect 374402 274046 374458 274102
rect 374526 274046 374582 274102
rect 374154 273922 374210 273978
rect 374278 273922 374334 273978
rect 374402 273922 374458 273978
rect 374526 273922 374582 273978
rect 351036 271682 351092 271738
rect 352716 269522 352772 269578
rect 351932 267182 351988 267238
rect 347788 265202 347844 265258
rect 347154 262294 347210 262350
rect 347278 262294 347334 262350
rect 347402 262294 347458 262350
rect 347526 262294 347582 262350
rect 347154 262170 347210 262226
rect 347278 262170 347334 262226
rect 347402 262170 347458 262226
rect 347526 262170 347582 262226
rect 347154 262046 347210 262102
rect 347278 262046 347334 262102
rect 347402 262046 347458 262102
rect 347526 262046 347582 262102
rect 347154 261922 347210 261978
rect 347278 261922 347334 261978
rect 347402 261922 347458 261978
rect 347526 261922 347582 261978
rect 351036 258722 351092 258778
rect 371878 262294 371934 262350
rect 372002 262294 372058 262350
rect 371878 262170 371934 262226
rect 372002 262170 372058 262226
rect 371878 262046 371934 262102
rect 372002 262046 372058 262102
rect 371878 261922 371934 261978
rect 372002 261922 372058 261978
rect 356518 256294 356574 256350
rect 356642 256294 356698 256350
rect 356518 256170 356574 256226
rect 356642 256170 356698 256226
rect 356518 256046 356574 256102
rect 356642 256046 356698 256102
rect 356518 255922 356574 255978
rect 356642 255922 356698 255978
rect 374154 256294 374210 256350
rect 374278 256294 374334 256350
rect 374402 256294 374458 256350
rect 374526 256294 374582 256350
rect 374154 256170 374210 256226
rect 374278 256170 374334 256226
rect 374402 256170 374458 256226
rect 374526 256170 374582 256226
rect 374154 256046 374210 256102
rect 374278 256046 374334 256102
rect 374402 256046 374458 256102
rect 374526 256046 374582 256102
rect 374154 255922 374210 255978
rect 374278 255922 374334 255978
rect 374402 255922 374458 255978
rect 374526 255922 374582 255978
rect 351036 250262 351092 250318
rect 347154 244294 347210 244350
rect 347278 244294 347334 244350
rect 347402 244294 347458 244350
rect 347526 244294 347582 244350
rect 347154 244170 347210 244226
rect 347278 244170 347334 244226
rect 347402 244170 347458 244226
rect 347526 244170 347582 244226
rect 347154 244046 347210 244102
rect 347278 244046 347334 244102
rect 347402 244046 347458 244102
rect 347526 244046 347582 244102
rect 347154 243922 347210 243978
rect 347278 243922 347334 243978
rect 347402 243922 347458 243978
rect 347526 243922 347582 243978
rect 343434 238294 343490 238350
rect 343558 238294 343614 238350
rect 343682 238294 343738 238350
rect 343806 238294 343862 238350
rect 343434 238170 343490 238226
rect 343558 238170 343614 238226
rect 343682 238170 343738 238226
rect 343806 238170 343862 238226
rect 343434 238046 343490 238102
rect 343558 238046 343614 238102
rect 343682 238046 343738 238102
rect 343806 238046 343862 238102
rect 343434 237922 343490 237978
rect 343558 237922 343614 237978
rect 343682 237922 343738 237978
rect 343806 237922 343862 237978
rect 334460 205082 334516 205138
rect 334460 203282 334516 203338
rect 334460 200762 334516 200818
rect 334460 200042 334516 200098
rect 334460 198242 334516 198298
rect 334460 196802 334516 196858
rect 334460 196622 334516 196678
rect 343434 220294 343490 220350
rect 343558 220294 343614 220350
rect 343682 220294 343738 220350
rect 343806 220294 343862 220350
rect 343434 220170 343490 220226
rect 343558 220170 343614 220226
rect 343682 220170 343738 220226
rect 343806 220170 343862 220226
rect 343434 220046 343490 220102
rect 343558 220046 343614 220102
rect 343682 220046 343738 220102
rect 343806 220046 343862 220102
rect 343434 219922 343490 219978
rect 343558 219922 343614 219978
rect 343682 219922 343738 219978
rect 343806 219922 343862 219978
rect 334460 195002 334516 195058
rect 334460 194822 334516 194878
rect 334460 193922 334516 193978
rect 334460 193202 334516 193258
rect 334460 192302 334516 192358
rect 347154 226294 347210 226350
rect 347278 226294 347334 226350
rect 347402 226294 347458 226350
rect 347526 226294 347582 226350
rect 347154 226170 347210 226226
rect 347278 226170 347334 226226
rect 347402 226170 347458 226226
rect 347526 226170 347582 226226
rect 347154 226046 347210 226102
rect 347278 226046 347334 226102
rect 347402 226046 347458 226102
rect 347526 226046 347582 226102
rect 347154 225922 347210 225978
rect 347278 225922 347334 225978
rect 347402 225922 347458 225978
rect 347526 225922 347582 225978
rect 374154 238294 374210 238350
rect 374278 238294 374334 238350
rect 374402 238294 374458 238350
rect 374526 238294 374582 238350
rect 374154 238170 374210 238226
rect 374278 238170 374334 238226
rect 374402 238170 374458 238226
rect 374526 238170 374582 238226
rect 374154 238046 374210 238102
rect 374278 238046 374334 238102
rect 374402 238046 374458 238102
rect 374526 238046 374582 238102
rect 374154 237922 374210 237978
rect 374278 237922 374334 237978
rect 374402 237922 374458 237978
rect 374526 237922 374582 237978
rect 374154 220294 374210 220350
rect 374278 220294 374334 220350
rect 374402 220294 374458 220350
rect 374526 220294 374582 220350
rect 374154 220170 374210 220226
rect 374278 220170 374334 220226
rect 374402 220170 374458 220226
rect 374526 220170 374582 220226
rect 374154 220046 374210 220102
rect 374278 220046 374334 220102
rect 374402 220046 374458 220102
rect 374526 220046 374582 220102
rect 374154 219922 374210 219978
rect 374278 219922 374334 219978
rect 374402 219922 374458 219978
rect 374526 219922 374582 219978
rect 347154 208294 347210 208350
rect 347278 208294 347334 208350
rect 347402 208294 347458 208350
rect 347526 208294 347582 208350
rect 347154 208170 347210 208226
rect 347278 208170 347334 208226
rect 347402 208170 347458 208226
rect 347526 208170 347582 208226
rect 347154 208046 347210 208102
rect 347278 208046 347334 208102
rect 347402 208046 347458 208102
rect 347526 208046 347582 208102
rect 347154 207922 347210 207978
rect 347278 207922 347334 207978
rect 347402 207922 347458 207978
rect 347526 207922 347582 207978
rect 343434 202294 343490 202350
rect 343558 202294 343614 202350
rect 343682 202294 343738 202350
rect 343806 202294 343862 202350
rect 343434 202170 343490 202226
rect 343558 202170 343614 202226
rect 343682 202170 343738 202226
rect 343806 202170 343862 202226
rect 343434 202046 343490 202102
rect 343558 202046 343614 202102
rect 343682 202046 343738 202102
rect 343806 202046 343862 202102
rect 343434 201922 343490 201978
rect 343558 201922 343614 201978
rect 343682 201922 343738 201978
rect 343806 201922 343862 201978
rect 335132 188882 335188 188938
rect 341852 187982 341908 188038
rect 336028 186362 336084 186418
rect 336140 187262 336196 187318
rect 342636 186182 342692 186238
rect 371878 208294 371934 208350
rect 372002 208294 372058 208350
rect 371878 208170 371934 208226
rect 372002 208170 372058 208226
rect 371878 208046 371934 208102
rect 372002 208046 372058 208102
rect 371878 207922 371934 207978
rect 372002 207922 372058 207978
rect 356518 202294 356574 202350
rect 356642 202294 356698 202350
rect 356518 202170 356574 202226
rect 356642 202170 356698 202226
rect 356518 202046 356574 202102
rect 356642 202046 356698 202102
rect 356518 201922 356574 201978
rect 356642 201922 356698 201978
rect 387238 400294 387294 400350
rect 387362 400294 387418 400350
rect 387238 400170 387294 400226
rect 387362 400170 387418 400226
rect 387238 400046 387294 400102
rect 387362 400046 387418 400102
rect 387238 399922 387294 399978
rect 387362 399922 387418 399978
rect 377874 388294 377930 388350
rect 377998 388294 378054 388350
rect 378122 388294 378178 388350
rect 378246 388294 378302 388350
rect 377874 388170 377930 388226
rect 377998 388170 378054 388226
rect 378122 388170 378178 388226
rect 378246 388170 378302 388226
rect 377874 388046 377930 388102
rect 377998 388046 378054 388102
rect 378122 388046 378178 388102
rect 378246 388046 378302 388102
rect 377874 387922 377930 387978
rect 377998 387922 378054 387978
rect 378122 387922 378178 387978
rect 378246 387922 378302 387978
rect 377874 370294 377930 370350
rect 377998 370294 378054 370350
rect 378122 370294 378178 370350
rect 378246 370294 378302 370350
rect 377874 370170 377930 370226
rect 377998 370170 378054 370226
rect 378122 370170 378178 370226
rect 378246 370170 378302 370226
rect 377874 370046 377930 370102
rect 377998 370046 378054 370102
rect 378122 370046 378178 370102
rect 378246 370046 378302 370102
rect 377874 369922 377930 369978
rect 377998 369922 378054 369978
rect 378122 369922 378178 369978
rect 378246 369922 378302 369978
rect 404874 418294 404930 418350
rect 404998 418294 405054 418350
rect 405122 418294 405178 418350
rect 405246 418294 405302 418350
rect 404874 418170 404930 418226
rect 404998 418170 405054 418226
rect 405122 418170 405178 418226
rect 405246 418170 405302 418226
rect 404874 418046 404930 418102
rect 404998 418046 405054 418102
rect 405122 418046 405178 418102
rect 405246 418046 405302 418102
rect 404874 417922 404930 417978
rect 404998 417922 405054 417978
rect 405122 417922 405178 417978
rect 405246 417922 405302 417978
rect 401436 409922 401492 409978
rect 401436 408122 401492 408178
rect 401212 397862 401268 397918
rect 401436 398942 401492 398998
rect 401324 397322 401380 397378
rect 401436 396242 401492 396298
rect 401324 393002 401380 393058
rect 408594 598116 408650 598172
rect 408718 598116 408774 598172
rect 408842 598116 408898 598172
rect 408966 598116 409022 598172
rect 408594 597992 408650 598048
rect 408718 597992 408774 598048
rect 408842 597992 408898 598048
rect 408966 597992 409022 598048
rect 408594 597868 408650 597924
rect 408718 597868 408774 597924
rect 408842 597868 408898 597924
rect 408966 597868 409022 597924
rect 408594 597744 408650 597800
rect 408718 597744 408774 597800
rect 408842 597744 408898 597800
rect 408966 597744 409022 597800
rect 408594 586294 408650 586350
rect 408718 586294 408774 586350
rect 408842 586294 408898 586350
rect 408966 586294 409022 586350
rect 408594 586170 408650 586226
rect 408718 586170 408774 586226
rect 408842 586170 408898 586226
rect 408966 586170 409022 586226
rect 408594 586046 408650 586102
rect 408718 586046 408774 586102
rect 408842 586046 408898 586102
rect 408966 586046 409022 586102
rect 408594 585922 408650 585978
rect 408718 585922 408774 585978
rect 408842 585922 408898 585978
rect 408966 585922 409022 585978
rect 408594 568294 408650 568350
rect 408718 568294 408774 568350
rect 408842 568294 408898 568350
rect 408966 568294 409022 568350
rect 408594 568170 408650 568226
rect 408718 568170 408774 568226
rect 408842 568170 408898 568226
rect 408966 568170 409022 568226
rect 408594 568046 408650 568102
rect 408718 568046 408774 568102
rect 408842 568046 408898 568102
rect 408966 568046 409022 568102
rect 408594 567922 408650 567978
rect 408718 567922 408774 567978
rect 408842 567922 408898 567978
rect 408966 567922 409022 567978
rect 435594 597156 435650 597212
rect 435718 597156 435774 597212
rect 435842 597156 435898 597212
rect 435966 597156 436022 597212
rect 435594 597032 435650 597088
rect 435718 597032 435774 597088
rect 435842 597032 435898 597088
rect 435966 597032 436022 597088
rect 435594 596908 435650 596964
rect 435718 596908 435774 596964
rect 435842 596908 435898 596964
rect 435966 596908 436022 596964
rect 435594 596784 435650 596840
rect 435718 596784 435774 596840
rect 435842 596784 435898 596840
rect 435966 596784 436022 596840
rect 435594 580294 435650 580350
rect 435718 580294 435774 580350
rect 435842 580294 435898 580350
rect 435966 580294 436022 580350
rect 435594 580170 435650 580226
rect 435718 580170 435774 580226
rect 435842 580170 435898 580226
rect 435966 580170 436022 580226
rect 435594 580046 435650 580102
rect 435718 580046 435774 580102
rect 435842 580046 435898 580102
rect 435966 580046 436022 580102
rect 435594 579922 435650 579978
rect 435718 579922 435774 579978
rect 435842 579922 435898 579978
rect 435966 579922 436022 579978
rect 418518 562294 418574 562350
rect 418642 562294 418698 562350
rect 418518 562170 418574 562226
rect 418642 562170 418698 562226
rect 418518 562046 418574 562102
rect 418642 562046 418698 562102
rect 418518 561922 418574 561978
rect 418642 561922 418698 561978
rect 435594 562294 435650 562350
rect 435718 562294 435774 562350
rect 435842 562294 435898 562350
rect 435966 562294 436022 562350
rect 435594 562170 435650 562226
rect 435718 562170 435774 562226
rect 435842 562170 435898 562226
rect 435966 562170 436022 562226
rect 435594 562046 435650 562102
rect 435718 562046 435774 562102
rect 435842 562046 435898 562102
rect 435966 562046 436022 562102
rect 435594 561922 435650 561978
rect 435718 561922 435774 561978
rect 435842 561922 435898 561978
rect 435966 561922 436022 561978
rect 414652 555182 414708 555238
rect 408594 550294 408650 550350
rect 408718 550294 408774 550350
rect 408842 550294 408898 550350
rect 408966 550294 409022 550350
rect 408594 550170 408650 550226
rect 408718 550170 408774 550226
rect 408842 550170 408898 550226
rect 408966 550170 409022 550226
rect 408594 550046 408650 550102
rect 408718 550046 408774 550102
rect 408842 550046 408898 550102
rect 408966 550046 409022 550102
rect 408594 549922 408650 549978
rect 408718 549922 408774 549978
rect 408842 549922 408898 549978
rect 408966 549922 409022 549978
rect 408594 532294 408650 532350
rect 408718 532294 408774 532350
rect 408842 532294 408898 532350
rect 408966 532294 409022 532350
rect 408594 532170 408650 532226
rect 408718 532170 408774 532226
rect 408842 532170 408898 532226
rect 408966 532170 409022 532226
rect 408594 532046 408650 532102
rect 408718 532046 408774 532102
rect 408842 532046 408898 532102
rect 408966 532046 409022 532102
rect 408594 531922 408650 531978
rect 408718 531922 408774 531978
rect 408842 531922 408898 531978
rect 408966 531922 409022 531978
rect 408594 514294 408650 514350
rect 408718 514294 408774 514350
rect 408842 514294 408898 514350
rect 408966 514294 409022 514350
rect 408594 514170 408650 514226
rect 408718 514170 408774 514226
rect 408842 514170 408898 514226
rect 408966 514170 409022 514226
rect 408594 514046 408650 514102
rect 408718 514046 408774 514102
rect 408842 514046 408898 514102
rect 408966 514046 409022 514102
rect 408594 513922 408650 513978
rect 408718 513922 408774 513978
rect 408842 513922 408898 513978
rect 408966 513922 409022 513978
rect 439314 598116 439370 598172
rect 439438 598116 439494 598172
rect 439562 598116 439618 598172
rect 439686 598116 439742 598172
rect 439314 597992 439370 598048
rect 439438 597992 439494 598048
rect 439562 597992 439618 598048
rect 439686 597992 439742 598048
rect 439314 597868 439370 597924
rect 439438 597868 439494 597924
rect 439562 597868 439618 597924
rect 439686 597868 439742 597924
rect 439314 597744 439370 597800
rect 439438 597744 439494 597800
rect 439562 597744 439618 597800
rect 439686 597744 439742 597800
rect 439314 586294 439370 586350
rect 439438 586294 439494 586350
rect 439562 586294 439618 586350
rect 439686 586294 439742 586350
rect 439314 586170 439370 586226
rect 439438 586170 439494 586226
rect 439562 586170 439618 586226
rect 439686 586170 439742 586226
rect 439314 586046 439370 586102
rect 439438 586046 439494 586102
rect 439562 586046 439618 586102
rect 439686 586046 439742 586102
rect 439314 585922 439370 585978
rect 439438 585922 439494 585978
rect 439562 585922 439618 585978
rect 439686 585922 439742 585978
rect 439314 568294 439370 568350
rect 439438 568294 439494 568350
rect 439562 568294 439618 568350
rect 439686 568294 439742 568350
rect 439314 568170 439370 568226
rect 439438 568170 439494 568226
rect 439562 568170 439618 568226
rect 439686 568170 439742 568226
rect 439314 568046 439370 568102
rect 439438 568046 439494 568102
rect 439562 568046 439618 568102
rect 439686 568046 439742 568102
rect 439314 567922 439370 567978
rect 439438 567922 439494 567978
rect 439562 567922 439618 567978
rect 439686 567922 439742 567978
rect 466314 597156 466370 597212
rect 466438 597156 466494 597212
rect 466562 597156 466618 597212
rect 466686 597156 466742 597212
rect 466314 597032 466370 597088
rect 466438 597032 466494 597088
rect 466562 597032 466618 597088
rect 466686 597032 466742 597088
rect 466314 596908 466370 596964
rect 466438 596908 466494 596964
rect 466562 596908 466618 596964
rect 466686 596908 466742 596964
rect 466314 596784 466370 596840
rect 466438 596784 466494 596840
rect 466562 596784 466618 596840
rect 466686 596784 466742 596840
rect 466314 580294 466370 580350
rect 466438 580294 466494 580350
rect 466562 580294 466618 580350
rect 466686 580294 466742 580350
rect 466314 580170 466370 580226
rect 466438 580170 466494 580226
rect 466562 580170 466618 580226
rect 466686 580170 466742 580226
rect 466314 580046 466370 580102
rect 466438 580046 466494 580102
rect 466562 580046 466618 580102
rect 466686 580046 466742 580102
rect 466314 579922 466370 579978
rect 466438 579922 466494 579978
rect 466562 579922 466618 579978
rect 466686 579922 466742 579978
rect 449238 562294 449294 562350
rect 449362 562294 449418 562350
rect 449238 562170 449294 562226
rect 449362 562170 449418 562226
rect 449238 562046 449294 562102
rect 449362 562046 449418 562102
rect 449238 561922 449294 561978
rect 449362 561922 449418 561978
rect 466314 562294 466370 562350
rect 466438 562294 466494 562350
rect 466562 562294 466618 562350
rect 466686 562294 466742 562350
rect 466314 562170 466370 562226
rect 466438 562170 466494 562226
rect 466562 562170 466618 562226
rect 466686 562170 466742 562226
rect 466314 562046 466370 562102
rect 466438 562046 466494 562102
rect 466562 562046 466618 562102
rect 466686 562046 466742 562102
rect 466314 561922 466370 561978
rect 466438 561922 466494 561978
rect 466562 561922 466618 561978
rect 466686 561922 466742 561978
rect 433878 550294 433934 550350
rect 434002 550294 434058 550350
rect 433878 550170 433934 550226
rect 434002 550170 434058 550226
rect 433878 550046 433934 550102
rect 434002 550046 434058 550102
rect 433878 549922 433934 549978
rect 434002 549922 434058 549978
rect 418518 544294 418574 544350
rect 418642 544294 418698 544350
rect 418518 544170 418574 544226
rect 418642 544170 418698 544226
rect 418518 544046 418574 544102
rect 418642 544046 418698 544102
rect 418518 543922 418574 543978
rect 418642 543922 418698 543978
rect 449238 544294 449294 544350
rect 449362 544294 449418 544350
rect 449238 544170 449294 544226
rect 449362 544170 449418 544226
rect 449238 544046 449294 544102
rect 449362 544046 449418 544102
rect 449238 543922 449294 543978
rect 449362 543922 449418 543978
rect 433878 532294 433934 532350
rect 434002 532294 434058 532350
rect 433878 532170 433934 532226
rect 434002 532170 434058 532226
rect 433878 532046 433934 532102
rect 434002 532046 434058 532102
rect 433878 531922 433934 531978
rect 434002 531922 434058 531978
rect 435594 526294 435650 526350
rect 435718 526294 435774 526350
rect 435842 526294 435898 526350
rect 435966 526294 436022 526350
rect 435594 526170 435650 526226
rect 435718 526170 435774 526226
rect 435842 526170 435898 526226
rect 435966 526170 436022 526226
rect 435594 526046 435650 526102
rect 435718 526046 435774 526102
rect 435842 526046 435898 526102
rect 435966 526046 436022 526102
rect 435594 525922 435650 525978
rect 435718 525922 435774 525978
rect 435842 525922 435898 525978
rect 435966 525922 436022 525978
rect 435594 508294 435650 508350
rect 435718 508294 435774 508350
rect 435842 508294 435898 508350
rect 435966 508294 436022 508350
rect 435594 508170 435650 508226
rect 435718 508170 435774 508226
rect 435842 508170 435898 508226
rect 435966 508170 436022 508226
rect 435594 508046 435650 508102
rect 435718 508046 435774 508102
rect 435842 508046 435898 508102
rect 435966 508046 436022 508102
rect 435594 507922 435650 507978
rect 435718 507922 435774 507978
rect 435842 507922 435898 507978
rect 435966 507922 436022 507978
rect 408594 496294 408650 496350
rect 408718 496294 408774 496350
rect 408842 496294 408898 496350
rect 408966 496294 409022 496350
rect 408594 496170 408650 496226
rect 408718 496170 408774 496226
rect 408842 496170 408898 496226
rect 408966 496170 409022 496226
rect 408594 496046 408650 496102
rect 408718 496046 408774 496102
rect 408842 496046 408898 496102
rect 408966 496046 409022 496102
rect 408594 495922 408650 495978
rect 408718 495922 408774 495978
rect 408842 495922 408898 495978
rect 408966 495922 409022 495978
rect 418518 490294 418574 490350
rect 418642 490294 418698 490350
rect 418518 490170 418574 490226
rect 418642 490170 418698 490226
rect 418518 490046 418574 490102
rect 418642 490046 418698 490102
rect 418518 489922 418574 489978
rect 418642 489922 418698 489978
rect 435594 490294 435650 490350
rect 435718 490294 435774 490350
rect 435842 490294 435898 490350
rect 435966 490294 436022 490350
rect 435594 490170 435650 490226
rect 435718 490170 435774 490226
rect 435842 490170 435898 490226
rect 435966 490170 436022 490226
rect 435594 490046 435650 490102
rect 435718 490046 435774 490102
rect 435842 490046 435898 490102
rect 435966 490046 436022 490102
rect 435594 489922 435650 489978
rect 435718 489922 435774 489978
rect 435842 489922 435898 489978
rect 435966 489922 436022 489978
rect 414652 483902 414708 483958
rect 408594 478294 408650 478350
rect 408718 478294 408774 478350
rect 408842 478294 408898 478350
rect 408966 478294 409022 478350
rect 408594 478170 408650 478226
rect 408718 478170 408774 478226
rect 408842 478170 408898 478226
rect 408966 478170 409022 478226
rect 408594 478046 408650 478102
rect 408718 478046 408774 478102
rect 408842 478046 408898 478102
rect 408966 478046 409022 478102
rect 408594 477922 408650 477978
rect 408718 477922 408774 477978
rect 408842 477922 408898 477978
rect 408966 477922 409022 477978
rect 408594 460294 408650 460350
rect 408718 460294 408774 460350
rect 408842 460294 408898 460350
rect 408966 460294 409022 460350
rect 408594 460170 408650 460226
rect 408718 460170 408774 460226
rect 408842 460170 408898 460226
rect 408966 460170 409022 460226
rect 408594 460046 408650 460102
rect 408718 460046 408774 460102
rect 408842 460046 408898 460102
rect 408966 460046 409022 460102
rect 408594 459922 408650 459978
rect 408718 459922 408774 459978
rect 408842 459922 408898 459978
rect 408966 459922 409022 459978
rect 433878 478294 433934 478350
rect 434002 478294 434058 478350
rect 433878 478170 433934 478226
rect 434002 478170 434058 478226
rect 433878 478046 433934 478102
rect 434002 478046 434058 478102
rect 439314 532294 439370 532350
rect 439438 532294 439494 532350
rect 439562 532294 439618 532350
rect 439686 532294 439742 532350
rect 439314 532170 439370 532226
rect 439438 532170 439494 532226
rect 439562 532170 439618 532226
rect 439686 532170 439742 532226
rect 439314 532046 439370 532102
rect 439438 532046 439494 532102
rect 439562 532046 439618 532102
rect 439686 532046 439742 532102
rect 439314 531922 439370 531978
rect 439438 531922 439494 531978
rect 439562 531922 439618 531978
rect 439686 531922 439742 531978
rect 439314 514294 439370 514350
rect 439438 514294 439494 514350
rect 439562 514294 439618 514350
rect 439686 514294 439742 514350
rect 439314 514170 439370 514226
rect 439438 514170 439494 514226
rect 439562 514170 439618 514226
rect 439686 514170 439742 514226
rect 439314 514046 439370 514102
rect 439438 514046 439494 514102
rect 439562 514046 439618 514102
rect 439686 514046 439742 514102
rect 439314 513922 439370 513978
rect 439438 513922 439494 513978
rect 439562 513922 439618 513978
rect 439686 513922 439742 513978
rect 466314 544294 466370 544350
rect 466438 544294 466494 544350
rect 466562 544294 466618 544350
rect 466686 544294 466742 544350
rect 466314 544170 466370 544226
rect 466438 544170 466494 544226
rect 466562 544170 466618 544226
rect 466686 544170 466742 544226
rect 466314 544046 466370 544102
rect 466438 544046 466494 544102
rect 466562 544046 466618 544102
rect 466686 544046 466742 544102
rect 466314 543922 466370 543978
rect 466438 543922 466494 543978
rect 466562 543922 466618 543978
rect 466686 543922 466742 543978
rect 466314 526294 466370 526350
rect 466438 526294 466494 526350
rect 466562 526294 466618 526350
rect 466686 526294 466742 526350
rect 466314 526170 466370 526226
rect 466438 526170 466494 526226
rect 466562 526170 466618 526226
rect 466686 526170 466742 526226
rect 466314 526046 466370 526102
rect 466438 526046 466494 526102
rect 466562 526046 466618 526102
rect 466686 526046 466742 526102
rect 466314 525922 466370 525978
rect 466438 525922 466494 525978
rect 466562 525922 466618 525978
rect 466686 525922 466742 525978
rect 466314 508294 466370 508350
rect 466438 508294 466494 508350
rect 466562 508294 466618 508350
rect 466686 508294 466742 508350
rect 466314 508170 466370 508226
rect 466438 508170 466494 508226
rect 466562 508170 466618 508226
rect 466686 508170 466742 508226
rect 466314 508046 466370 508102
rect 466438 508046 466494 508102
rect 466562 508046 466618 508102
rect 466686 508046 466742 508102
rect 466314 507922 466370 507978
rect 466438 507922 466494 507978
rect 466562 507922 466618 507978
rect 466686 507922 466742 507978
rect 439314 496294 439370 496350
rect 439438 496294 439494 496350
rect 439562 496294 439618 496350
rect 439686 496294 439742 496350
rect 439314 496170 439370 496226
rect 439438 496170 439494 496226
rect 439562 496170 439618 496226
rect 439686 496170 439742 496226
rect 439314 496046 439370 496102
rect 439438 496046 439494 496102
rect 439562 496046 439618 496102
rect 439686 496046 439742 496102
rect 439314 495922 439370 495978
rect 439438 495922 439494 495978
rect 439562 495922 439618 495978
rect 439686 495922 439742 495978
rect 449238 490294 449294 490350
rect 449362 490294 449418 490350
rect 449238 490170 449294 490226
rect 449362 490170 449418 490226
rect 449238 490046 449294 490102
rect 449362 490046 449418 490102
rect 449238 489922 449294 489978
rect 449362 489922 449418 489978
rect 439314 478294 439370 478350
rect 439438 478294 439494 478350
rect 439562 478294 439618 478350
rect 439686 478294 439742 478350
rect 439314 478170 439370 478226
rect 439438 478170 439494 478226
rect 439562 478170 439618 478226
rect 439686 478170 439742 478226
rect 433878 477922 433934 477978
rect 434002 477922 434058 477978
rect 439314 478046 439370 478102
rect 439438 478046 439494 478102
rect 439562 478046 439618 478102
rect 439686 478046 439742 478102
rect 439314 477922 439370 477978
rect 439438 477922 439494 477978
rect 439562 477922 439618 477978
rect 439686 477922 439742 477978
rect 418518 472294 418574 472350
rect 418642 472294 418698 472350
rect 418518 472170 418574 472226
rect 418642 472170 418698 472226
rect 418518 472046 418574 472102
rect 418642 472046 418698 472102
rect 418518 471922 418574 471978
rect 418642 471922 418698 471978
rect 435594 472004 435650 472060
rect 435718 472004 435774 472060
rect 435842 472004 435898 472060
rect 435966 472004 436022 472060
rect 435594 471880 435650 471936
rect 435718 471880 435774 471936
rect 435842 471880 435898 471936
rect 435966 471880 436022 471936
rect 433878 460294 433934 460350
rect 434002 460294 434058 460350
rect 433878 460170 433934 460226
rect 434002 460170 434058 460226
rect 433878 460046 433934 460102
rect 434002 460046 434058 460102
rect 433878 459922 433934 459978
rect 434002 459922 434058 459978
rect 435594 454294 435650 454350
rect 435718 454294 435774 454350
rect 435842 454294 435898 454350
rect 435966 454294 436022 454350
rect 435594 454170 435650 454226
rect 435718 454170 435774 454226
rect 435842 454170 435898 454226
rect 435966 454170 436022 454226
rect 435594 454046 435650 454102
rect 435718 454046 435774 454102
rect 435842 454046 435898 454102
rect 435966 454046 436022 454102
rect 435594 453922 435650 453978
rect 435718 453922 435774 453978
rect 435842 453922 435898 453978
rect 435966 453922 436022 453978
rect 408594 442294 408650 442350
rect 408718 442294 408774 442350
rect 408842 442294 408898 442350
rect 408966 442294 409022 442350
rect 408594 442170 408650 442226
rect 408718 442170 408774 442226
rect 408842 442170 408898 442226
rect 408966 442170 409022 442226
rect 408594 442046 408650 442102
rect 408718 442046 408774 442102
rect 408842 442046 408898 442102
rect 408966 442046 409022 442102
rect 408594 441922 408650 441978
rect 408718 441922 408774 441978
rect 408842 441922 408898 441978
rect 408966 441922 409022 441978
rect 408594 424294 408650 424350
rect 408718 424294 408774 424350
rect 408842 424294 408898 424350
rect 408966 424294 409022 424350
rect 408594 424170 408650 424226
rect 408718 424170 408774 424226
rect 408842 424170 408898 424226
rect 408966 424170 409022 424226
rect 408594 424046 408650 424102
rect 408718 424046 408774 424102
rect 408842 424046 408898 424102
rect 408966 424046 409022 424102
rect 408594 423922 408650 423978
rect 408718 423922 408774 423978
rect 408842 423922 408898 423978
rect 408966 423922 409022 423978
rect 435594 436294 435650 436350
rect 435718 436294 435774 436350
rect 435842 436294 435898 436350
rect 435966 436294 436022 436350
rect 435594 436170 435650 436226
rect 435718 436170 435774 436226
rect 435842 436170 435898 436226
rect 435966 436170 436022 436226
rect 435594 436046 435650 436102
rect 435718 436046 435774 436102
rect 435842 436046 435898 436102
rect 435966 436046 436022 436102
rect 435594 435922 435650 435978
rect 435718 435922 435774 435978
rect 435842 435922 435898 435978
rect 435966 435922 436022 435978
rect 408594 406294 408650 406350
rect 408718 406294 408774 406350
rect 408842 406294 408898 406350
rect 408966 406294 409022 406350
rect 408594 406170 408650 406226
rect 408718 406170 408774 406226
rect 408842 406170 408898 406226
rect 408966 406170 409022 406226
rect 404874 400294 404930 400350
rect 404998 400294 405054 400350
rect 405122 400294 405178 400350
rect 405246 400294 405302 400350
rect 404874 400170 404930 400226
rect 404998 400170 405054 400226
rect 405122 400170 405178 400226
rect 405246 400170 405302 400226
rect 404874 400046 404930 400102
rect 404998 400046 405054 400102
rect 405122 400046 405178 400102
rect 405246 400046 405302 400102
rect 404874 399922 404930 399978
rect 404998 399922 405054 399978
rect 405122 399922 405178 399978
rect 405246 399922 405302 399978
rect 406588 399662 406644 399718
rect 408594 406046 408650 406102
rect 408718 406046 408774 406102
rect 408842 406046 408898 406102
rect 408966 406046 409022 406102
rect 408594 405922 408650 405978
rect 408718 405922 408774 405978
rect 408842 405922 408898 405978
rect 408966 405922 409022 405978
rect 404874 382294 404930 382350
rect 404998 382294 405054 382350
rect 405122 382294 405178 382350
rect 405246 382294 405302 382350
rect 404874 382170 404930 382226
rect 404998 382170 405054 382226
rect 405122 382170 405178 382226
rect 405246 382170 405302 382226
rect 404874 382046 404930 382102
rect 404998 382046 405054 382102
rect 405122 382046 405178 382102
rect 405246 382046 405302 382102
rect 404874 381922 404930 381978
rect 404998 381922 405054 381978
rect 405122 381922 405178 381978
rect 405246 381922 405302 381978
rect 404874 364294 404930 364350
rect 404998 364294 405054 364350
rect 405122 364294 405178 364350
rect 405246 364294 405302 364350
rect 404874 364170 404930 364226
rect 404998 364170 405054 364226
rect 405122 364170 405178 364226
rect 405246 364170 405302 364226
rect 404874 364046 404930 364102
rect 404998 364046 405054 364102
rect 405122 364046 405178 364102
rect 405246 364046 405302 364102
rect 404874 363922 404930 363978
rect 404998 363922 405054 363978
rect 405122 363922 405178 363978
rect 405246 363922 405302 363978
rect 377874 352294 377930 352350
rect 377998 352294 378054 352350
rect 378122 352294 378178 352350
rect 378246 352294 378302 352350
rect 377874 352170 377930 352226
rect 377998 352170 378054 352226
rect 378122 352170 378178 352226
rect 378246 352170 378302 352226
rect 377874 352046 377930 352102
rect 377998 352046 378054 352102
rect 378122 352046 378178 352102
rect 378246 352046 378302 352102
rect 377874 351922 377930 351978
rect 377998 351922 378054 351978
rect 378122 351922 378178 351978
rect 378246 351922 378302 351978
rect 393372 349262 393428 349318
rect 394828 348542 394884 348598
rect 387238 346294 387294 346350
rect 387362 346294 387418 346350
rect 387238 346170 387294 346226
rect 387362 346170 387418 346226
rect 387238 346046 387294 346102
rect 387362 346046 387418 346102
rect 387238 345922 387294 345978
rect 387362 345922 387418 345978
rect 394828 344222 394884 344278
rect 404874 346294 404930 346350
rect 404998 346294 405054 346350
rect 405122 346294 405178 346350
rect 405246 346294 405302 346350
rect 404874 346170 404930 346226
rect 404998 346170 405054 346226
rect 405122 346170 405178 346226
rect 405246 346170 405302 346226
rect 404874 346046 404930 346102
rect 404998 346046 405054 346102
rect 405122 346046 405178 346102
rect 405246 346046 405302 346102
rect 404874 345922 404930 345978
rect 404998 345922 405054 345978
rect 405122 345922 405178 345978
rect 405246 345922 405302 345978
rect 393372 339182 393428 339238
rect 377874 334294 377930 334350
rect 377998 334294 378054 334350
rect 378122 334294 378178 334350
rect 378246 334294 378302 334350
rect 377874 334170 377930 334226
rect 377998 334170 378054 334226
rect 378122 334170 378178 334226
rect 378246 334170 378302 334226
rect 377874 334046 377930 334102
rect 377998 334046 378054 334102
rect 378122 334046 378178 334102
rect 378246 334046 378302 334102
rect 377874 333922 377930 333978
rect 377998 333922 378054 333978
rect 378122 333922 378178 333978
rect 378246 333922 378302 333978
rect 393148 336302 393204 336358
rect 393484 333602 393540 333658
rect 393372 332522 393428 332578
rect 393148 331802 393204 331858
rect 393260 329462 393316 329518
rect 387238 328294 387294 328350
rect 387362 328294 387418 328350
rect 387238 328170 387294 328226
rect 387362 328170 387418 328226
rect 387238 328046 387294 328102
rect 387362 328046 387418 328102
rect 387238 327922 387294 327978
rect 387362 327922 387418 327978
rect 377874 316294 377930 316350
rect 377998 316294 378054 316350
rect 378122 316294 378178 316350
rect 378246 316294 378302 316350
rect 377874 316170 377930 316226
rect 377998 316170 378054 316226
rect 378122 316170 378178 316226
rect 378246 316170 378302 316226
rect 377874 316046 377930 316102
rect 377998 316046 378054 316102
rect 378122 316046 378178 316102
rect 378246 316046 378302 316102
rect 377874 315922 377930 315978
rect 377998 315922 378054 315978
rect 378122 315922 378178 315978
rect 378246 315922 378302 315978
rect 404460 339722 404516 339778
rect 394828 338462 394884 338518
rect 394828 337562 394884 337618
rect 396508 337922 396564 337978
rect 396508 336842 396564 336898
rect 394828 332522 394884 332578
rect 394940 330722 394996 330778
rect 394828 327482 394884 327538
rect 394044 327302 394100 327358
rect 399756 336122 399812 336178
rect 404572 337742 404628 337798
rect 404572 335942 404628 335998
rect 404460 335042 404516 335098
rect 403228 334682 403284 334738
rect 403228 330002 403284 330058
rect 418518 418294 418574 418350
rect 418642 418294 418698 418350
rect 418518 418170 418574 418226
rect 418642 418170 418698 418226
rect 418518 418046 418574 418102
rect 418642 418046 418698 418102
rect 418518 417922 418574 417978
rect 418642 417922 418698 417978
rect 449238 472294 449294 472350
rect 449362 472294 449418 472350
rect 449238 472170 449294 472226
rect 449362 472170 449418 472226
rect 449238 472046 449294 472102
rect 449362 472046 449418 472102
rect 449238 471922 449294 471978
rect 449362 471922 449418 471978
rect 439314 460294 439370 460350
rect 439438 460294 439494 460350
rect 439562 460294 439618 460350
rect 439686 460294 439742 460350
rect 439314 460170 439370 460226
rect 439438 460170 439494 460226
rect 439562 460170 439618 460226
rect 439686 460170 439742 460226
rect 439314 460046 439370 460102
rect 439438 460046 439494 460102
rect 439562 460046 439618 460102
rect 439686 460046 439742 460102
rect 439314 459922 439370 459978
rect 439438 459922 439494 459978
rect 439562 459922 439618 459978
rect 439686 459922 439742 459978
rect 439314 442294 439370 442350
rect 439438 442294 439494 442350
rect 439562 442294 439618 442350
rect 439686 442294 439742 442350
rect 439314 442170 439370 442226
rect 439438 442170 439494 442226
rect 439562 442170 439618 442226
rect 439686 442170 439742 442226
rect 439314 442046 439370 442102
rect 439438 442046 439494 442102
rect 439562 442046 439618 442102
rect 439686 442046 439742 442102
rect 439314 441922 439370 441978
rect 439438 441922 439494 441978
rect 439562 441922 439618 441978
rect 439686 441922 439742 441978
rect 435594 418294 435650 418350
rect 435718 418294 435774 418350
rect 435842 418294 435898 418350
rect 435966 418294 436022 418350
rect 435594 418170 435650 418226
rect 435718 418170 435774 418226
rect 435842 418170 435898 418226
rect 435966 418170 436022 418226
rect 435594 418046 435650 418102
rect 435718 418046 435774 418102
rect 435842 418046 435898 418102
rect 435966 418046 436022 418102
rect 435594 417922 435650 417978
rect 435718 417922 435774 417978
rect 435842 417922 435898 417978
rect 435966 417922 436022 417978
rect 414092 413702 414148 413758
rect 411516 411542 411572 411598
rect 411180 406682 411236 406738
rect 411068 402362 411124 402418
rect 414652 413342 414708 413398
rect 428876 412082 428932 412138
rect 466314 490294 466370 490350
rect 466438 490294 466494 490350
rect 466562 490294 466618 490350
rect 466686 490294 466742 490350
rect 466314 490170 466370 490226
rect 466438 490170 466494 490226
rect 466562 490170 466618 490226
rect 466686 490170 466742 490226
rect 466314 490046 466370 490102
rect 466438 490046 466494 490102
rect 466562 490046 466618 490102
rect 466686 490046 466742 490102
rect 466314 489922 466370 489978
rect 466438 489922 466494 489978
rect 466562 489922 466618 489978
rect 466686 489922 466742 489978
rect 462812 462842 462868 462898
rect 470034 598116 470090 598172
rect 470158 598116 470214 598172
rect 470282 598116 470338 598172
rect 470406 598116 470462 598172
rect 470034 597992 470090 598048
rect 470158 597992 470214 598048
rect 470282 597992 470338 598048
rect 470406 597992 470462 598048
rect 470034 597868 470090 597924
rect 470158 597868 470214 597924
rect 470282 597868 470338 597924
rect 470406 597868 470462 597924
rect 470034 597744 470090 597800
rect 470158 597744 470214 597800
rect 470282 597744 470338 597800
rect 470406 597744 470462 597800
rect 470034 586294 470090 586350
rect 470158 586294 470214 586350
rect 470282 586294 470338 586350
rect 470406 586294 470462 586350
rect 470034 586170 470090 586226
rect 470158 586170 470214 586226
rect 470282 586170 470338 586226
rect 470406 586170 470462 586226
rect 470034 586046 470090 586102
rect 470158 586046 470214 586102
rect 470282 586046 470338 586102
rect 470406 586046 470462 586102
rect 470034 585922 470090 585978
rect 470158 585922 470214 585978
rect 470282 585922 470338 585978
rect 470406 585922 470462 585978
rect 470034 568294 470090 568350
rect 470158 568294 470214 568350
rect 470282 568294 470338 568350
rect 470406 568294 470462 568350
rect 470034 568170 470090 568226
rect 470158 568170 470214 568226
rect 470282 568170 470338 568226
rect 470406 568170 470462 568226
rect 470034 568046 470090 568102
rect 470158 568046 470214 568102
rect 470282 568046 470338 568102
rect 470406 568046 470462 568102
rect 470034 567922 470090 567978
rect 470158 567922 470214 567978
rect 470282 567922 470338 567978
rect 470406 567922 470462 567978
rect 497034 597156 497090 597212
rect 497158 597156 497214 597212
rect 497282 597156 497338 597212
rect 497406 597156 497462 597212
rect 497034 597032 497090 597088
rect 497158 597032 497214 597088
rect 497282 597032 497338 597088
rect 497406 597032 497462 597088
rect 497034 596908 497090 596964
rect 497158 596908 497214 596964
rect 497282 596908 497338 596964
rect 497406 596908 497462 596964
rect 497034 596784 497090 596840
rect 497158 596784 497214 596840
rect 497282 596784 497338 596840
rect 497406 596784 497462 596840
rect 497034 580294 497090 580350
rect 497158 580294 497214 580350
rect 497282 580294 497338 580350
rect 497406 580294 497462 580350
rect 497034 580170 497090 580226
rect 497158 580170 497214 580226
rect 497282 580170 497338 580226
rect 497406 580170 497462 580226
rect 497034 580046 497090 580102
rect 497158 580046 497214 580102
rect 497282 580046 497338 580102
rect 497406 580046 497462 580102
rect 497034 579922 497090 579978
rect 497158 579922 497214 579978
rect 497282 579922 497338 579978
rect 497406 579922 497462 579978
rect 480518 562294 480574 562350
rect 480642 562294 480698 562350
rect 480518 562170 480574 562226
rect 480642 562170 480698 562226
rect 480518 562046 480574 562102
rect 480642 562046 480698 562102
rect 480518 561922 480574 561978
rect 480642 561922 480698 561978
rect 497034 562294 497090 562350
rect 497158 562294 497214 562350
rect 497282 562294 497338 562350
rect 497406 562294 497462 562350
rect 497034 562170 497090 562226
rect 497158 562170 497214 562226
rect 497282 562170 497338 562226
rect 497406 562170 497462 562226
rect 497034 562046 497090 562102
rect 497158 562046 497214 562102
rect 497282 562046 497338 562102
rect 497406 562046 497462 562102
rect 497034 561922 497090 561978
rect 497158 561922 497214 561978
rect 497282 561922 497338 561978
rect 497406 561922 497462 561978
rect 500754 598116 500810 598172
rect 500878 598116 500934 598172
rect 501002 598116 501058 598172
rect 501126 598116 501182 598172
rect 500754 597992 500810 598048
rect 500878 597992 500934 598048
rect 501002 597992 501058 598048
rect 501126 597992 501182 598048
rect 500754 597868 500810 597924
rect 500878 597868 500934 597924
rect 501002 597868 501058 597924
rect 501126 597868 501182 597924
rect 500754 597744 500810 597800
rect 500878 597744 500934 597800
rect 501002 597744 501058 597800
rect 501126 597744 501182 597800
rect 500754 586294 500810 586350
rect 500878 586294 500934 586350
rect 501002 586294 501058 586350
rect 501126 586294 501182 586350
rect 500754 586170 500810 586226
rect 500878 586170 500934 586226
rect 501002 586170 501058 586226
rect 501126 586170 501182 586226
rect 500754 586046 500810 586102
rect 500878 586046 500934 586102
rect 501002 586046 501058 586102
rect 501126 586046 501182 586102
rect 500754 585922 500810 585978
rect 500878 585922 500934 585978
rect 501002 585922 501058 585978
rect 501126 585922 501182 585978
rect 500754 568294 500810 568350
rect 500878 568294 500934 568350
rect 501002 568294 501058 568350
rect 501126 568294 501182 568350
rect 500754 568170 500810 568226
rect 500878 568170 500934 568226
rect 501002 568170 501058 568226
rect 501126 568170 501182 568226
rect 500754 568046 500810 568102
rect 500878 568046 500934 568102
rect 501002 568046 501058 568102
rect 501126 568046 501182 568102
rect 500754 567922 500810 567978
rect 500878 567922 500934 567978
rect 501002 567922 501058 567978
rect 501126 567922 501182 567978
rect 527754 597156 527810 597212
rect 527878 597156 527934 597212
rect 528002 597156 528058 597212
rect 528126 597156 528182 597212
rect 527754 597032 527810 597088
rect 527878 597032 527934 597088
rect 528002 597032 528058 597088
rect 528126 597032 528182 597088
rect 527754 596908 527810 596964
rect 527878 596908 527934 596964
rect 528002 596908 528058 596964
rect 528126 596908 528182 596964
rect 527754 596784 527810 596840
rect 527878 596784 527934 596840
rect 528002 596784 528058 596840
rect 528126 596784 528182 596840
rect 527754 580294 527810 580350
rect 527878 580294 527934 580350
rect 528002 580294 528058 580350
rect 528126 580294 528182 580350
rect 527754 580170 527810 580226
rect 527878 580170 527934 580226
rect 528002 580170 528058 580226
rect 528126 580170 528182 580226
rect 527754 580046 527810 580102
rect 527878 580046 527934 580102
rect 528002 580046 528058 580102
rect 528126 580046 528182 580102
rect 527754 579922 527810 579978
rect 527878 579922 527934 579978
rect 528002 579922 528058 579978
rect 528126 579922 528182 579978
rect 511238 562294 511294 562350
rect 511362 562294 511418 562350
rect 511238 562170 511294 562226
rect 511362 562170 511418 562226
rect 511238 562046 511294 562102
rect 511362 562046 511418 562102
rect 511238 561922 511294 561978
rect 511362 561922 511418 561978
rect 527754 562294 527810 562350
rect 527878 562294 527934 562350
rect 528002 562294 528058 562350
rect 528126 562294 528182 562350
rect 527754 562170 527810 562226
rect 527878 562170 527934 562226
rect 528002 562170 528058 562226
rect 528126 562170 528182 562226
rect 527754 562046 527810 562102
rect 527878 562046 527934 562102
rect 528002 562046 528058 562102
rect 528126 562046 528182 562102
rect 527754 561922 527810 561978
rect 527878 561922 527934 561978
rect 528002 561922 528058 561978
rect 528126 561922 528182 561978
rect 473676 555212 473732 555238
rect 473676 555182 473732 555212
rect 476028 554642 476084 554698
rect 519036 554462 519092 554518
rect 470034 550294 470090 550350
rect 470158 550294 470214 550350
rect 470282 550294 470338 550350
rect 470406 550294 470462 550350
rect 470034 550170 470090 550226
rect 470158 550170 470214 550226
rect 470282 550170 470338 550226
rect 470406 550170 470462 550226
rect 470034 550046 470090 550102
rect 470158 550046 470214 550102
rect 470282 550046 470338 550102
rect 470406 550046 470462 550102
rect 470034 549922 470090 549978
rect 470158 549922 470214 549978
rect 470282 549922 470338 549978
rect 470406 549922 470462 549978
rect 470034 532294 470090 532350
rect 470158 532294 470214 532350
rect 470282 532294 470338 532350
rect 470406 532294 470462 532350
rect 470034 532170 470090 532226
rect 470158 532170 470214 532226
rect 470282 532170 470338 532226
rect 470406 532170 470462 532226
rect 470034 532046 470090 532102
rect 470158 532046 470214 532102
rect 470282 532046 470338 532102
rect 470406 532046 470462 532102
rect 470034 531922 470090 531978
rect 470158 531922 470214 531978
rect 470282 531922 470338 531978
rect 470406 531922 470462 531978
rect 470034 514294 470090 514350
rect 470158 514294 470214 514350
rect 470282 514294 470338 514350
rect 470406 514294 470462 514350
rect 470034 514170 470090 514226
rect 470158 514170 470214 514226
rect 470282 514170 470338 514226
rect 470406 514170 470462 514226
rect 470034 514046 470090 514102
rect 470158 514046 470214 514102
rect 470282 514046 470338 514102
rect 470406 514046 470462 514102
rect 470034 513922 470090 513978
rect 470158 513922 470214 513978
rect 470282 513922 470338 513978
rect 470406 513922 470462 513978
rect 495878 550294 495934 550350
rect 496002 550294 496058 550350
rect 495878 550170 495934 550226
rect 496002 550170 496058 550226
rect 495878 550046 495934 550102
rect 496002 550046 496058 550102
rect 495878 549922 495934 549978
rect 496002 549922 496058 549978
rect 480518 544294 480574 544350
rect 480642 544294 480698 544350
rect 480518 544170 480574 544226
rect 480642 544170 480698 544226
rect 480518 544046 480574 544102
rect 480642 544046 480698 544102
rect 480518 543922 480574 543978
rect 480642 543922 480698 543978
rect 497034 544294 497090 544350
rect 497158 544294 497214 544350
rect 497282 544294 497338 544350
rect 497406 544294 497462 544350
rect 497034 544170 497090 544226
rect 497158 544170 497214 544226
rect 497282 544170 497338 544226
rect 497406 544170 497462 544226
rect 497034 544046 497090 544102
rect 497158 544046 497214 544102
rect 497282 544046 497338 544102
rect 497406 544046 497462 544102
rect 497034 543922 497090 543978
rect 497158 543922 497214 543978
rect 497282 543922 497338 543978
rect 497406 543922 497462 543978
rect 495878 532294 495934 532350
rect 496002 532294 496058 532350
rect 495878 532170 495934 532226
rect 496002 532170 496058 532226
rect 495878 532046 495934 532102
rect 496002 532046 496058 532102
rect 495878 531922 495934 531978
rect 496002 531922 496058 531978
rect 497034 526294 497090 526350
rect 497158 526294 497214 526350
rect 497282 526294 497338 526350
rect 497406 526294 497462 526350
rect 497034 526170 497090 526226
rect 497158 526170 497214 526226
rect 497282 526170 497338 526226
rect 497406 526170 497462 526226
rect 497034 526046 497090 526102
rect 497158 526046 497214 526102
rect 497282 526046 497338 526102
rect 497406 526046 497462 526102
rect 497034 525922 497090 525978
rect 497158 525922 497214 525978
rect 497282 525922 497338 525978
rect 497406 525922 497462 525978
rect 497034 508294 497090 508350
rect 497158 508294 497214 508350
rect 497282 508294 497338 508350
rect 497406 508294 497462 508350
rect 497034 508170 497090 508226
rect 497158 508170 497214 508226
rect 497282 508170 497338 508226
rect 497406 508170 497462 508226
rect 497034 508046 497090 508102
rect 497158 508046 497214 508102
rect 497282 508046 497338 508102
rect 497406 508046 497462 508102
rect 497034 507922 497090 507978
rect 497158 507922 497214 507978
rect 497282 507922 497338 507978
rect 497406 507922 497462 507978
rect 470034 496294 470090 496350
rect 470158 496294 470214 496350
rect 470282 496294 470338 496350
rect 470406 496294 470462 496350
rect 470034 496170 470090 496226
rect 470158 496170 470214 496226
rect 470282 496170 470338 496226
rect 470406 496170 470462 496226
rect 470034 496046 470090 496102
rect 470158 496046 470214 496102
rect 470282 496046 470338 496102
rect 470406 496046 470462 496102
rect 470034 495922 470090 495978
rect 470158 495922 470214 495978
rect 470282 495922 470338 495978
rect 470406 495922 470462 495978
rect 480518 490294 480574 490350
rect 480642 490294 480698 490350
rect 480518 490170 480574 490226
rect 480642 490170 480698 490226
rect 480518 490046 480574 490102
rect 480642 490046 480698 490102
rect 480518 489922 480574 489978
rect 480642 489922 480698 489978
rect 497034 490294 497090 490350
rect 497158 490294 497214 490350
rect 497282 490294 497338 490350
rect 497406 490294 497462 490350
rect 497034 490170 497090 490226
rect 497158 490170 497214 490226
rect 497282 490170 497338 490226
rect 497406 490170 497462 490226
rect 497034 490046 497090 490102
rect 497158 490046 497214 490102
rect 497282 490046 497338 490102
rect 497406 490046 497462 490102
rect 497034 489922 497090 489978
rect 497158 489922 497214 489978
rect 497282 489922 497338 489978
rect 497406 489922 497462 489978
rect 476028 484622 476084 484678
rect 473676 483902 473732 483958
rect 472220 480482 472276 480538
rect 470034 478294 470090 478350
rect 470158 478294 470214 478350
rect 470282 478294 470338 478350
rect 470406 478294 470462 478350
rect 470034 478170 470090 478226
rect 470158 478170 470214 478226
rect 470282 478170 470338 478226
rect 470406 478170 470462 478226
rect 470034 478046 470090 478102
rect 470158 478046 470214 478102
rect 470282 478046 470338 478102
rect 470406 478046 470462 478102
rect 466314 472294 466370 472350
rect 466438 472294 466494 472350
rect 466562 472294 466618 472350
rect 466686 472294 466742 472350
rect 466314 472170 466370 472226
rect 466438 472170 466494 472226
rect 466562 472170 466618 472226
rect 466686 472170 466742 472226
rect 466314 472046 466370 472102
rect 466438 472046 466494 472102
rect 466562 472046 466618 472102
rect 466686 472046 466742 472102
rect 466314 471922 466370 471978
rect 466438 471922 466494 471978
rect 466562 471922 466618 471978
rect 466686 471922 466742 471978
rect 466314 454294 466370 454350
rect 466438 454294 466494 454350
rect 466562 454294 466618 454350
rect 466686 454294 466742 454350
rect 466314 454170 466370 454226
rect 466438 454170 466494 454226
rect 466562 454170 466618 454226
rect 466686 454170 466742 454226
rect 466314 454046 466370 454102
rect 466438 454046 466494 454102
rect 466562 454046 466618 454102
rect 466686 454046 466742 454102
rect 466314 453922 466370 453978
rect 466438 453922 466494 453978
rect 466562 453922 466618 453978
rect 466686 453922 466742 453978
rect 466314 436294 466370 436350
rect 466438 436294 466494 436350
rect 466562 436294 466618 436350
rect 466686 436294 466742 436350
rect 466314 436170 466370 436226
rect 466438 436170 466494 436226
rect 466562 436170 466618 436226
rect 466686 436170 466742 436226
rect 466314 436046 466370 436102
rect 466438 436046 466494 436102
rect 466562 436046 466618 436102
rect 466686 436046 466742 436102
rect 466314 435922 466370 435978
rect 466438 435922 466494 435978
rect 466562 435922 466618 435978
rect 466686 435922 466742 435978
rect 439314 424294 439370 424350
rect 439438 424294 439494 424350
rect 439562 424294 439618 424350
rect 439686 424294 439742 424350
rect 439314 424170 439370 424226
rect 439438 424170 439494 424226
rect 439562 424170 439618 424226
rect 439686 424170 439742 424226
rect 439314 424046 439370 424102
rect 439438 424046 439494 424102
rect 439562 424046 439618 424102
rect 439686 424046 439742 424102
rect 439314 423922 439370 423978
rect 439438 423922 439494 423978
rect 439562 423922 439618 423978
rect 439686 423922 439742 423978
rect 449238 418294 449294 418350
rect 449362 418294 449418 418350
rect 449238 418170 449294 418226
rect 449362 418170 449418 418226
rect 449238 418046 449294 418102
rect 449362 418046 449418 418102
rect 449238 417922 449294 417978
rect 449362 417922 449418 417978
rect 470034 477922 470090 477978
rect 470158 477922 470214 477978
rect 470282 477922 470338 477978
rect 470406 477922 470462 477978
rect 470034 460294 470090 460350
rect 470158 460294 470214 460350
rect 470282 460294 470338 460350
rect 470406 460294 470462 460350
rect 470034 460170 470090 460226
rect 470158 460170 470214 460226
rect 470282 460170 470338 460226
rect 470406 460170 470462 460226
rect 470034 460046 470090 460102
rect 470158 460046 470214 460102
rect 470282 460046 470338 460102
rect 470406 460046 470462 460102
rect 470034 459922 470090 459978
rect 470158 459922 470214 459978
rect 470282 459922 470338 459978
rect 470406 459922 470462 459978
rect 495878 478294 495934 478350
rect 496002 478294 496058 478350
rect 495878 478170 495934 478226
rect 496002 478170 496058 478226
rect 495878 478046 495934 478102
rect 496002 478046 496058 478102
rect 495878 477922 495934 477978
rect 496002 477922 496058 477978
rect 500754 550294 500810 550350
rect 500878 550294 500934 550350
rect 501002 550294 501058 550350
rect 501126 550294 501182 550350
rect 500754 550170 500810 550226
rect 500878 550170 500934 550226
rect 501002 550170 501058 550226
rect 501126 550170 501182 550226
rect 500754 550046 500810 550102
rect 500878 550046 500934 550102
rect 501002 550046 501058 550102
rect 501126 550046 501182 550102
rect 500754 549922 500810 549978
rect 500878 549922 500934 549978
rect 501002 549922 501058 549978
rect 501126 549922 501182 549978
rect 511238 544294 511294 544350
rect 511362 544294 511418 544350
rect 511238 544170 511294 544226
rect 511362 544170 511418 544226
rect 511238 544046 511294 544102
rect 511362 544046 511418 544102
rect 511238 543922 511294 543978
rect 511362 543922 511418 543978
rect 500754 532294 500810 532350
rect 500878 532294 500934 532350
rect 501002 532294 501058 532350
rect 501126 532294 501182 532350
rect 500754 532170 500810 532226
rect 500878 532170 500934 532226
rect 501002 532170 501058 532226
rect 501126 532170 501182 532226
rect 500754 532046 500810 532102
rect 500878 532046 500934 532102
rect 501002 532046 501058 532102
rect 501126 532046 501182 532102
rect 500754 531922 500810 531978
rect 500878 531922 500934 531978
rect 501002 531922 501058 531978
rect 501126 531922 501182 531978
rect 500754 514294 500810 514350
rect 500878 514294 500934 514350
rect 501002 514294 501058 514350
rect 501126 514294 501182 514350
rect 500754 514170 500810 514226
rect 500878 514170 500934 514226
rect 501002 514170 501058 514226
rect 501126 514170 501182 514226
rect 500754 514046 500810 514102
rect 500878 514046 500934 514102
rect 501002 514046 501058 514102
rect 501126 514046 501182 514102
rect 500754 513922 500810 513978
rect 500878 513922 500934 513978
rect 501002 513922 501058 513978
rect 501126 513922 501182 513978
rect 527754 544294 527810 544350
rect 527878 544294 527934 544350
rect 528002 544294 528058 544350
rect 528126 544294 528182 544350
rect 527754 544170 527810 544226
rect 527878 544170 527934 544226
rect 528002 544170 528058 544226
rect 528126 544170 528182 544226
rect 527754 544046 527810 544102
rect 527878 544046 527934 544102
rect 528002 544046 528058 544102
rect 528126 544046 528182 544102
rect 527754 543922 527810 543978
rect 527878 543922 527934 543978
rect 528002 543922 528058 543978
rect 528126 543922 528182 543978
rect 527754 526294 527810 526350
rect 527878 526294 527934 526350
rect 528002 526294 528058 526350
rect 528126 526294 528182 526350
rect 527754 526170 527810 526226
rect 527878 526170 527934 526226
rect 528002 526170 528058 526226
rect 528126 526170 528182 526226
rect 527754 526046 527810 526102
rect 527878 526046 527934 526102
rect 528002 526046 528058 526102
rect 528126 526046 528182 526102
rect 527754 525922 527810 525978
rect 527878 525922 527934 525978
rect 528002 525922 528058 525978
rect 528126 525922 528182 525978
rect 527754 508294 527810 508350
rect 527878 508294 527934 508350
rect 528002 508294 528058 508350
rect 528126 508294 528182 508350
rect 527754 508170 527810 508226
rect 527878 508170 527934 508226
rect 528002 508170 528058 508226
rect 528126 508170 528182 508226
rect 527754 508046 527810 508102
rect 527878 508046 527934 508102
rect 528002 508046 528058 508102
rect 528126 508046 528182 508102
rect 527754 507922 527810 507978
rect 527878 507922 527934 507978
rect 528002 507922 528058 507978
rect 528126 507922 528182 507978
rect 500754 496294 500810 496350
rect 500878 496294 500934 496350
rect 501002 496294 501058 496350
rect 501126 496294 501182 496350
rect 500754 496170 500810 496226
rect 500878 496170 500934 496226
rect 501002 496170 501058 496226
rect 501126 496170 501182 496226
rect 500754 496046 500810 496102
rect 500878 496046 500934 496102
rect 501002 496046 501058 496102
rect 501126 496046 501182 496102
rect 500754 495922 500810 495978
rect 500878 495922 500934 495978
rect 501002 495922 501058 495978
rect 501126 495922 501182 495978
rect 511238 490294 511294 490350
rect 511362 490294 511418 490350
rect 511238 490170 511294 490226
rect 511362 490170 511418 490226
rect 511238 490046 511294 490102
rect 511362 490046 511418 490102
rect 511238 489922 511294 489978
rect 511362 489922 511418 489978
rect 527754 490294 527810 490350
rect 527878 490294 527934 490350
rect 528002 490294 528058 490350
rect 528126 490294 528182 490350
rect 527754 490170 527810 490226
rect 527878 490170 527934 490226
rect 528002 490170 528058 490226
rect 528126 490170 528182 490226
rect 527754 490046 527810 490102
rect 527878 490046 527934 490102
rect 528002 490046 528058 490102
rect 528126 490046 528182 490102
rect 527754 489922 527810 489978
rect 527878 489922 527934 489978
rect 528002 489922 528058 489978
rect 528126 489922 528182 489978
rect 500754 478294 500810 478350
rect 500878 478294 500934 478350
rect 501002 478294 501058 478350
rect 501126 478294 501182 478350
rect 500754 478170 500810 478226
rect 500878 478170 500934 478226
rect 501002 478170 501058 478226
rect 501126 478170 501182 478226
rect 500754 478046 500810 478102
rect 500878 478046 500934 478102
rect 501002 478046 501058 478102
rect 501126 478046 501182 478102
rect 500754 477922 500810 477978
rect 500878 477922 500934 477978
rect 501002 477922 501058 477978
rect 501126 477922 501182 477978
rect 480518 472294 480574 472350
rect 480642 472294 480698 472350
rect 480518 472170 480574 472226
rect 480642 472170 480698 472226
rect 480518 472046 480574 472102
rect 480642 472046 480698 472102
rect 480518 471922 480574 471978
rect 480642 471922 480698 471978
rect 473116 465182 473172 465238
rect 495878 460294 495934 460350
rect 496002 460294 496058 460350
rect 495878 460170 495934 460226
rect 496002 460170 496058 460226
rect 495878 460046 495934 460102
rect 496002 460046 496058 460102
rect 495878 459922 495934 459978
rect 496002 459922 496058 459978
rect 497034 454294 497090 454350
rect 497158 454294 497214 454350
rect 497282 454294 497338 454350
rect 497406 454294 497462 454350
rect 497034 454170 497090 454226
rect 497158 454170 497214 454226
rect 497282 454170 497338 454226
rect 497406 454170 497462 454226
rect 497034 454046 497090 454102
rect 497158 454046 497214 454102
rect 497282 454046 497338 454102
rect 497406 454046 497462 454102
rect 497034 453922 497090 453978
rect 497158 453922 497214 453978
rect 497282 453922 497338 453978
rect 497406 453922 497462 453978
rect 470034 442294 470090 442350
rect 470158 442294 470214 442350
rect 470282 442294 470338 442350
rect 470406 442294 470462 442350
rect 470034 442170 470090 442226
rect 470158 442170 470214 442226
rect 470282 442170 470338 442226
rect 470406 442170 470462 442226
rect 470034 442046 470090 442102
rect 470158 442046 470214 442102
rect 470282 442046 470338 442102
rect 470406 442046 470462 442102
rect 470034 441922 470090 441978
rect 470158 441922 470214 441978
rect 470282 441922 470338 441978
rect 470406 441922 470462 441978
rect 466314 418294 466370 418350
rect 466438 418294 466494 418350
rect 466562 418294 466618 418350
rect 466686 418294 466742 418350
rect 466314 418170 466370 418226
rect 466438 418170 466494 418226
rect 466562 418170 466618 418226
rect 466686 418170 466742 418226
rect 466314 418046 466370 418102
rect 466438 418046 466494 418102
rect 466562 418046 466618 418102
rect 466686 418046 466742 418102
rect 466314 417922 466370 417978
rect 466438 417922 466494 417978
rect 466562 417922 466618 417978
rect 466686 417922 466742 417978
rect 440972 411902 441028 411958
rect 428876 407402 428932 407458
rect 440972 407402 441028 407458
rect 433878 406294 433934 406350
rect 434002 406294 434058 406350
rect 433878 406170 433934 406226
rect 434002 406170 434058 406226
rect 433878 406046 433934 406102
rect 434002 406046 434058 406102
rect 433878 405922 433934 405978
rect 434002 405922 434058 405978
rect 414092 402902 414148 402958
rect 418518 400294 418574 400350
rect 418642 400294 418698 400350
rect 418518 400170 418574 400226
rect 418642 400170 418698 400226
rect 418518 400046 418574 400102
rect 418642 400046 418698 400102
rect 418518 399922 418574 399978
rect 418642 399922 418698 399978
rect 435594 400294 435650 400350
rect 435718 400294 435774 400350
rect 435842 400294 435898 400350
rect 435966 400294 436022 400350
rect 435594 400170 435650 400226
rect 435718 400170 435774 400226
rect 435842 400170 435898 400226
rect 435966 400170 436022 400226
rect 435594 400046 435650 400102
rect 435718 400046 435774 400102
rect 435842 400046 435898 400102
rect 435966 400046 436022 400102
rect 435594 399922 435650 399978
rect 435718 399922 435774 399978
rect 435842 399922 435898 399978
rect 435966 399922 436022 399978
rect 411180 398042 411236 398098
rect 410732 394442 410788 394498
rect 408594 388294 408650 388350
rect 408718 388294 408774 388350
rect 408842 388294 408898 388350
rect 408966 388294 409022 388350
rect 433836 388333 433892 388389
rect 433940 388333 433996 388389
rect 434044 388333 434100 388389
rect 408594 388170 408650 388226
rect 408718 388170 408774 388226
rect 408842 388170 408898 388226
rect 408966 388170 409022 388226
rect 408594 388046 408650 388102
rect 408718 388046 408774 388102
rect 408842 388046 408898 388102
rect 408966 388046 409022 388102
rect 408594 387922 408650 387978
rect 408718 387922 408774 387978
rect 408842 387922 408898 387978
rect 408966 387922 409022 387978
rect 408594 370294 408650 370350
rect 408718 370294 408774 370350
rect 408842 370294 408898 370350
rect 408966 370294 409022 370350
rect 408594 370170 408650 370226
rect 408718 370170 408774 370226
rect 408842 370170 408898 370226
rect 408966 370170 409022 370226
rect 408594 370046 408650 370102
rect 408718 370046 408774 370102
rect 408842 370046 408898 370102
rect 408966 370046 409022 370102
rect 408594 369922 408650 369978
rect 408718 369922 408774 369978
rect 408842 369922 408898 369978
rect 408966 369922 409022 369978
rect 435594 382294 435650 382350
rect 435718 382294 435774 382350
rect 435842 382294 435898 382350
rect 435966 382294 436022 382350
rect 435594 382170 435650 382226
rect 435718 382170 435774 382226
rect 435842 382170 435898 382226
rect 435966 382170 436022 382226
rect 435594 382046 435650 382102
rect 435718 382046 435774 382102
rect 435842 382046 435898 382102
rect 435966 382046 436022 382102
rect 435594 381922 435650 381978
rect 435718 381922 435774 381978
rect 435842 381922 435898 381978
rect 435966 381922 436022 381978
rect 435594 364294 435650 364350
rect 435718 364294 435774 364350
rect 435842 364294 435898 364350
rect 435966 364294 436022 364350
rect 435594 364170 435650 364226
rect 435718 364170 435774 364226
rect 435842 364170 435898 364226
rect 435966 364170 436022 364226
rect 435594 364046 435650 364102
rect 435718 364046 435774 364102
rect 435842 364046 435898 364102
rect 435966 364046 436022 364102
rect 435594 363922 435650 363978
rect 435718 363922 435774 363978
rect 435842 363922 435898 363978
rect 435966 363922 436022 363978
rect 408594 352294 408650 352350
rect 408718 352294 408774 352350
rect 408842 352294 408898 352350
rect 408966 352294 409022 352350
rect 408594 352170 408650 352226
rect 408718 352170 408774 352226
rect 408842 352170 408898 352226
rect 408966 352170 409022 352226
rect 408594 352046 408650 352102
rect 408718 352046 408774 352102
rect 408842 352046 408898 352102
rect 408966 352046 409022 352102
rect 408594 351922 408650 351978
rect 408718 351922 408774 351978
rect 408842 351922 408898 351978
rect 408966 351922 409022 351978
rect 407372 341522 407428 341578
rect 433878 352294 433934 352350
rect 434002 352294 434058 352350
rect 433878 352170 433934 352226
rect 434002 352170 434058 352226
rect 433878 352046 433934 352102
rect 434002 352046 434058 352102
rect 433878 351922 433934 351978
rect 434002 351922 434058 351978
rect 418518 346294 418574 346350
rect 418642 346294 418698 346350
rect 418518 346170 418574 346226
rect 418642 346170 418698 346226
rect 418518 346046 418574 346102
rect 418642 346046 418698 346102
rect 418518 345922 418574 345978
rect 418642 345922 418698 345978
rect 435594 346294 435650 346350
rect 435718 346294 435774 346350
rect 435842 346294 435898 346350
rect 435966 346294 436022 346350
rect 435594 346170 435650 346226
rect 435718 346170 435774 346226
rect 435842 346170 435898 346226
rect 435966 346170 436022 346226
rect 435594 346046 435650 346102
rect 435718 346046 435774 346102
rect 435842 346046 435898 346102
rect 435966 346046 436022 346102
rect 435594 345922 435650 345978
rect 435718 345922 435774 345978
rect 435842 345922 435898 345978
rect 435966 345922 436022 345978
rect 414652 341162 414708 341218
rect 408594 334294 408650 334350
rect 408718 334294 408774 334350
rect 408842 334294 408898 334350
rect 408966 334294 409022 334350
rect 408594 334170 408650 334226
rect 408718 334170 408774 334226
rect 408842 334170 408898 334226
rect 408966 334170 409022 334226
rect 408594 334046 408650 334102
rect 408718 334046 408774 334102
rect 408842 334046 408898 334102
rect 408966 334046 409022 334102
rect 408594 333922 408650 333978
rect 408718 333922 408774 333978
rect 408842 333922 408898 333978
rect 408966 333922 409022 333978
rect 404874 328294 404930 328350
rect 404998 328294 405054 328350
rect 405122 328294 405178 328350
rect 405246 328294 405302 328350
rect 404874 328170 404930 328226
rect 404998 328170 405054 328226
rect 405122 328170 405178 328226
rect 405246 328170 405302 328226
rect 404874 328046 404930 328102
rect 404998 328046 405054 328102
rect 405122 328046 405178 328102
rect 405246 328046 405302 328102
rect 404874 327922 404930 327978
rect 404998 327922 405054 327978
rect 405122 327922 405178 327978
rect 405246 327922 405302 327978
rect 404572 326762 404628 326818
rect 404572 320822 404628 320878
rect 404874 310294 404930 310350
rect 404998 310294 405054 310350
rect 405122 310294 405178 310350
rect 405246 310294 405302 310350
rect 404874 310170 404930 310226
rect 404998 310170 405054 310226
rect 405122 310170 405178 310226
rect 405246 310170 405302 310226
rect 404874 310046 404930 310102
rect 404998 310046 405054 310102
rect 405122 310046 405178 310102
rect 405246 310046 405302 310102
rect 404874 309922 404930 309978
rect 404998 309922 405054 309978
rect 405122 309922 405178 309978
rect 405246 309922 405302 309978
rect 377874 298294 377930 298350
rect 377998 298294 378054 298350
rect 378122 298294 378178 298350
rect 378246 298294 378302 298350
rect 377874 298170 377930 298226
rect 377998 298170 378054 298226
rect 378122 298170 378178 298226
rect 378246 298170 378302 298226
rect 377874 298046 377930 298102
rect 377998 298046 378054 298102
rect 378122 298046 378178 298102
rect 378246 298046 378302 298102
rect 377874 297922 377930 297978
rect 377998 297922 378054 297978
rect 378122 297922 378178 297978
rect 378246 297922 378302 297978
rect 377874 280294 377930 280350
rect 377998 280294 378054 280350
rect 378122 280294 378178 280350
rect 378246 280294 378302 280350
rect 377874 280170 377930 280226
rect 377998 280170 378054 280226
rect 378122 280170 378178 280226
rect 378246 280170 378302 280226
rect 377874 280046 377930 280102
rect 377998 280046 378054 280102
rect 378122 280046 378178 280102
rect 378246 280046 378302 280102
rect 377874 279922 377930 279978
rect 377998 279922 378054 279978
rect 378122 279922 378178 279978
rect 378246 279922 378302 279978
rect 404874 292294 404930 292350
rect 404998 292294 405054 292350
rect 405122 292294 405178 292350
rect 405246 292294 405302 292350
rect 404874 292170 404930 292226
rect 404998 292170 405054 292226
rect 405122 292170 405178 292226
rect 405246 292170 405302 292226
rect 404874 292046 404930 292102
rect 404998 292046 405054 292102
rect 405122 292046 405178 292102
rect 405246 292046 405302 292102
rect 404874 291922 404930 291978
rect 404998 291922 405054 291978
rect 405122 291922 405178 291978
rect 405246 291922 405302 291978
rect 394828 275642 394884 275698
rect 387238 274294 387294 274350
rect 387362 274294 387418 274350
rect 387238 274170 387294 274226
rect 387362 274170 387418 274226
rect 387238 274046 387294 274102
rect 387362 274046 387418 274102
rect 387238 273922 387294 273978
rect 387362 273922 387418 273978
rect 404874 274294 404930 274350
rect 404998 274294 405054 274350
rect 405122 274294 405178 274350
rect 405246 274294 405302 274350
rect 404874 274170 404930 274226
rect 404998 274170 405054 274226
rect 405122 274170 405178 274226
rect 405246 274170 405302 274226
rect 404874 274046 404930 274102
rect 404998 274046 405054 274102
rect 405122 274046 405178 274102
rect 405246 274046 405302 274102
rect 404874 273922 404930 273978
rect 404998 273922 405054 273978
rect 405122 273922 405178 273978
rect 405246 273922 405302 273978
rect 396620 272942 396676 272998
rect 394828 271322 394884 271378
rect 395612 272222 395668 272278
rect 394828 269702 394884 269758
rect 393820 268982 393876 269038
rect 393484 268802 393540 268858
rect 377874 262294 377930 262350
rect 377998 262294 378054 262350
rect 378122 262294 378178 262350
rect 378246 262294 378302 262350
rect 377874 262170 377930 262226
rect 377998 262170 378054 262226
rect 378122 262170 378178 262226
rect 378246 262170 378302 262226
rect 377874 262046 377930 262102
rect 377998 262046 378054 262102
rect 378122 262046 378178 262102
rect 378246 262046 378302 262102
rect 377874 261922 377930 261978
rect 377998 261922 378054 261978
rect 378122 261922 378178 261978
rect 378246 261922 378302 261978
rect 393260 267362 393316 267418
rect 393372 266642 393428 266698
rect 393372 264852 393428 264898
rect 393372 264842 393428 264852
rect 393596 266642 393652 266698
rect 393596 263582 393652 263638
rect 393820 260342 393876 260398
rect 393148 258902 393204 258958
rect 393148 258362 393204 258418
rect 387238 256294 387294 256350
rect 387362 256294 387418 256350
rect 387238 256170 387294 256226
rect 387362 256170 387418 256226
rect 387238 256046 387294 256102
rect 387362 256046 387418 256102
rect 387238 255922 387294 255978
rect 387362 255922 387418 255978
rect 377874 244294 377930 244350
rect 377998 244294 378054 244350
rect 378122 244294 378178 244350
rect 378246 244294 378302 244350
rect 377874 244170 377930 244226
rect 377998 244170 378054 244226
rect 378122 244170 378178 244226
rect 378246 244170 378302 244226
rect 377874 244046 377930 244102
rect 377998 244046 378054 244102
rect 378122 244046 378178 244102
rect 378246 244046 378302 244102
rect 377874 243922 377930 243978
rect 377998 243922 378054 243978
rect 378122 243922 378178 243978
rect 378246 243922 378302 243978
rect 396844 271682 396900 271738
rect 396956 271502 397012 271558
rect 398972 254942 399028 254998
rect 404012 250082 404068 250138
rect 433878 334294 433934 334350
rect 434002 334294 434058 334350
rect 433878 334170 433934 334226
rect 434002 334170 434058 334226
rect 433878 334046 433934 334102
rect 434002 334046 434058 334102
rect 433878 333922 433934 333978
rect 434002 333922 434058 333978
rect 418518 328294 418574 328350
rect 418642 328294 418698 328350
rect 418518 328170 418574 328226
rect 418642 328170 418698 328226
rect 418518 328046 418574 328102
rect 418642 328046 418698 328102
rect 418518 327922 418574 327978
rect 418642 327922 418698 327978
rect 435594 328294 435650 328350
rect 435718 328294 435774 328350
rect 435842 328294 435898 328350
rect 435966 328294 436022 328350
rect 435594 328170 435650 328226
rect 435718 328170 435774 328226
rect 435842 328170 435898 328226
rect 435966 328170 436022 328226
rect 435594 328046 435650 328102
rect 435718 328046 435774 328102
rect 435842 328046 435898 328102
rect 435966 328046 436022 328102
rect 435594 327922 435650 327978
rect 435718 327922 435774 327978
rect 435842 327922 435898 327978
rect 435966 327922 436022 327978
rect 408594 316294 408650 316350
rect 408718 316294 408774 316350
rect 408842 316294 408898 316350
rect 408966 316294 409022 316350
rect 408594 316170 408650 316226
rect 408718 316170 408774 316226
rect 408842 316170 408898 316226
rect 408966 316170 409022 316226
rect 408594 316046 408650 316102
rect 408718 316046 408774 316102
rect 408842 316046 408898 316102
rect 408966 316046 409022 316102
rect 408594 315922 408650 315978
rect 408718 315922 408774 315978
rect 408842 315922 408898 315978
rect 408966 315922 409022 315978
rect 408594 298294 408650 298350
rect 408718 298294 408774 298350
rect 408842 298294 408898 298350
rect 408966 298294 409022 298350
rect 408594 298170 408650 298226
rect 408718 298170 408774 298226
rect 408842 298170 408898 298226
rect 408966 298170 409022 298226
rect 408594 298046 408650 298102
rect 408718 298046 408774 298102
rect 408842 298046 408898 298102
rect 408966 298046 409022 298102
rect 408594 297922 408650 297978
rect 408718 297922 408774 297978
rect 408842 297922 408898 297978
rect 408966 297922 409022 297978
rect 435594 310294 435650 310350
rect 435718 310294 435774 310350
rect 435842 310294 435898 310350
rect 435966 310294 436022 310350
rect 435594 310170 435650 310226
rect 435718 310170 435774 310226
rect 435842 310170 435898 310226
rect 435966 310170 436022 310226
rect 435594 310046 435650 310102
rect 435718 310046 435774 310102
rect 435842 310046 435898 310102
rect 435966 310046 436022 310102
rect 435594 309922 435650 309978
rect 435718 309922 435774 309978
rect 435842 309922 435898 309978
rect 435966 309922 436022 309978
rect 435594 292294 435650 292350
rect 435718 292294 435774 292350
rect 435842 292294 435898 292350
rect 435966 292294 436022 292350
rect 435594 292170 435650 292226
rect 435718 292170 435774 292226
rect 435842 292170 435898 292226
rect 435966 292170 436022 292226
rect 435594 292046 435650 292102
rect 435718 292046 435774 292102
rect 435842 292046 435898 292102
rect 435966 292046 436022 292102
rect 435594 291922 435650 291978
rect 435718 291922 435774 291978
rect 435842 291922 435898 291978
rect 435966 291922 436022 291978
rect 408594 280294 408650 280350
rect 408718 280294 408774 280350
rect 408842 280294 408898 280350
rect 408966 280294 409022 280350
rect 408594 280170 408650 280226
rect 408718 280170 408774 280226
rect 408842 280170 408898 280226
rect 408966 280170 409022 280226
rect 408594 280046 408650 280102
rect 408718 280046 408774 280102
rect 408842 280046 408898 280102
rect 408966 280046 409022 280102
rect 408594 279922 408650 279978
rect 408718 279922 408774 279978
rect 408842 279922 408898 279978
rect 408966 279922 409022 279978
rect 404874 256294 404930 256350
rect 404998 256294 405054 256350
rect 405122 256294 405178 256350
rect 405246 256294 405302 256350
rect 404874 256170 404930 256226
rect 404998 256170 405054 256226
rect 405122 256170 405178 256226
rect 405246 256170 405302 256226
rect 404874 256046 404930 256102
rect 404998 256046 405054 256102
rect 405122 256046 405178 256102
rect 405246 256046 405302 256102
rect 404874 255922 404930 255978
rect 404998 255922 405054 255978
rect 405122 255922 405178 255978
rect 405246 255922 405302 255978
rect 402332 248462 402388 248518
rect 407372 251702 407428 251758
rect 433878 280294 433934 280350
rect 434002 280294 434058 280350
rect 433878 280170 433934 280226
rect 434002 280170 434058 280226
rect 433878 280046 433934 280102
rect 434002 280046 434058 280102
rect 433878 279922 433934 279978
rect 434002 279922 434058 279978
rect 418518 274294 418574 274350
rect 418642 274294 418698 274350
rect 418518 274170 418574 274226
rect 418642 274170 418698 274226
rect 418518 274046 418574 274102
rect 418642 274046 418698 274102
rect 418518 273922 418574 273978
rect 418642 273922 418698 273978
rect 435594 274294 435650 274350
rect 435718 274294 435774 274350
rect 435842 274294 435898 274350
rect 435966 274294 436022 274350
rect 435594 274170 435650 274226
rect 435718 274170 435774 274226
rect 435842 274170 435898 274226
rect 435966 274170 436022 274226
rect 435594 274046 435650 274102
rect 435718 274046 435774 274102
rect 435842 274046 435898 274102
rect 435966 274046 436022 274102
rect 435594 273922 435650 273978
rect 435718 273922 435774 273978
rect 435842 273922 435898 273978
rect 435966 273922 436022 273978
rect 414652 269556 414708 269578
rect 414652 269522 414708 269556
rect 428316 268802 428372 268858
rect 408594 262294 408650 262350
rect 408718 262294 408774 262350
rect 408842 262294 408898 262350
rect 408966 262294 409022 262350
rect 408594 262170 408650 262226
rect 408718 262170 408774 262226
rect 408842 262170 408898 262226
rect 408966 262170 409022 262226
rect 408594 262046 408650 262102
rect 408718 262046 408774 262102
rect 408842 262046 408898 262102
rect 408966 262046 409022 262102
rect 408594 261922 408650 261978
rect 408718 261922 408774 261978
rect 408842 261922 408898 261978
rect 408966 261922 409022 261978
rect 404874 238294 404930 238350
rect 404998 238294 405054 238350
rect 405122 238294 405178 238350
rect 405246 238294 405302 238350
rect 404874 238170 404930 238226
rect 404998 238170 405054 238226
rect 405122 238170 405178 238226
rect 405246 238170 405302 238226
rect 404874 238046 404930 238102
rect 404998 238046 405054 238102
rect 405122 238046 405178 238102
rect 405246 238046 405302 238102
rect 404874 237922 404930 237978
rect 404998 237922 405054 237978
rect 405122 237922 405178 237978
rect 405246 237922 405302 237978
rect 377874 226294 377930 226350
rect 377998 226294 378054 226350
rect 378122 226294 378178 226350
rect 378246 226294 378302 226350
rect 377874 226170 377930 226226
rect 377998 226170 378054 226226
rect 378122 226170 378178 226226
rect 378246 226170 378302 226226
rect 377874 226046 377930 226102
rect 377998 226046 378054 226102
rect 378122 226046 378178 226102
rect 378246 226046 378302 226102
rect 377874 225922 377930 225978
rect 377998 225922 378054 225978
rect 378122 225922 378178 225978
rect 378246 225922 378302 225978
rect 374154 202294 374210 202350
rect 374278 202294 374334 202350
rect 374402 202294 374458 202350
rect 374526 202294 374582 202350
rect 374154 202170 374210 202226
rect 374278 202170 374334 202226
rect 374402 202170 374458 202226
rect 374526 202170 374582 202226
rect 374154 202046 374210 202102
rect 374278 202046 374334 202102
rect 374402 202046 374458 202102
rect 374526 202046 374582 202102
rect 374154 201922 374210 201978
rect 374278 201922 374334 201978
rect 374402 201922 374458 201978
rect 374526 201922 374582 201978
rect 352716 198962 352772 199018
rect 351820 195182 351876 195238
rect 347154 190294 347210 190350
rect 347278 190294 347334 190350
rect 347402 190294 347458 190350
rect 347526 190294 347582 190350
rect 347154 190170 347210 190226
rect 347278 190170 347334 190226
rect 347402 190170 347458 190226
rect 347526 190170 347582 190226
rect 347154 190046 347210 190102
rect 347278 190046 347334 190102
rect 347402 190046 347458 190102
rect 347526 190046 347582 190102
rect 347154 189922 347210 189978
rect 347278 189922 347334 189978
rect 347402 189922 347458 189978
rect 347526 189922 347582 189978
rect 343434 184294 343490 184350
rect 343558 184294 343614 184350
rect 343682 184294 343738 184350
rect 343806 184294 343862 184350
rect 343434 184170 343490 184226
rect 343558 184170 343614 184226
rect 343682 184170 343738 184226
rect 343806 184170 343862 184226
rect 343434 184046 343490 184102
rect 343558 184046 343614 184102
rect 343682 184046 343738 184102
rect 343806 184046 343862 184102
rect 343434 183922 343490 183978
rect 343558 183922 343614 183978
rect 343682 183922 343738 183978
rect 343806 183922 343862 183978
rect 343434 166294 343490 166350
rect 343558 166294 343614 166350
rect 343682 166294 343738 166350
rect 343806 166294 343862 166350
rect 343434 166170 343490 166226
rect 343558 166170 343614 166226
rect 343682 166170 343738 166226
rect 343806 166170 343862 166226
rect 343434 166046 343490 166102
rect 343558 166046 343614 166102
rect 343682 166046 343738 166102
rect 343806 166046 343862 166102
rect 343434 165922 343490 165978
rect 343558 165922 343614 165978
rect 343682 165922 343738 165978
rect 343806 165922 343862 165978
rect 334460 133442 334516 133498
rect 334460 131282 334516 131338
rect 334460 131102 334516 131158
rect 334460 126782 334516 126838
rect 334460 125162 334516 125218
rect 343434 148294 343490 148350
rect 343558 148294 343614 148350
rect 343682 148294 343738 148350
rect 343806 148294 343862 148350
rect 343434 148170 343490 148226
rect 343558 148170 343614 148226
rect 343682 148170 343738 148226
rect 343806 148170 343862 148226
rect 343434 148046 343490 148102
rect 343558 148046 343614 148102
rect 343682 148046 343738 148102
rect 343806 148046 343862 148102
rect 343434 147922 343490 147978
rect 343558 147922 343614 147978
rect 343682 147922 343738 147978
rect 343806 147922 343862 147978
rect 347788 192482 347844 192538
rect 371878 190294 371934 190350
rect 372002 190294 372058 190350
rect 371878 190170 371934 190226
rect 372002 190170 372058 190226
rect 371878 190046 371934 190102
rect 372002 190046 372058 190102
rect 371878 189922 371934 189978
rect 372002 189922 372058 189978
rect 356518 184294 356574 184350
rect 356642 184294 356698 184350
rect 356518 184170 356574 184226
rect 356642 184170 356698 184226
rect 356518 184046 356574 184102
rect 356642 184046 356698 184102
rect 356518 183922 356574 183978
rect 356642 183922 356698 183978
rect 374154 184294 374210 184350
rect 374278 184294 374334 184350
rect 374402 184294 374458 184350
rect 374526 184294 374582 184350
rect 374154 184170 374210 184226
rect 374278 184170 374334 184226
rect 374402 184170 374458 184226
rect 374526 184170 374582 184226
rect 374154 184046 374210 184102
rect 374278 184046 374334 184102
rect 374402 184046 374458 184102
rect 374526 184046 374582 184102
rect 374154 183922 374210 183978
rect 374278 183922 374334 183978
rect 374402 183922 374458 183978
rect 374526 183922 374582 183978
rect 347154 172294 347210 172350
rect 347278 172294 347334 172350
rect 347402 172294 347458 172350
rect 347526 172294 347582 172350
rect 347154 172170 347210 172226
rect 347278 172170 347334 172226
rect 347402 172170 347458 172226
rect 347526 172170 347582 172226
rect 347154 172046 347210 172102
rect 347278 172046 347334 172102
rect 347402 172046 347458 172102
rect 347526 172046 347582 172102
rect 347154 171922 347210 171978
rect 347278 171922 347334 171978
rect 347402 171922 347458 171978
rect 347526 171922 347582 171978
rect 347154 154294 347210 154350
rect 347278 154294 347334 154350
rect 347402 154294 347458 154350
rect 347526 154294 347582 154350
rect 347154 154170 347210 154226
rect 347278 154170 347334 154226
rect 347402 154170 347458 154226
rect 347526 154170 347582 154226
rect 347154 154046 347210 154102
rect 347278 154046 347334 154102
rect 347402 154046 347458 154102
rect 347526 154046 347582 154102
rect 347154 153922 347210 153978
rect 347278 153922 347334 153978
rect 347402 153922 347458 153978
rect 347526 153922 347582 153978
rect 374154 166294 374210 166350
rect 374278 166294 374334 166350
rect 374402 166294 374458 166350
rect 374526 166294 374582 166350
rect 374154 166170 374210 166226
rect 374278 166170 374334 166226
rect 374402 166170 374458 166226
rect 374526 166170 374582 166226
rect 374154 166046 374210 166102
rect 374278 166046 374334 166102
rect 374402 166046 374458 166102
rect 374526 166046 374582 166102
rect 374154 165922 374210 165978
rect 374278 165922 374334 165978
rect 374402 165922 374458 165978
rect 374526 165922 374582 165978
rect 374154 148294 374210 148350
rect 374278 148294 374334 148350
rect 374402 148294 374458 148350
rect 374526 148294 374582 148350
rect 374154 148170 374210 148226
rect 374278 148170 374334 148226
rect 374402 148170 374458 148226
rect 374526 148170 374582 148226
rect 374154 148046 374210 148102
rect 374278 148046 374334 148102
rect 374402 148046 374458 148102
rect 374526 148046 374582 148102
rect 374154 147922 374210 147978
rect 374278 147922 374334 147978
rect 374402 147922 374458 147978
rect 374526 147922 374582 147978
rect 347154 136294 347210 136350
rect 347278 136294 347334 136350
rect 347402 136294 347458 136350
rect 347526 136294 347582 136350
rect 347154 136170 347210 136226
rect 347278 136170 347334 136226
rect 347402 136170 347458 136226
rect 347526 136170 347582 136226
rect 347154 136046 347210 136102
rect 347278 136046 347334 136102
rect 347402 136046 347458 136102
rect 347526 136046 347582 136102
rect 347154 135922 347210 135978
rect 347278 135922 347334 135978
rect 347402 135922 347458 135978
rect 347526 135922 347582 135978
rect 343434 130294 343490 130350
rect 343558 130294 343614 130350
rect 343682 130294 343738 130350
rect 343806 130294 343862 130350
rect 343434 130170 343490 130226
rect 343558 130170 343614 130226
rect 343682 130170 343738 130226
rect 343806 130170 343862 130226
rect 338492 124262 338548 124318
rect 272518 58294 272574 58350
rect 272642 58294 272698 58350
rect 272518 58170 272574 58226
rect 272642 58170 272698 58226
rect 272518 58046 272574 58102
rect 272642 58046 272698 58102
rect 272518 57922 272574 57978
rect 272642 57922 272698 57978
rect 281994 58294 282050 58350
rect 282118 58294 282174 58350
rect 282242 58294 282298 58350
rect 282366 58294 282422 58350
rect 281994 58170 282050 58226
rect 282118 58170 282174 58226
rect 282242 58170 282298 58226
rect 282366 58170 282422 58226
rect 281994 58046 282050 58102
rect 282118 58046 282174 58102
rect 282242 58046 282298 58102
rect 282366 58046 282422 58102
rect 281994 57922 282050 57978
rect 282118 57922 282174 57978
rect 282242 57922 282298 57978
rect 282366 57922 282422 57978
rect 270060 55502 270116 55558
rect 254994 46294 255050 46350
rect 255118 46294 255174 46350
rect 255242 46294 255298 46350
rect 255366 46294 255422 46350
rect 254994 46170 255050 46226
rect 255118 46170 255174 46226
rect 255242 46170 255298 46226
rect 255366 46170 255422 46226
rect 254994 46046 255050 46102
rect 255118 46046 255174 46102
rect 255242 46046 255298 46102
rect 255366 46046 255422 46102
rect 254994 45922 255050 45978
rect 255118 45922 255174 45978
rect 255242 45922 255298 45978
rect 255366 45922 255422 45978
rect 251274 40294 251330 40350
rect 251398 40294 251454 40350
rect 251522 40294 251578 40350
rect 251646 40294 251702 40350
rect 251274 40170 251330 40226
rect 251398 40170 251454 40226
rect 251522 40170 251578 40226
rect 251646 40170 251702 40226
rect 251274 40046 251330 40102
rect 251398 40046 251454 40102
rect 251522 40046 251578 40102
rect 251646 40046 251702 40102
rect 251274 39922 251330 39978
rect 251398 39922 251454 39978
rect 251522 39922 251578 39978
rect 251646 39922 251702 39978
rect 224274 28294 224330 28350
rect 224398 28294 224454 28350
rect 224522 28294 224578 28350
rect 224646 28294 224702 28350
rect 224274 28170 224330 28226
rect 224398 28170 224454 28226
rect 224522 28170 224578 28226
rect 224646 28170 224702 28226
rect 224274 28046 224330 28102
rect 224398 28046 224454 28102
rect 224522 28046 224578 28102
rect 224646 28046 224702 28102
rect 224274 27922 224330 27978
rect 224398 27922 224454 27978
rect 224522 27922 224578 27978
rect 224646 27922 224702 27978
rect 224274 10294 224330 10350
rect 224398 10294 224454 10350
rect 224522 10294 224578 10350
rect 224646 10294 224702 10350
rect 224274 10170 224330 10226
rect 224398 10170 224454 10226
rect 224522 10170 224578 10226
rect 224646 10170 224702 10226
rect 224274 10046 224330 10102
rect 224398 10046 224454 10102
rect 224522 10046 224578 10102
rect 224646 10046 224702 10102
rect 224274 9922 224330 9978
rect 224398 9922 224454 9978
rect 224522 9922 224578 9978
rect 224646 9922 224702 9978
rect 224274 -1176 224330 -1120
rect 224398 -1176 224454 -1120
rect 224522 -1176 224578 -1120
rect 224646 -1176 224702 -1120
rect 224274 -1300 224330 -1244
rect 224398 -1300 224454 -1244
rect 224522 -1300 224578 -1244
rect 224646 -1300 224702 -1244
rect 224274 -1424 224330 -1368
rect 224398 -1424 224454 -1368
rect 224522 -1424 224578 -1368
rect 224646 -1424 224702 -1368
rect 224274 -1548 224330 -1492
rect 224398 -1548 224454 -1492
rect 224522 -1548 224578 -1492
rect 224646 -1548 224702 -1492
rect 251274 22294 251330 22350
rect 251398 22294 251454 22350
rect 251522 22294 251578 22350
rect 251646 22294 251702 22350
rect 251274 22170 251330 22226
rect 251398 22170 251454 22226
rect 251522 22170 251578 22226
rect 251646 22170 251702 22226
rect 251274 22046 251330 22102
rect 251398 22046 251454 22102
rect 251522 22046 251578 22102
rect 251646 22046 251702 22102
rect 251274 21922 251330 21978
rect 251398 21922 251454 21978
rect 251522 21922 251578 21978
rect 251646 21922 251702 21978
rect 251274 4294 251330 4350
rect 251398 4294 251454 4350
rect 251522 4294 251578 4350
rect 251646 4294 251702 4350
rect 251274 4170 251330 4226
rect 251398 4170 251454 4226
rect 251522 4170 251578 4226
rect 251646 4170 251702 4226
rect 251274 4046 251330 4102
rect 251398 4046 251454 4102
rect 251522 4046 251578 4102
rect 251646 4046 251702 4102
rect 251274 3922 251330 3978
rect 251398 3922 251454 3978
rect 251522 3922 251578 3978
rect 251646 3922 251702 3978
rect 251274 -216 251330 -160
rect 251398 -216 251454 -160
rect 251522 -216 251578 -160
rect 251646 -216 251702 -160
rect 251274 -340 251330 -284
rect 251398 -340 251454 -284
rect 251522 -340 251578 -284
rect 251646 -340 251702 -284
rect 251274 -464 251330 -408
rect 251398 -464 251454 -408
rect 251522 -464 251578 -408
rect 251646 -464 251702 -408
rect 251274 -588 251330 -532
rect 251398 -588 251454 -532
rect 251522 -588 251578 -532
rect 251646 -588 251702 -532
rect 272518 40294 272574 40350
rect 272642 40294 272698 40350
rect 272518 40170 272574 40226
rect 272642 40170 272698 40226
rect 272518 40046 272574 40102
rect 272642 40046 272698 40102
rect 272518 39922 272574 39978
rect 272642 39922 272698 39978
rect 281994 40294 282050 40350
rect 282118 40294 282174 40350
rect 282242 40294 282298 40350
rect 282366 40294 282422 40350
rect 281994 40170 282050 40226
rect 282118 40170 282174 40226
rect 282242 40170 282298 40226
rect 282366 40170 282422 40226
rect 281994 40046 282050 40102
rect 282118 40046 282174 40102
rect 282242 40046 282298 40102
rect 282366 40046 282422 40102
rect 281994 39922 282050 39978
rect 282118 39922 282174 39978
rect 282242 39922 282298 39978
rect 282366 39922 282422 39978
rect 254994 28294 255050 28350
rect 255118 28294 255174 28350
rect 255242 28294 255298 28350
rect 255366 28294 255422 28350
rect 254994 28170 255050 28226
rect 255118 28170 255174 28226
rect 255242 28170 255298 28226
rect 255366 28170 255422 28226
rect 254994 28046 255050 28102
rect 255118 28046 255174 28102
rect 255242 28046 255298 28102
rect 255366 28046 255422 28102
rect 254994 27922 255050 27978
rect 255118 27922 255174 27978
rect 255242 27922 255298 27978
rect 255366 27922 255422 27978
rect 254994 10294 255050 10350
rect 255118 10294 255174 10350
rect 255242 10294 255298 10350
rect 255366 10294 255422 10350
rect 254994 10170 255050 10226
rect 255118 10170 255174 10226
rect 255242 10170 255298 10226
rect 255366 10170 255422 10226
rect 254994 10046 255050 10102
rect 255118 10046 255174 10102
rect 255242 10046 255298 10102
rect 255366 10046 255422 10102
rect 254994 9922 255050 9978
rect 255118 9922 255174 9978
rect 255242 9922 255298 9978
rect 255366 9922 255422 9978
rect 254994 -1176 255050 -1120
rect 255118 -1176 255174 -1120
rect 255242 -1176 255298 -1120
rect 255366 -1176 255422 -1120
rect 254994 -1300 255050 -1244
rect 255118 -1300 255174 -1244
rect 255242 -1300 255298 -1244
rect 255366 -1300 255422 -1244
rect 254994 -1424 255050 -1368
rect 255118 -1424 255174 -1368
rect 255242 -1424 255298 -1368
rect 255366 -1424 255422 -1368
rect 254994 -1548 255050 -1492
rect 255118 -1548 255174 -1492
rect 255242 -1548 255298 -1492
rect 255366 -1548 255422 -1492
rect 281994 22294 282050 22350
rect 282118 22294 282174 22350
rect 282242 22294 282298 22350
rect 282366 22294 282422 22350
rect 281994 22170 282050 22226
rect 282118 22170 282174 22226
rect 282242 22170 282298 22226
rect 282366 22170 282422 22226
rect 281994 22046 282050 22102
rect 282118 22046 282174 22102
rect 282242 22046 282298 22102
rect 282366 22046 282422 22102
rect 281994 21922 282050 21978
rect 282118 21922 282174 21978
rect 282242 21922 282298 21978
rect 282366 21922 282422 21978
rect 281994 4294 282050 4350
rect 282118 4294 282174 4350
rect 282242 4294 282298 4350
rect 282366 4294 282422 4350
rect 281994 4170 282050 4226
rect 282118 4170 282174 4226
rect 282242 4170 282298 4226
rect 282366 4170 282422 4226
rect 281994 4046 282050 4102
rect 282118 4046 282174 4102
rect 282242 4046 282298 4102
rect 282366 4046 282422 4102
rect 281994 3922 282050 3978
rect 282118 3922 282174 3978
rect 282242 3922 282298 3978
rect 282366 3922 282422 3978
rect 281994 -216 282050 -160
rect 282118 -216 282174 -160
rect 282242 -216 282298 -160
rect 282366 -216 282422 -160
rect 281994 -340 282050 -284
rect 282118 -340 282174 -284
rect 282242 -340 282298 -284
rect 282366 -340 282422 -284
rect 281994 -464 282050 -408
rect 282118 -464 282174 -408
rect 282242 -464 282298 -408
rect 282366 -464 282422 -408
rect 281994 -588 282050 -532
rect 282118 -588 282174 -532
rect 282242 -588 282298 -532
rect 282366 -588 282422 -532
rect 285714 64294 285770 64350
rect 285838 64294 285894 64350
rect 285962 64294 286018 64350
rect 286086 64294 286142 64350
rect 285714 64170 285770 64226
rect 285838 64170 285894 64226
rect 285962 64170 286018 64226
rect 286086 64170 286142 64226
rect 285714 64046 285770 64102
rect 285838 64046 285894 64102
rect 285962 64046 286018 64102
rect 286086 64046 286142 64102
rect 285714 63922 285770 63978
rect 285838 63922 285894 63978
rect 285962 63922 286018 63978
rect 286086 63922 286142 63978
rect 287878 64294 287934 64350
rect 288002 64294 288058 64350
rect 287878 64170 287934 64226
rect 288002 64170 288058 64226
rect 287878 64046 287934 64102
rect 288002 64046 288058 64102
rect 287878 63922 287934 63978
rect 288002 63922 288058 63978
rect 303238 58294 303294 58350
rect 303362 58294 303418 58350
rect 303238 58170 303294 58226
rect 303362 58170 303418 58226
rect 303238 58046 303294 58102
rect 303362 58046 303418 58102
rect 303238 57922 303294 57978
rect 303362 57922 303418 57978
rect 312714 58294 312770 58350
rect 312838 58294 312894 58350
rect 312962 58294 313018 58350
rect 313086 58294 313142 58350
rect 312714 58170 312770 58226
rect 312838 58170 312894 58226
rect 312962 58170 313018 58226
rect 313086 58170 313142 58226
rect 312714 58046 312770 58102
rect 312838 58046 312894 58102
rect 312962 58046 313018 58102
rect 313086 58046 313142 58102
rect 312714 57922 312770 57978
rect 312838 57922 312894 57978
rect 312962 57922 313018 57978
rect 313086 57922 313142 57978
rect 285714 46294 285770 46350
rect 285838 46294 285894 46350
rect 285962 46294 286018 46350
rect 286086 46294 286142 46350
rect 285714 46170 285770 46226
rect 285838 46170 285894 46226
rect 285962 46170 286018 46226
rect 286086 46170 286142 46226
rect 285714 46046 285770 46102
rect 285838 46046 285894 46102
rect 285962 46046 286018 46102
rect 286086 46046 286142 46102
rect 285714 45922 285770 45978
rect 285838 45922 285894 45978
rect 285962 45922 286018 45978
rect 286086 45922 286142 45978
rect 287878 46294 287934 46350
rect 288002 46294 288058 46350
rect 287878 46170 287934 46226
rect 288002 46170 288058 46226
rect 287878 46046 287934 46102
rect 288002 46046 288058 46102
rect 287878 45922 287934 45978
rect 288002 45922 288058 45978
rect 303238 40294 303294 40350
rect 303362 40294 303418 40350
rect 303238 40170 303294 40226
rect 303362 40170 303418 40226
rect 303238 40046 303294 40102
rect 303362 40046 303418 40102
rect 303238 39922 303294 39978
rect 303362 39922 303418 39978
rect 312714 40294 312770 40350
rect 312838 40294 312894 40350
rect 312962 40294 313018 40350
rect 313086 40294 313142 40350
rect 312714 40170 312770 40226
rect 312838 40170 312894 40226
rect 312962 40170 313018 40226
rect 313086 40170 313142 40226
rect 312714 40046 312770 40102
rect 312838 40046 312894 40102
rect 312962 40046 313018 40102
rect 313086 40046 313142 40102
rect 312714 39922 312770 39978
rect 312838 39922 312894 39978
rect 312962 39922 313018 39978
rect 313086 39922 313142 39978
rect 285714 28294 285770 28350
rect 285838 28294 285894 28350
rect 285962 28294 286018 28350
rect 286086 28294 286142 28350
rect 285714 28170 285770 28226
rect 285838 28170 285894 28226
rect 285962 28170 286018 28226
rect 286086 28170 286142 28226
rect 285714 28046 285770 28102
rect 285838 28046 285894 28102
rect 285962 28046 286018 28102
rect 286086 28046 286142 28102
rect 285714 27922 285770 27978
rect 285838 27922 285894 27978
rect 285962 27922 286018 27978
rect 286086 27922 286142 27978
rect 285714 10294 285770 10350
rect 285838 10294 285894 10350
rect 285962 10294 286018 10350
rect 286086 10294 286142 10350
rect 285714 10170 285770 10226
rect 285838 10170 285894 10226
rect 285962 10170 286018 10226
rect 286086 10170 286142 10226
rect 285714 10046 285770 10102
rect 285838 10046 285894 10102
rect 285962 10046 286018 10102
rect 286086 10046 286142 10102
rect 285714 9922 285770 9978
rect 285838 9922 285894 9978
rect 285962 9922 286018 9978
rect 286086 9922 286142 9978
rect 285714 -1176 285770 -1120
rect 285838 -1176 285894 -1120
rect 285962 -1176 286018 -1120
rect 286086 -1176 286142 -1120
rect 285714 -1300 285770 -1244
rect 285838 -1300 285894 -1244
rect 285962 -1300 286018 -1244
rect 286086 -1300 286142 -1244
rect 285714 -1424 285770 -1368
rect 285838 -1424 285894 -1368
rect 285962 -1424 286018 -1368
rect 286086 -1424 286142 -1368
rect 285714 -1548 285770 -1492
rect 285838 -1548 285894 -1492
rect 285962 -1548 286018 -1492
rect 286086 -1548 286142 -1492
rect 312714 22294 312770 22350
rect 312838 22294 312894 22350
rect 312962 22294 313018 22350
rect 313086 22294 313142 22350
rect 312714 22170 312770 22226
rect 312838 22170 312894 22226
rect 312962 22170 313018 22226
rect 313086 22170 313142 22226
rect 312714 22046 312770 22102
rect 312838 22046 312894 22102
rect 312962 22046 313018 22102
rect 313086 22046 313142 22102
rect 312714 21922 312770 21978
rect 312838 21922 312894 21978
rect 312962 21922 313018 21978
rect 313086 21922 313142 21978
rect 312714 4294 312770 4350
rect 312838 4294 312894 4350
rect 312962 4294 313018 4350
rect 313086 4294 313142 4350
rect 312714 4170 312770 4226
rect 312838 4170 312894 4226
rect 312962 4170 313018 4226
rect 313086 4170 313142 4226
rect 312714 4046 312770 4102
rect 312838 4046 312894 4102
rect 312962 4046 313018 4102
rect 313086 4046 313142 4102
rect 312714 3922 312770 3978
rect 312838 3922 312894 3978
rect 312962 3922 313018 3978
rect 313086 3922 313142 3978
rect 312714 -216 312770 -160
rect 312838 -216 312894 -160
rect 312962 -216 313018 -160
rect 313086 -216 313142 -160
rect 312714 -340 312770 -284
rect 312838 -340 312894 -284
rect 312962 -340 313018 -284
rect 313086 -340 313142 -284
rect 312714 -464 312770 -408
rect 312838 -464 312894 -408
rect 312962 -464 313018 -408
rect 313086 -464 313142 -408
rect 312714 -588 312770 -532
rect 312838 -588 312894 -532
rect 312962 -588 313018 -532
rect 313086 -588 313142 -532
rect 316434 64294 316490 64350
rect 316558 64294 316614 64350
rect 316682 64294 316738 64350
rect 316806 64294 316862 64350
rect 316434 64170 316490 64226
rect 316558 64170 316614 64226
rect 316682 64170 316738 64226
rect 316806 64170 316862 64226
rect 316434 64046 316490 64102
rect 316558 64046 316614 64102
rect 316682 64046 316738 64102
rect 316806 64046 316862 64102
rect 316434 63922 316490 63978
rect 316558 63922 316614 63978
rect 316682 63922 316738 63978
rect 316806 63922 316862 63978
rect 318598 64294 318654 64350
rect 318722 64294 318778 64350
rect 318598 64170 318654 64226
rect 318722 64170 318778 64226
rect 318598 64046 318654 64102
rect 318722 64046 318778 64102
rect 318598 63922 318654 63978
rect 318722 63922 318778 63978
rect 343434 130046 343490 130102
rect 343558 130046 343614 130102
rect 343682 130046 343738 130102
rect 343806 130046 343862 130102
rect 343434 129922 343490 129978
rect 343558 129922 343614 129978
rect 343682 129922 343738 129978
rect 343806 129922 343862 129978
rect 345212 122462 345268 122518
rect 343434 112294 343490 112350
rect 343558 112294 343614 112350
rect 343682 112294 343738 112350
rect 343806 112294 343862 112350
rect 343434 112170 343490 112226
rect 343558 112170 343614 112226
rect 343682 112170 343738 112226
rect 343806 112170 343862 112226
rect 343434 112046 343490 112102
rect 343558 112046 343614 112102
rect 343682 112046 343738 112102
rect 343806 112046 343862 112102
rect 343434 111922 343490 111978
rect 343558 111922 343614 111978
rect 343682 111922 343738 111978
rect 343806 111922 343862 111978
rect 343434 94294 343490 94350
rect 343558 94294 343614 94350
rect 343682 94294 343738 94350
rect 343806 94294 343862 94350
rect 343434 94170 343490 94226
rect 343558 94170 343614 94226
rect 343682 94170 343738 94226
rect 343806 94170 343862 94226
rect 343434 94046 343490 94102
rect 343558 94046 343614 94102
rect 343682 94046 343738 94102
rect 343806 94046 343862 94102
rect 343434 93922 343490 93978
rect 343558 93922 343614 93978
rect 343682 93922 343738 93978
rect 343806 93922 343862 93978
rect 343434 76294 343490 76350
rect 343558 76294 343614 76350
rect 343682 76294 343738 76350
rect 343806 76294 343862 76350
rect 343434 76170 343490 76226
rect 343558 76170 343614 76226
rect 343682 76170 343738 76226
rect 343806 76170 343862 76226
rect 343434 76046 343490 76102
rect 343558 76046 343614 76102
rect 343682 76046 343738 76102
rect 343806 76046 343862 76102
rect 343434 75922 343490 75978
rect 343558 75922 343614 75978
rect 343682 75922 343738 75978
rect 343806 75922 343862 75978
rect 343434 58294 343490 58350
rect 343558 58294 343614 58350
rect 343682 58294 343738 58350
rect 343806 58294 343862 58350
rect 343434 58170 343490 58226
rect 343558 58170 343614 58226
rect 343682 58170 343738 58226
rect 343806 58170 343862 58226
rect 343434 58046 343490 58102
rect 343558 58046 343614 58102
rect 343682 58046 343738 58102
rect 343806 58046 343862 58102
rect 343434 57922 343490 57978
rect 343558 57922 343614 57978
rect 343682 57922 343738 57978
rect 343806 57922 343862 57978
rect 316434 46294 316490 46350
rect 316558 46294 316614 46350
rect 316682 46294 316738 46350
rect 316806 46294 316862 46350
rect 316434 46170 316490 46226
rect 316558 46170 316614 46226
rect 316682 46170 316738 46226
rect 316806 46170 316862 46226
rect 316434 46046 316490 46102
rect 316558 46046 316614 46102
rect 316682 46046 316738 46102
rect 316806 46046 316862 46102
rect 316434 45922 316490 45978
rect 316558 45922 316614 45978
rect 316682 45922 316738 45978
rect 316806 45922 316862 45978
rect 318598 46294 318654 46350
rect 318722 46294 318778 46350
rect 318598 46170 318654 46226
rect 318722 46170 318778 46226
rect 318598 46046 318654 46102
rect 318722 46046 318778 46102
rect 318598 45922 318654 45978
rect 318722 45922 318778 45978
rect 316434 28294 316490 28350
rect 316558 28294 316614 28350
rect 316682 28294 316738 28350
rect 316806 28294 316862 28350
rect 316434 28170 316490 28226
rect 316558 28170 316614 28226
rect 316682 28170 316738 28226
rect 316806 28170 316862 28226
rect 316434 28046 316490 28102
rect 316558 28046 316614 28102
rect 316682 28046 316738 28102
rect 316806 28046 316862 28102
rect 316434 27922 316490 27978
rect 316558 27922 316614 27978
rect 316682 27922 316738 27978
rect 316806 27922 316862 27978
rect 316434 10294 316490 10350
rect 316558 10294 316614 10350
rect 316682 10294 316738 10350
rect 316806 10294 316862 10350
rect 316434 10170 316490 10226
rect 316558 10170 316614 10226
rect 316682 10170 316738 10226
rect 316806 10170 316862 10226
rect 316434 10046 316490 10102
rect 316558 10046 316614 10102
rect 316682 10046 316738 10102
rect 316806 10046 316862 10102
rect 316434 9922 316490 9978
rect 316558 9922 316614 9978
rect 316682 9922 316738 9978
rect 316806 9922 316862 9978
rect 316434 -1176 316490 -1120
rect 316558 -1176 316614 -1120
rect 316682 -1176 316738 -1120
rect 316806 -1176 316862 -1120
rect 316434 -1300 316490 -1244
rect 316558 -1300 316614 -1244
rect 316682 -1300 316738 -1244
rect 316806 -1300 316862 -1244
rect 316434 -1424 316490 -1368
rect 316558 -1424 316614 -1368
rect 316682 -1424 316738 -1368
rect 316806 -1424 316862 -1368
rect 316434 -1548 316490 -1492
rect 316558 -1548 316614 -1492
rect 316682 -1548 316738 -1492
rect 316806 -1548 316862 -1492
rect 371878 136294 371934 136350
rect 372002 136294 372058 136350
rect 371878 136170 371934 136226
rect 372002 136170 372058 136226
rect 371878 136046 371934 136102
rect 372002 136046 372058 136102
rect 371878 135922 371934 135978
rect 372002 135922 372058 135978
rect 347154 118294 347210 118350
rect 347278 118294 347334 118350
rect 347402 118294 347458 118350
rect 347526 118294 347582 118350
rect 347154 118170 347210 118226
rect 347278 118170 347334 118226
rect 347402 118170 347458 118226
rect 347526 118170 347582 118226
rect 347154 118046 347210 118102
rect 347278 118046 347334 118102
rect 347402 118046 347458 118102
rect 347526 118046 347582 118102
rect 347154 117922 347210 117978
rect 347278 117922 347334 117978
rect 347402 117922 347458 117978
rect 347526 117922 347582 117978
rect 347154 100294 347210 100350
rect 347278 100294 347334 100350
rect 347402 100294 347458 100350
rect 347526 100294 347582 100350
rect 347154 100170 347210 100226
rect 347278 100170 347334 100226
rect 347402 100170 347458 100226
rect 347526 100170 347582 100226
rect 347154 100046 347210 100102
rect 347278 100046 347334 100102
rect 347402 100046 347458 100102
rect 347526 100046 347582 100102
rect 347154 99922 347210 99978
rect 347278 99922 347334 99978
rect 347402 99922 347458 99978
rect 347526 99922 347582 99978
rect 347154 82294 347210 82350
rect 347278 82294 347334 82350
rect 347402 82294 347458 82350
rect 347526 82294 347582 82350
rect 347154 82170 347210 82226
rect 347278 82170 347334 82226
rect 347402 82170 347458 82226
rect 347526 82170 347582 82226
rect 347154 82046 347210 82102
rect 347278 82046 347334 82102
rect 347402 82046 347458 82102
rect 347526 82046 347582 82102
rect 347154 81922 347210 81978
rect 347278 81922 347334 81978
rect 347402 81922 347458 81978
rect 347526 81922 347582 81978
rect 356518 130294 356574 130350
rect 356642 130294 356698 130350
rect 356518 130170 356574 130226
rect 356642 130170 356698 130226
rect 356518 130046 356574 130102
rect 356642 130046 356698 130102
rect 356518 129922 356574 129978
rect 356642 129922 356698 129978
rect 374154 130294 374210 130350
rect 374278 130294 374334 130350
rect 374402 130294 374458 130350
rect 374526 130294 374582 130350
rect 374154 130170 374210 130226
rect 374278 130170 374334 130226
rect 374402 130170 374458 130226
rect 374526 130170 374582 130226
rect 374154 130046 374210 130102
rect 374278 130046 374334 130102
rect 374402 130046 374458 130102
rect 374526 130046 374582 130102
rect 374154 129922 374210 129978
rect 374278 129922 374334 129978
rect 374402 129922 374458 129978
rect 374526 129922 374582 129978
rect 352716 128402 352772 128458
rect 351932 120842 351988 120898
rect 377874 208294 377930 208350
rect 377998 208294 378054 208350
rect 378122 208294 378178 208350
rect 378246 208294 378302 208350
rect 377874 208170 377930 208226
rect 377998 208170 378054 208226
rect 378122 208170 378178 208226
rect 378246 208170 378302 208226
rect 377874 208046 377930 208102
rect 377998 208046 378054 208102
rect 378122 208046 378178 208102
rect 378246 208046 378302 208102
rect 377874 207922 377930 207978
rect 377998 207922 378054 207978
rect 378122 207922 378178 207978
rect 378246 207922 378302 207978
rect 387238 202294 387294 202350
rect 387362 202294 387418 202350
rect 387238 202170 387294 202226
rect 387362 202170 387418 202226
rect 387238 202046 387294 202102
rect 387362 202046 387418 202102
rect 387238 201922 387294 201978
rect 387362 201922 387418 201978
rect 377874 190294 377930 190350
rect 377998 190294 378054 190350
rect 378122 190294 378178 190350
rect 378246 190294 378302 190350
rect 377874 190170 377930 190226
rect 377998 190170 378054 190226
rect 378122 190170 378178 190226
rect 378246 190170 378302 190226
rect 377874 190046 377930 190102
rect 377998 190046 378054 190102
rect 378122 190046 378178 190102
rect 378246 190046 378302 190102
rect 377874 189922 377930 189978
rect 377998 189922 378054 189978
rect 378122 189922 378178 189978
rect 378246 189922 378302 189978
rect 404874 220294 404930 220350
rect 404998 220294 405054 220350
rect 405122 220294 405178 220350
rect 405246 220294 405302 220350
rect 404874 220170 404930 220226
rect 404998 220170 405054 220226
rect 405122 220170 405178 220226
rect 405246 220170 405302 220226
rect 404874 220046 404930 220102
rect 404998 220046 405054 220102
rect 405122 220046 405178 220102
rect 405246 220046 405302 220102
rect 404874 219922 404930 219978
rect 404998 219922 405054 219978
rect 405122 219922 405178 219978
rect 405246 219922 405302 219978
rect 394828 188882 394884 188938
rect 429212 267362 429268 267418
rect 429212 266282 429268 266338
rect 428316 265382 428372 265438
rect 428428 263762 428484 263818
rect 433878 262294 433934 262350
rect 434002 262294 434058 262350
rect 433878 262170 433934 262226
rect 434002 262170 434058 262226
rect 433878 262046 433934 262102
rect 434002 262046 434058 262102
rect 433878 261922 433934 261978
rect 434002 261922 434058 261978
rect 428428 260342 428484 260398
rect 418518 256294 418574 256350
rect 418642 256294 418698 256350
rect 418518 256170 418574 256226
rect 418642 256170 418698 256226
rect 418518 256046 418574 256102
rect 418642 256046 418698 256102
rect 418518 255922 418574 255978
rect 418642 255922 418698 255978
rect 435594 256294 435650 256350
rect 435718 256294 435774 256350
rect 435842 256294 435898 256350
rect 435966 256294 436022 256350
rect 435594 256170 435650 256226
rect 435718 256170 435774 256226
rect 435842 256170 435898 256226
rect 435966 256170 436022 256226
rect 435594 256046 435650 256102
rect 435718 256046 435774 256102
rect 435842 256046 435898 256102
rect 435966 256046 436022 256102
rect 435594 255922 435650 255978
rect 435718 255922 435774 255978
rect 435842 255922 435898 255978
rect 435966 255922 436022 255978
rect 408594 244294 408650 244350
rect 408718 244294 408774 244350
rect 408842 244294 408898 244350
rect 408966 244294 409022 244350
rect 408594 244170 408650 244226
rect 408718 244170 408774 244226
rect 408842 244170 408898 244226
rect 408966 244170 409022 244226
rect 408594 244046 408650 244102
rect 408718 244046 408774 244102
rect 408842 244046 408898 244102
rect 408966 244046 409022 244102
rect 408594 243922 408650 243978
rect 408718 243922 408774 243978
rect 408842 243922 408898 243978
rect 408966 243922 409022 243978
rect 435594 238294 435650 238350
rect 435718 238294 435774 238350
rect 435842 238294 435898 238350
rect 435966 238294 436022 238350
rect 435594 238170 435650 238226
rect 435718 238170 435774 238226
rect 435842 238170 435898 238226
rect 435966 238170 436022 238226
rect 435594 238046 435650 238102
rect 435718 238046 435774 238102
rect 435842 238046 435898 238102
rect 435966 238046 436022 238102
rect 435594 237922 435650 237978
rect 435718 237922 435774 237978
rect 435842 237922 435898 237978
rect 435966 237922 436022 237978
rect 408594 226294 408650 226350
rect 408718 226294 408774 226350
rect 408842 226294 408898 226350
rect 408966 226294 409022 226350
rect 408594 226170 408650 226226
rect 408718 226170 408774 226226
rect 408842 226170 408898 226226
rect 408966 226170 409022 226226
rect 408594 226046 408650 226102
rect 408718 226046 408774 226102
rect 408842 226046 408898 226102
rect 408966 226046 409022 226102
rect 408594 225922 408650 225978
rect 408718 225922 408774 225978
rect 408842 225922 408898 225978
rect 408966 225922 409022 225978
rect 404874 202294 404930 202350
rect 404998 202294 405054 202350
rect 405122 202294 405178 202350
rect 405246 202294 405302 202350
rect 404874 202170 404930 202226
rect 404998 202170 405054 202226
rect 405122 202170 405178 202226
rect 405246 202170 405302 202226
rect 404874 202046 404930 202102
rect 404998 202046 405054 202102
rect 405122 202046 405178 202102
rect 405246 202046 405302 202102
rect 404874 201922 404930 201978
rect 404998 201922 405054 201978
rect 405122 201922 405178 201978
rect 405246 201922 405302 201978
rect 403116 198422 403172 198478
rect 401436 198242 401492 198298
rect 401436 195722 401492 195778
rect 403116 194822 403172 194878
rect 403228 195002 403284 195058
rect 403228 189602 403284 189658
rect 396508 187262 396564 187318
rect 393260 186182 393316 186238
rect 387238 184294 387294 184350
rect 387362 184294 387418 184350
rect 387238 184170 387294 184226
rect 387362 184170 387418 184226
rect 387238 184046 387294 184102
rect 387362 184046 387418 184102
rect 387238 183922 387294 183978
rect 387362 183922 387418 183978
rect 408594 208294 408650 208350
rect 408718 208294 408774 208350
rect 408842 208294 408898 208350
rect 408966 208294 409022 208350
rect 408594 208170 408650 208226
rect 408718 208170 408774 208226
rect 408842 208170 408898 208226
rect 408966 208170 409022 208226
rect 408594 208046 408650 208102
rect 408718 208046 408774 208102
rect 408842 208046 408898 208102
rect 408966 208046 409022 208102
rect 408594 207922 408650 207978
rect 408718 207922 408774 207978
rect 408842 207922 408898 207978
rect 408966 207922 409022 207978
rect 404874 184294 404930 184350
rect 404998 184294 405054 184350
rect 405122 184294 405178 184350
rect 405246 184294 405302 184350
rect 404874 184170 404930 184226
rect 404998 184170 405054 184226
rect 405122 184170 405178 184226
rect 405246 184170 405302 184226
rect 404874 184046 404930 184102
rect 404998 184046 405054 184102
rect 405122 184046 405178 184102
rect 405246 184046 405302 184102
rect 404874 183922 404930 183978
rect 404998 183922 405054 183978
rect 405122 183922 405178 183978
rect 405246 183922 405302 183978
rect 377874 172294 377930 172350
rect 377998 172294 378054 172350
rect 378122 172294 378178 172350
rect 378246 172294 378302 172350
rect 377874 172170 377930 172226
rect 377998 172170 378054 172226
rect 378122 172170 378178 172226
rect 378246 172170 378302 172226
rect 377874 172046 377930 172102
rect 377998 172046 378054 172102
rect 378122 172046 378178 172102
rect 378246 172046 378302 172102
rect 377874 171922 377930 171978
rect 377998 171922 378054 171978
rect 378122 171922 378178 171978
rect 378246 171922 378302 171978
rect 377874 154294 377930 154350
rect 377998 154294 378054 154350
rect 378122 154294 378178 154350
rect 378246 154294 378302 154350
rect 377874 154170 377930 154226
rect 377998 154170 378054 154226
rect 378122 154170 378178 154226
rect 378246 154170 378302 154226
rect 377874 154046 377930 154102
rect 377998 154046 378054 154102
rect 378122 154046 378178 154102
rect 378246 154046 378302 154102
rect 377874 153922 377930 153978
rect 377998 153922 378054 153978
rect 378122 153922 378178 153978
rect 378246 153922 378302 153978
rect 404874 166294 404930 166350
rect 404998 166294 405054 166350
rect 405122 166294 405178 166350
rect 405246 166294 405302 166350
rect 404874 166170 404930 166226
rect 404998 166170 405054 166226
rect 405122 166170 405178 166226
rect 405246 166170 405302 166226
rect 404874 166046 404930 166102
rect 404998 166046 405054 166102
rect 405122 166046 405178 166102
rect 405246 166046 405302 166102
rect 404874 165922 404930 165978
rect 404998 165922 405054 165978
rect 405122 165922 405178 165978
rect 405246 165922 405302 165978
rect 377874 136294 377930 136350
rect 377998 136294 378054 136350
rect 378122 136294 378178 136350
rect 378246 136294 378302 136350
rect 377874 136170 377930 136226
rect 377998 136170 378054 136226
rect 378122 136170 378178 136226
rect 378246 136170 378302 136226
rect 377874 136046 377930 136102
rect 377998 136046 378054 136102
rect 378122 136046 378178 136102
rect 378246 136046 378302 136102
rect 377874 135922 377930 135978
rect 377998 135922 378054 135978
rect 378122 135922 378178 135978
rect 378246 135922 378302 135978
rect 371878 118294 371934 118350
rect 372002 118294 372058 118350
rect 371878 118170 371934 118226
rect 372002 118170 372058 118226
rect 371878 118046 371934 118102
rect 372002 118046 372058 118102
rect 371878 117922 371934 117978
rect 372002 117922 372058 117978
rect 387238 130294 387294 130350
rect 387362 130294 387418 130350
rect 387238 130170 387294 130226
rect 387362 130170 387418 130226
rect 387238 130046 387294 130102
rect 387362 130046 387418 130102
rect 387238 129922 387294 129978
rect 387362 129922 387418 129978
rect 393260 126644 393316 126658
rect 393260 126602 393316 126644
rect 393372 125342 393428 125398
rect 404874 148294 404930 148350
rect 404998 148294 405054 148350
rect 405122 148294 405178 148350
rect 405246 148294 405302 148350
rect 404874 148170 404930 148226
rect 404998 148170 405054 148226
rect 405122 148170 405178 148226
rect 405246 148170 405302 148226
rect 404874 148046 404930 148102
rect 404998 148046 405054 148102
rect 405122 148046 405178 148102
rect 405246 148046 405302 148102
rect 404874 147922 404930 147978
rect 404998 147922 405054 147978
rect 405122 147922 405178 147978
rect 405246 147922 405302 147978
rect 377874 118294 377930 118350
rect 377998 118294 378054 118350
rect 378122 118294 378178 118350
rect 378246 118294 378302 118350
rect 377874 118170 377930 118226
rect 377998 118170 378054 118226
rect 378122 118170 378178 118226
rect 378246 118170 378302 118226
rect 377874 118046 377930 118102
rect 377998 118046 378054 118102
rect 378122 118046 378178 118102
rect 378246 118046 378302 118102
rect 377874 117922 377930 117978
rect 377998 117922 378054 117978
rect 378122 117922 378178 117978
rect 378246 117922 378302 117978
rect 356518 112294 356574 112350
rect 356642 112294 356698 112350
rect 356518 112170 356574 112226
rect 356642 112170 356698 112226
rect 356518 112046 356574 112102
rect 356642 112046 356698 112102
rect 356518 111922 356574 111978
rect 356642 111922 356698 111978
rect 374154 112294 374210 112350
rect 374278 112294 374334 112350
rect 374402 112294 374458 112350
rect 374526 112294 374582 112350
rect 374154 112170 374210 112226
rect 374278 112170 374334 112226
rect 374402 112170 374458 112226
rect 374526 112170 374582 112226
rect 374154 112046 374210 112102
rect 374278 112046 374334 112102
rect 374402 112046 374458 112102
rect 374526 112046 374582 112102
rect 374154 111922 374210 111978
rect 374278 111922 374334 111978
rect 374402 111922 374458 111978
rect 374526 111922 374582 111978
rect 374154 94294 374210 94350
rect 374278 94294 374334 94350
rect 374402 94294 374458 94350
rect 374526 94294 374582 94350
rect 374154 94170 374210 94226
rect 374278 94170 374334 94226
rect 374402 94170 374458 94226
rect 374526 94170 374582 94226
rect 374154 94046 374210 94102
rect 374278 94046 374334 94102
rect 374402 94046 374458 94102
rect 374526 94046 374582 94102
rect 374154 93922 374210 93978
rect 374278 93922 374334 93978
rect 374402 93922 374458 93978
rect 374526 93922 374582 93978
rect 374154 76294 374210 76350
rect 374278 76294 374334 76350
rect 374402 76294 374458 76350
rect 374526 76294 374582 76350
rect 374154 76170 374210 76226
rect 374278 76170 374334 76226
rect 374402 76170 374458 76226
rect 374526 76170 374582 76226
rect 374154 76046 374210 76102
rect 374278 76046 374334 76102
rect 374402 76046 374458 76102
rect 374526 76046 374582 76102
rect 374154 75922 374210 75978
rect 374278 75922 374334 75978
rect 374402 75922 374458 75978
rect 374526 75922 374582 75978
rect 347154 64294 347210 64350
rect 347278 64294 347334 64350
rect 347402 64294 347458 64350
rect 347526 64294 347582 64350
rect 347154 64170 347210 64226
rect 347278 64170 347334 64226
rect 347402 64170 347458 64226
rect 347526 64170 347582 64226
rect 347154 64046 347210 64102
rect 347278 64046 347334 64102
rect 347402 64046 347458 64102
rect 347526 64046 347582 64102
rect 347154 63922 347210 63978
rect 347278 63922 347334 63978
rect 347402 63922 347458 63978
rect 347526 63922 347582 63978
rect 343434 40294 343490 40350
rect 343558 40294 343614 40350
rect 343682 40294 343738 40350
rect 343806 40294 343862 40350
rect 343434 40170 343490 40226
rect 343558 40170 343614 40226
rect 343682 40170 343738 40226
rect 343806 40170 343862 40226
rect 343434 40046 343490 40102
rect 343558 40046 343614 40102
rect 343682 40046 343738 40102
rect 343806 40046 343862 40102
rect 343434 39922 343490 39978
rect 343558 39922 343614 39978
rect 343682 39922 343738 39978
rect 343806 39922 343862 39978
rect 343434 22294 343490 22350
rect 343558 22294 343614 22350
rect 343682 22294 343738 22350
rect 343806 22294 343862 22350
rect 343434 22170 343490 22226
rect 343558 22170 343614 22226
rect 343682 22170 343738 22226
rect 343806 22170 343862 22226
rect 343434 22046 343490 22102
rect 343558 22046 343614 22102
rect 343682 22046 343738 22102
rect 343806 22046 343862 22102
rect 343434 21922 343490 21978
rect 343558 21922 343614 21978
rect 343682 21922 343738 21978
rect 343806 21922 343862 21978
rect 343434 4294 343490 4350
rect 343558 4294 343614 4350
rect 343682 4294 343738 4350
rect 343806 4294 343862 4350
rect 343434 4170 343490 4226
rect 343558 4170 343614 4226
rect 343682 4170 343738 4226
rect 343806 4170 343862 4226
rect 343434 4046 343490 4102
rect 343558 4046 343614 4102
rect 343682 4046 343738 4102
rect 343806 4046 343862 4102
rect 343434 3922 343490 3978
rect 343558 3922 343614 3978
rect 343682 3922 343738 3978
rect 343806 3922 343862 3978
rect 343434 -216 343490 -160
rect 343558 -216 343614 -160
rect 343682 -216 343738 -160
rect 343806 -216 343862 -160
rect 343434 -340 343490 -284
rect 343558 -340 343614 -284
rect 343682 -340 343738 -284
rect 343806 -340 343862 -284
rect 343434 -464 343490 -408
rect 343558 -464 343614 -408
rect 343682 -464 343738 -408
rect 343806 -464 343862 -408
rect 343434 -588 343490 -532
rect 343558 -588 343614 -532
rect 343682 -588 343738 -532
rect 343806 -588 343862 -532
rect 371878 64294 371934 64350
rect 372002 64294 372058 64350
rect 371878 64170 371934 64226
rect 372002 64170 372058 64226
rect 371878 64046 371934 64102
rect 372002 64046 372058 64102
rect 371878 63922 371934 63978
rect 372002 63922 372058 63978
rect 356518 58294 356574 58350
rect 356642 58294 356698 58350
rect 356518 58170 356574 58226
rect 356642 58170 356698 58226
rect 356518 58046 356574 58102
rect 356642 58046 356698 58102
rect 356518 57922 356574 57978
rect 356642 57922 356698 57978
rect 374154 58294 374210 58350
rect 374278 58294 374334 58350
rect 374402 58294 374458 58350
rect 374526 58294 374582 58350
rect 374154 58170 374210 58226
rect 374278 58170 374334 58226
rect 374402 58170 374458 58226
rect 374526 58170 374582 58226
rect 374154 58046 374210 58102
rect 374278 58046 374334 58102
rect 374402 58046 374458 58102
rect 374526 58046 374582 58102
rect 374154 57922 374210 57978
rect 374278 57922 374334 57978
rect 374402 57922 374458 57978
rect 374526 57922 374582 57978
rect 349356 56222 349412 56278
rect 352716 56222 352772 56278
rect 347154 46294 347210 46350
rect 347278 46294 347334 46350
rect 347402 46294 347458 46350
rect 347526 46294 347582 46350
rect 347154 46170 347210 46226
rect 347278 46170 347334 46226
rect 347402 46170 347458 46226
rect 347526 46170 347582 46226
rect 347154 46046 347210 46102
rect 347278 46046 347334 46102
rect 347402 46046 347458 46102
rect 347526 46046 347582 46102
rect 347154 45922 347210 45978
rect 347278 45922 347334 45978
rect 347402 45922 347458 45978
rect 347526 45922 347582 45978
rect 371878 46294 371934 46350
rect 372002 46294 372058 46350
rect 371878 46170 371934 46226
rect 372002 46170 372058 46226
rect 371878 46046 371934 46102
rect 372002 46046 372058 46102
rect 371878 45922 371934 45978
rect 372002 45922 372058 45978
rect 356518 40294 356574 40350
rect 356642 40294 356698 40350
rect 356518 40170 356574 40226
rect 356642 40170 356698 40226
rect 356518 40046 356574 40102
rect 356642 40046 356698 40102
rect 356518 39922 356574 39978
rect 356642 39922 356698 39978
rect 374154 40294 374210 40350
rect 374278 40294 374334 40350
rect 374402 40294 374458 40350
rect 374526 40294 374582 40350
rect 374154 40170 374210 40226
rect 374278 40170 374334 40226
rect 374402 40170 374458 40226
rect 374526 40170 374582 40226
rect 374154 40046 374210 40102
rect 374278 40046 374334 40102
rect 374402 40046 374458 40102
rect 374526 40046 374582 40102
rect 374154 39922 374210 39978
rect 374278 39922 374334 39978
rect 374402 39922 374458 39978
rect 374526 39922 374582 39978
rect 347154 28294 347210 28350
rect 347278 28294 347334 28350
rect 347402 28294 347458 28350
rect 347526 28294 347582 28350
rect 347154 28170 347210 28226
rect 347278 28170 347334 28226
rect 347402 28170 347458 28226
rect 347526 28170 347582 28226
rect 347154 28046 347210 28102
rect 347278 28046 347334 28102
rect 347402 28046 347458 28102
rect 347526 28046 347582 28102
rect 347154 27922 347210 27978
rect 347278 27922 347334 27978
rect 347402 27922 347458 27978
rect 347526 27922 347582 27978
rect 347154 10294 347210 10350
rect 347278 10294 347334 10350
rect 347402 10294 347458 10350
rect 347526 10294 347582 10350
rect 347154 10170 347210 10226
rect 347278 10170 347334 10226
rect 347402 10170 347458 10226
rect 347526 10170 347582 10226
rect 347154 10046 347210 10102
rect 347278 10046 347334 10102
rect 347402 10046 347458 10102
rect 347526 10046 347582 10102
rect 347154 9922 347210 9978
rect 347278 9922 347334 9978
rect 347402 9922 347458 9978
rect 347526 9922 347582 9978
rect 347154 -1176 347210 -1120
rect 347278 -1176 347334 -1120
rect 347402 -1176 347458 -1120
rect 347526 -1176 347582 -1120
rect 347154 -1300 347210 -1244
rect 347278 -1300 347334 -1244
rect 347402 -1300 347458 -1244
rect 347526 -1300 347582 -1244
rect 347154 -1424 347210 -1368
rect 347278 -1424 347334 -1368
rect 347402 -1424 347458 -1368
rect 347526 -1424 347582 -1368
rect 347154 -1548 347210 -1492
rect 347278 -1548 347334 -1492
rect 347402 -1548 347458 -1492
rect 347526 -1548 347582 -1492
rect 374154 22294 374210 22350
rect 374278 22294 374334 22350
rect 374402 22294 374458 22350
rect 374526 22294 374582 22350
rect 374154 22170 374210 22226
rect 374278 22170 374334 22226
rect 374402 22170 374458 22226
rect 374526 22170 374582 22226
rect 374154 22046 374210 22102
rect 374278 22046 374334 22102
rect 374402 22046 374458 22102
rect 374526 22046 374582 22102
rect 374154 21922 374210 21978
rect 374278 21922 374334 21978
rect 374402 21922 374458 21978
rect 374526 21922 374582 21978
rect 374154 4294 374210 4350
rect 374278 4294 374334 4350
rect 374402 4294 374458 4350
rect 374526 4294 374582 4350
rect 374154 4170 374210 4226
rect 374278 4170 374334 4226
rect 374402 4170 374458 4226
rect 374526 4170 374582 4226
rect 374154 4046 374210 4102
rect 374278 4046 374334 4102
rect 374402 4046 374458 4102
rect 374526 4046 374582 4102
rect 374154 3922 374210 3978
rect 374278 3922 374334 3978
rect 374402 3922 374458 3978
rect 374526 3922 374582 3978
rect 374154 -216 374210 -160
rect 374278 -216 374334 -160
rect 374402 -216 374458 -160
rect 374526 -216 374582 -160
rect 374154 -340 374210 -284
rect 374278 -340 374334 -284
rect 374402 -340 374458 -284
rect 374526 -340 374582 -284
rect 374154 -464 374210 -408
rect 374278 -464 374334 -408
rect 374402 -464 374458 -408
rect 374526 -464 374582 -408
rect 374154 -588 374210 -532
rect 374278 -588 374334 -532
rect 374402 -588 374458 -532
rect 374526 -588 374582 -532
rect 400652 131282 400708 131338
rect 400652 125882 400708 125938
rect 404012 131102 404068 131158
rect 404874 130294 404930 130350
rect 404998 130294 405054 130350
rect 405122 130294 405178 130350
rect 405246 130294 405302 130350
rect 404874 130170 404930 130226
rect 404998 130170 405054 130226
rect 405122 130170 405178 130226
rect 405246 130170 405302 130226
rect 404874 130046 404930 130102
rect 404998 130046 405054 130102
rect 405122 130046 405178 130102
rect 405246 130046 405302 130102
rect 404874 129922 404930 129978
rect 404998 129922 405054 129978
rect 405122 129922 405178 129978
rect 405246 129922 405302 129978
rect 387238 112294 387294 112350
rect 387362 112294 387418 112350
rect 387238 112170 387294 112226
rect 387362 112170 387418 112226
rect 387238 112046 387294 112102
rect 387362 112046 387418 112102
rect 387238 111922 387294 111978
rect 387362 111922 387418 111978
rect 404874 112294 404930 112350
rect 404998 112294 405054 112350
rect 405122 112294 405178 112350
rect 405246 112294 405302 112350
rect 404874 112170 404930 112226
rect 404998 112170 405054 112226
rect 405122 112170 405178 112226
rect 405246 112170 405302 112226
rect 404874 112046 404930 112102
rect 404998 112046 405054 112102
rect 405122 112046 405178 112102
rect 405246 112046 405302 112102
rect 404874 111922 404930 111978
rect 404998 111922 405054 111978
rect 405122 111922 405178 111978
rect 405246 111922 405302 111978
rect 377874 100294 377930 100350
rect 377998 100294 378054 100350
rect 378122 100294 378178 100350
rect 378246 100294 378302 100350
rect 377874 100170 377930 100226
rect 377998 100170 378054 100226
rect 378122 100170 378178 100226
rect 378246 100170 378302 100226
rect 377874 100046 377930 100102
rect 377998 100046 378054 100102
rect 378122 100046 378178 100102
rect 378246 100046 378302 100102
rect 377874 99922 377930 99978
rect 377998 99922 378054 99978
rect 378122 99922 378178 99978
rect 378246 99922 378302 99978
rect 377874 82294 377930 82350
rect 377998 82294 378054 82350
rect 378122 82294 378178 82350
rect 378246 82294 378302 82350
rect 377874 82170 377930 82226
rect 377998 82170 378054 82226
rect 378122 82170 378178 82226
rect 378246 82170 378302 82226
rect 377874 82046 377930 82102
rect 377998 82046 378054 82102
rect 378122 82046 378178 82102
rect 378246 82046 378302 82102
rect 377874 81922 377930 81978
rect 377998 81922 378054 81978
rect 378122 81922 378178 81978
rect 378246 81922 378302 81978
rect 377874 64294 377930 64350
rect 377998 64294 378054 64350
rect 378122 64294 378178 64350
rect 378246 64294 378302 64350
rect 377874 64170 377930 64226
rect 377998 64170 378054 64226
rect 378122 64170 378178 64226
rect 378246 64170 378302 64226
rect 377874 64046 377930 64102
rect 377998 64046 378054 64102
rect 378122 64046 378178 64102
rect 378246 64046 378302 64102
rect 377874 63922 377930 63978
rect 377998 63922 378054 63978
rect 378122 63922 378178 63978
rect 378246 63922 378302 63978
rect 387238 58294 387294 58350
rect 387362 58294 387418 58350
rect 387238 58170 387294 58226
rect 387362 58170 387418 58226
rect 387238 58046 387294 58102
rect 387362 58046 387418 58102
rect 387238 57922 387294 57978
rect 387362 57922 387418 57978
rect 377874 46294 377930 46350
rect 377998 46294 378054 46350
rect 378122 46294 378178 46350
rect 378246 46294 378302 46350
rect 377874 46170 377930 46226
rect 377998 46170 378054 46226
rect 378122 46170 378178 46226
rect 378246 46170 378302 46226
rect 377874 46046 377930 46102
rect 377998 46046 378054 46102
rect 378122 46046 378178 46102
rect 378246 46046 378302 46102
rect 377874 45922 377930 45978
rect 377998 45922 378054 45978
rect 378122 45922 378178 45978
rect 378246 45922 378302 45978
rect 404874 94294 404930 94350
rect 404998 94294 405054 94350
rect 405122 94294 405178 94350
rect 405246 94294 405302 94350
rect 404874 94170 404930 94226
rect 404998 94170 405054 94226
rect 405122 94170 405178 94226
rect 405246 94170 405302 94226
rect 404874 94046 404930 94102
rect 404998 94046 405054 94102
rect 405122 94046 405178 94102
rect 405246 94046 405302 94102
rect 404874 93922 404930 93978
rect 404998 93922 405054 93978
rect 405122 93922 405178 93978
rect 405246 93922 405302 93978
rect 404874 76294 404930 76350
rect 404998 76294 405054 76350
rect 405122 76294 405178 76350
rect 405246 76294 405302 76350
rect 404874 76170 404930 76226
rect 404998 76170 405054 76226
rect 405122 76170 405178 76226
rect 405246 76170 405302 76226
rect 404874 76046 404930 76102
rect 404998 76046 405054 76102
rect 405122 76046 405178 76102
rect 405246 76046 405302 76102
rect 404874 75922 404930 75978
rect 404998 75922 405054 75978
rect 405122 75922 405178 75978
rect 405246 75922 405302 75978
rect 404874 58294 404930 58350
rect 404998 58294 405054 58350
rect 405122 58294 405178 58350
rect 405246 58294 405302 58350
rect 404874 58170 404930 58226
rect 404998 58170 405054 58226
rect 405122 58170 405178 58226
rect 405246 58170 405302 58226
rect 404874 58046 404930 58102
rect 404998 58046 405054 58102
rect 405122 58046 405178 58102
rect 405246 58046 405302 58102
rect 404874 57922 404930 57978
rect 404998 57922 405054 57978
rect 405122 57922 405178 57978
rect 405246 57922 405302 57978
rect 387238 40294 387294 40350
rect 387362 40294 387418 40350
rect 387238 40170 387294 40226
rect 387362 40170 387418 40226
rect 387238 40046 387294 40102
rect 387362 40046 387418 40102
rect 387238 39922 387294 39978
rect 387362 39922 387418 39978
rect 404874 40294 404930 40350
rect 404998 40294 405054 40350
rect 405122 40294 405178 40350
rect 405246 40294 405302 40350
rect 404874 40170 404930 40226
rect 404998 40170 405054 40226
rect 405122 40170 405178 40226
rect 405246 40170 405302 40226
rect 404874 40046 404930 40102
rect 404998 40046 405054 40102
rect 405122 40046 405178 40102
rect 405246 40046 405302 40102
rect 404874 39922 404930 39978
rect 404998 39922 405054 39978
rect 405122 39922 405178 39978
rect 405246 39922 405302 39978
rect 377874 28294 377930 28350
rect 377998 28294 378054 28350
rect 378122 28294 378178 28350
rect 378246 28294 378302 28350
rect 377874 28170 377930 28226
rect 377998 28170 378054 28226
rect 378122 28170 378178 28226
rect 378246 28170 378302 28226
rect 377874 28046 377930 28102
rect 377998 28046 378054 28102
rect 378122 28046 378178 28102
rect 378246 28046 378302 28102
rect 377874 27922 377930 27978
rect 377998 27922 378054 27978
rect 378122 27922 378178 27978
rect 378246 27922 378302 27978
rect 377874 10294 377930 10350
rect 377998 10294 378054 10350
rect 378122 10294 378178 10350
rect 378246 10294 378302 10350
rect 377874 10170 377930 10226
rect 377998 10170 378054 10226
rect 378122 10170 378178 10226
rect 378246 10170 378302 10226
rect 377874 10046 377930 10102
rect 377998 10046 378054 10102
rect 378122 10046 378178 10102
rect 378246 10046 378302 10102
rect 377874 9922 377930 9978
rect 377998 9922 378054 9978
rect 378122 9922 378178 9978
rect 378246 9922 378302 9978
rect 377874 -1176 377930 -1120
rect 377998 -1176 378054 -1120
rect 378122 -1176 378178 -1120
rect 378246 -1176 378302 -1120
rect 377874 -1300 377930 -1244
rect 377998 -1300 378054 -1244
rect 378122 -1300 378178 -1244
rect 378246 -1300 378302 -1244
rect 377874 -1424 377930 -1368
rect 377998 -1424 378054 -1368
rect 378122 -1424 378178 -1368
rect 378246 -1424 378302 -1368
rect 377874 -1548 377930 -1492
rect 377998 -1548 378054 -1492
rect 378122 -1548 378178 -1492
rect 378246 -1548 378302 -1492
rect 404874 22294 404930 22350
rect 404998 22294 405054 22350
rect 405122 22294 405178 22350
rect 405246 22294 405302 22350
rect 404874 22170 404930 22226
rect 404998 22170 405054 22226
rect 405122 22170 405178 22226
rect 405246 22170 405302 22226
rect 404874 22046 404930 22102
rect 404998 22046 405054 22102
rect 405122 22046 405178 22102
rect 405246 22046 405302 22102
rect 404874 21922 404930 21978
rect 404998 21922 405054 21978
rect 405122 21922 405178 21978
rect 405246 21922 405302 21978
rect 404874 4294 404930 4350
rect 404998 4294 405054 4350
rect 405122 4294 405178 4350
rect 405246 4294 405302 4350
rect 404874 4170 404930 4226
rect 404998 4170 405054 4226
rect 405122 4170 405178 4226
rect 405246 4170 405302 4226
rect 404874 4046 404930 4102
rect 404998 4046 405054 4102
rect 405122 4046 405178 4102
rect 405246 4046 405302 4102
rect 404874 3922 404930 3978
rect 404998 3922 405054 3978
rect 405122 3922 405178 3978
rect 405246 3922 405302 3978
rect 404874 -216 404930 -160
rect 404998 -216 405054 -160
rect 405122 -216 405178 -160
rect 405246 -216 405302 -160
rect 404874 -340 404930 -284
rect 404998 -340 405054 -284
rect 405122 -340 405178 -284
rect 405246 -340 405302 -284
rect 404874 -464 404930 -408
rect 404998 -464 405054 -408
rect 405122 -464 405178 -408
rect 405246 -464 405302 -408
rect 404874 -588 404930 -532
rect 404998 -588 405054 -532
rect 405122 -588 405178 -532
rect 405246 -588 405302 -532
rect 435594 220294 435650 220350
rect 435718 220294 435774 220350
rect 435842 220294 435898 220350
rect 435966 220294 436022 220350
rect 435594 220170 435650 220226
rect 435718 220170 435774 220226
rect 435842 220170 435898 220226
rect 435966 220170 436022 220226
rect 435594 220046 435650 220102
rect 435718 220046 435774 220102
rect 435842 220046 435898 220102
rect 435966 220046 436022 220102
rect 435594 219922 435650 219978
rect 435718 219922 435774 219978
rect 435842 219922 435898 219978
rect 435966 219922 436022 219978
rect 433878 208294 433934 208350
rect 434002 208294 434058 208350
rect 433878 208170 433934 208226
rect 434002 208170 434058 208226
rect 433878 208046 433934 208102
rect 434002 208046 434058 208102
rect 433878 207922 433934 207978
rect 434002 207922 434058 207978
rect 418518 202294 418574 202350
rect 418642 202294 418698 202350
rect 418518 202170 418574 202226
rect 418642 202170 418698 202226
rect 418518 202046 418574 202102
rect 418642 202046 418698 202102
rect 418518 201922 418574 201978
rect 418642 201922 418698 201978
rect 435594 202294 435650 202350
rect 435718 202294 435774 202350
rect 435842 202294 435898 202350
rect 435966 202294 436022 202350
rect 435594 202170 435650 202226
rect 435718 202170 435774 202226
rect 435842 202170 435898 202226
rect 435966 202170 436022 202226
rect 435594 202046 435650 202102
rect 435718 202046 435774 202102
rect 435842 202046 435898 202102
rect 435966 202046 436022 202102
rect 435594 201922 435650 201978
rect 435718 201922 435774 201978
rect 435842 201922 435898 201978
rect 435966 201922 436022 201978
rect 414652 198242 414708 198298
rect 411180 195188 411236 195238
rect 411180 195182 411236 195188
rect 411292 192482 411348 192538
rect 411180 192302 411236 192358
rect 408594 190294 408650 190350
rect 408718 190294 408774 190350
rect 408842 190294 408898 190350
rect 408966 190294 409022 190350
rect 408594 190170 408650 190226
rect 408718 190170 408774 190226
rect 408842 190170 408898 190226
rect 408966 190170 409022 190226
rect 408594 190046 408650 190102
rect 408718 190046 408774 190102
rect 408842 190046 408898 190102
rect 408966 190046 409022 190102
rect 408594 189922 408650 189978
rect 408718 189922 408774 189978
rect 408842 189922 408898 189978
rect 408966 189922 409022 189978
rect 433878 190294 433934 190350
rect 434002 190294 434058 190350
rect 433878 190170 433934 190226
rect 434002 190170 434058 190226
rect 433878 190046 433934 190102
rect 434002 190046 434058 190102
rect 433878 189922 433934 189978
rect 434002 189922 434058 189978
rect 418518 184294 418574 184350
rect 418642 184294 418698 184350
rect 418518 184170 418574 184226
rect 418642 184170 418698 184226
rect 418518 184046 418574 184102
rect 418642 184046 418698 184102
rect 418518 183922 418574 183978
rect 418642 183922 418698 183978
rect 435594 184294 435650 184350
rect 435718 184294 435774 184350
rect 435842 184294 435898 184350
rect 435966 184294 436022 184350
rect 435594 184170 435650 184226
rect 435718 184170 435774 184226
rect 435842 184170 435898 184226
rect 435966 184170 436022 184226
rect 435594 184046 435650 184102
rect 435718 184046 435774 184102
rect 435842 184046 435898 184102
rect 435966 184046 436022 184102
rect 435594 183922 435650 183978
rect 435718 183922 435774 183978
rect 435842 183922 435898 183978
rect 435966 183922 436022 183978
rect 408594 172294 408650 172350
rect 408718 172294 408774 172350
rect 408842 172294 408898 172350
rect 408966 172294 409022 172350
rect 408594 172170 408650 172226
rect 408718 172170 408774 172226
rect 408842 172170 408898 172226
rect 408966 172170 409022 172226
rect 408594 172046 408650 172102
rect 408718 172046 408774 172102
rect 408842 172046 408898 172102
rect 408966 172046 409022 172102
rect 408594 171922 408650 171978
rect 408718 171922 408774 171978
rect 408842 171922 408898 171978
rect 408966 171922 409022 171978
rect 435594 166294 435650 166350
rect 435718 166294 435774 166350
rect 435842 166294 435898 166350
rect 435966 166294 436022 166350
rect 435594 166170 435650 166226
rect 435718 166170 435774 166226
rect 435842 166170 435898 166226
rect 435966 166170 436022 166226
rect 435594 166046 435650 166102
rect 435718 166046 435774 166102
rect 435842 166046 435898 166102
rect 435966 166046 436022 166102
rect 435594 165922 435650 165978
rect 435718 165922 435774 165978
rect 435842 165922 435898 165978
rect 435966 165922 436022 165978
rect 408594 154294 408650 154350
rect 408718 154294 408774 154350
rect 408842 154294 408898 154350
rect 408966 154294 409022 154350
rect 408594 154170 408650 154226
rect 408718 154170 408774 154226
rect 408842 154170 408898 154226
rect 408966 154170 409022 154226
rect 408594 154046 408650 154102
rect 408718 154046 408774 154102
rect 408842 154046 408898 154102
rect 408966 154046 409022 154102
rect 408594 153922 408650 153978
rect 408718 153922 408774 153978
rect 408842 153922 408898 153978
rect 408966 153922 409022 153978
rect 408594 136294 408650 136350
rect 408718 136294 408774 136350
rect 408842 136294 408898 136350
rect 408966 136294 409022 136350
rect 408594 136170 408650 136226
rect 408718 136170 408774 136226
rect 408842 136170 408898 136226
rect 408966 136170 409022 136226
rect 408594 136046 408650 136102
rect 408718 136046 408774 136102
rect 408842 136046 408898 136102
rect 408966 136046 409022 136102
rect 408594 135922 408650 135978
rect 408718 135922 408774 135978
rect 408842 135922 408898 135978
rect 408966 135922 409022 135978
rect 408594 118294 408650 118350
rect 408718 118294 408774 118350
rect 408842 118294 408898 118350
rect 408966 118294 409022 118350
rect 408594 118170 408650 118226
rect 408718 118170 408774 118226
rect 408842 118170 408898 118226
rect 408966 118170 409022 118226
rect 408594 118046 408650 118102
rect 408718 118046 408774 118102
rect 408842 118046 408898 118102
rect 408966 118046 409022 118102
rect 408594 117922 408650 117978
rect 408718 117922 408774 117978
rect 408842 117922 408898 117978
rect 408966 117922 409022 117978
rect 435594 148294 435650 148350
rect 435718 148294 435774 148350
rect 435842 148294 435898 148350
rect 435966 148294 436022 148350
rect 435594 148170 435650 148226
rect 435718 148170 435774 148226
rect 435842 148170 435898 148226
rect 435966 148170 436022 148226
rect 435594 148046 435650 148102
rect 435718 148046 435774 148102
rect 435842 148046 435898 148102
rect 435966 148046 436022 148102
rect 435594 147922 435650 147978
rect 435718 147922 435774 147978
rect 435842 147922 435898 147978
rect 435966 147922 436022 147978
rect 433878 136294 433934 136350
rect 434002 136294 434058 136350
rect 433878 136170 433934 136226
rect 434002 136170 434058 136226
rect 433878 136046 433934 136102
rect 434002 136046 434058 136102
rect 433878 135922 433934 135978
rect 434002 135922 434058 135978
rect 418518 130294 418574 130350
rect 418642 130294 418698 130350
rect 418518 130170 418574 130226
rect 418642 130170 418698 130226
rect 418518 130046 418574 130102
rect 418642 130046 418698 130102
rect 418518 129922 418574 129978
rect 418642 129922 418698 129978
rect 435594 130294 435650 130350
rect 435718 130294 435774 130350
rect 435842 130294 435898 130350
rect 435966 130294 436022 130350
rect 435594 130170 435650 130226
rect 435718 130170 435774 130226
rect 435842 130170 435898 130226
rect 435966 130170 436022 130226
rect 435594 130046 435650 130102
rect 435718 130046 435774 130102
rect 435842 130046 435898 130102
rect 435966 130046 436022 130102
rect 435594 129922 435650 129978
rect 435718 129922 435774 129978
rect 435842 129922 435898 129978
rect 435966 129922 436022 129978
rect 411516 128402 411572 128458
rect 411180 122462 411236 122518
rect 449238 400294 449294 400350
rect 449362 400294 449418 400350
rect 449238 400170 449294 400226
rect 449362 400170 449418 400226
rect 449238 400046 449294 400102
rect 449362 400046 449418 400102
rect 449238 399922 449294 399978
rect 449362 399922 449418 399978
rect 439314 388294 439370 388350
rect 439438 388294 439494 388350
rect 439562 388294 439618 388350
rect 439686 388294 439742 388350
rect 439314 388170 439370 388226
rect 439438 388170 439494 388226
rect 439562 388170 439618 388226
rect 439686 388170 439742 388226
rect 439314 388046 439370 388102
rect 439438 388046 439494 388102
rect 439562 388046 439618 388102
rect 439686 388046 439742 388102
rect 439314 387922 439370 387978
rect 439438 387922 439494 387978
rect 439562 387922 439618 387978
rect 439686 387922 439742 387978
rect 439314 370294 439370 370350
rect 439438 370294 439494 370350
rect 439562 370294 439618 370350
rect 439686 370294 439742 370350
rect 439314 370170 439370 370226
rect 439438 370170 439494 370226
rect 439562 370170 439618 370226
rect 439686 370170 439742 370226
rect 439314 370046 439370 370102
rect 439438 370046 439494 370102
rect 439562 370046 439618 370102
rect 439686 370046 439742 370102
rect 439314 369922 439370 369978
rect 439438 369922 439494 369978
rect 439562 369922 439618 369978
rect 439686 369922 439742 369978
rect 455532 394622 455588 394678
rect 455532 391562 455588 391618
rect 456988 396422 457044 396478
rect 458668 398942 458724 398998
rect 458892 397322 458948 397378
rect 461132 403082 461188 403138
rect 470034 424294 470090 424350
rect 470158 424294 470214 424350
rect 470282 424294 470338 424350
rect 470406 424294 470462 424350
rect 470034 424170 470090 424226
rect 470158 424170 470214 424226
rect 470282 424170 470338 424226
rect 470406 424170 470462 424226
rect 470034 424046 470090 424102
rect 470158 424046 470214 424102
rect 470282 424046 470338 424102
rect 470406 424046 470462 424102
rect 470034 423922 470090 423978
rect 470158 423922 470214 423978
rect 470282 423922 470338 423978
rect 470406 423922 470462 423978
rect 466314 400294 466370 400350
rect 466438 400294 466494 400350
rect 466562 400294 466618 400350
rect 466686 400294 466742 400350
rect 466314 400170 466370 400226
rect 466438 400170 466494 400226
rect 466562 400170 466618 400226
rect 466686 400170 466742 400226
rect 466314 400046 466370 400102
rect 466438 400046 466494 400102
rect 466562 400046 466618 400102
rect 466686 400046 466742 400102
rect 466314 399922 466370 399978
rect 466438 399922 466494 399978
rect 466562 399922 466618 399978
rect 466686 399922 466742 399978
rect 466314 382294 466370 382350
rect 466438 382294 466494 382350
rect 466562 382294 466618 382350
rect 466686 382294 466742 382350
rect 466314 382170 466370 382226
rect 466438 382170 466494 382226
rect 466562 382170 466618 382226
rect 466686 382170 466742 382226
rect 466314 382046 466370 382102
rect 466438 382046 466494 382102
rect 466562 382046 466618 382102
rect 466686 382046 466742 382102
rect 466314 381922 466370 381978
rect 466438 381922 466494 381978
rect 466562 381922 466618 381978
rect 466686 381922 466742 381978
rect 439314 352294 439370 352350
rect 439438 352294 439494 352350
rect 439562 352294 439618 352350
rect 439686 352294 439742 352350
rect 439314 352170 439370 352226
rect 439438 352170 439494 352226
rect 439562 352170 439618 352226
rect 439686 352170 439742 352226
rect 439314 352046 439370 352102
rect 439438 352046 439494 352102
rect 439562 352046 439618 352102
rect 439686 352046 439742 352102
rect 439314 351922 439370 351978
rect 439438 351922 439494 351978
rect 439562 351922 439618 351978
rect 439686 351922 439742 351978
rect 497034 436294 497090 436350
rect 497158 436294 497214 436350
rect 497282 436294 497338 436350
rect 497406 436294 497462 436350
rect 497034 436170 497090 436226
rect 497158 436170 497214 436226
rect 497282 436170 497338 436226
rect 497406 436170 497462 436226
rect 497034 436046 497090 436102
rect 497158 436046 497214 436102
rect 497282 436046 497338 436102
rect 497406 436046 497462 436102
rect 497034 435922 497090 435978
rect 497158 435922 497214 435978
rect 497282 435922 497338 435978
rect 497406 435922 497462 435978
rect 472108 420002 472164 420058
rect 480518 418294 480574 418350
rect 480642 418294 480698 418350
rect 480518 418170 480574 418226
rect 480642 418170 480698 418226
rect 480518 418046 480574 418102
rect 480642 418046 480698 418102
rect 480518 417922 480574 417978
rect 480642 417922 480698 417978
rect 497034 418294 497090 418350
rect 497158 418294 497214 418350
rect 497282 418294 497338 418350
rect 497406 418294 497462 418350
rect 497034 418170 497090 418226
rect 497158 418170 497214 418226
rect 497282 418170 497338 418226
rect 497406 418170 497462 418226
rect 497034 418046 497090 418102
rect 497158 418046 497214 418102
rect 497282 418046 497338 418102
rect 497406 418046 497462 418102
rect 497034 417922 497090 417978
rect 497158 417922 497214 417978
rect 497282 417922 497338 417978
rect 497406 417922 497462 417978
rect 472108 413342 472164 413398
rect 472108 412132 472164 412138
rect 472108 412082 472164 412132
rect 470034 406294 470090 406350
rect 470158 406294 470214 406350
rect 470282 406294 470338 406350
rect 470406 406294 470462 406350
rect 470034 406170 470090 406226
rect 470158 406170 470214 406226
rect 470282 406170 470338 406226
rect 470406 406170 470462 406226
rect 470034 406046 470090 406102
rect 470158 406046 470214 406102
rect 470282 406046 470338 406102
rect 470406 406046 470462 406102
rect 470034 405922 470090 405978
rect 470158 405922 470214 405978
rect 470282 405922 470338 405978
rect 470406 405922 470462 405978
rect 472108 404702 472164 404758
rect 470034 388294 470090 388350
rect 470158 388294 470214 388350
rect 470282 388294 470338 388350
rect 470406 388294 470462 388350
rect 470034 388170 470090 388226
rect 470158 388170 470214 388226
rect 470282 388170 470338 388226
rect 470406 388170 470462 388226
rect 470034 388046 470090 388102
rect 470158 388046 470214 388102
rect 470282 388046 470338 388102
rect 470406 388046 470462 388102
rect 470034 387922 470090 387978
rect 470158 387922 470214 387978
rect 470282 387922 470338 387978
rect 470406 387922 470462 387978
rect 466314 364294 466370 364350
rect 466438 364294 466494 364350
rect 466562 364294 466618 364350
rect 466686 364294 466742 364350
rect 466314 364170 466370 364226
rect 466438 364170 466494 364226
rect 466562 364170 466618 364226
rect 466686 364170 466742 364226
rect 466314 364046 466370 364102
rect 466438 364046 466494 364102
rect 466562 364046 466618 364102
rect 466686 364046 466742 364102
rect 466314 363922 466370 363978
rect 466438 363922 466494 363978
rect 466562 363922 466618 363978
rect 466686 363922 466742 363978
rect 449238 346294 449294 346350
rect 449362 346294 449418 346350
rect 449238 346170 449294 346226
rect 449362 346170 449418 346226
rect 449238 346046 449294 346102
rect 449362 346046 449418 346102
rect 449238 345922 449294 345978
rect 449362 345922 449418 345978
rect 466314 346294 466370 346350
rect 466438 346294 466494 346350
rect 466562 346294 466618 346350
rect 466686 346294 466742 346350
rect 466314 346170 466370 346226
rect 466438 346170 466494 346226
rect 466562 346170 466618 346226
rect 466686 346170 466742 346226
rect 466314 346046 466370 346102
rect 466438 346046 466494 346102
rect 466562 346046 466618 346102
rect 466686 346046 466742 346102
rect 466314 345922 466370 345978
rect 466438 345922 466494 345978
rect 466562 345922 466618 345978
rect 466686 345922 466742 345978
rect 460236 344402 460292 344458
rect 460236 340082 460292 340138
rect 461132 341342 461188 341398
rect 455420 339722 455476 339778
rect 455420 339362 455476 339418
rect 455308 337742 455364 337798
rect 455532 338822 455588 338878
rect 455308 337022 455364 337078
rect 455644 336482 455700 336538
rect 439314 334294 439370 334350
rect 439438 334294 439494 334350
rect 439562 334294 439618 334350
rect 439686 334294 439742 334350
rect 439314 334170 439370 334226
rect 439438 334170 439494 334226
rect 439562 334170 439618 334226
rect 439686 334170 439742 334226
rect 439314 334046 439370 334102
rect 439438 334046 439494 334102
rect 439562 334046 439618 334102
rect 439686 334046 439742 334102
rect 439314 333922 439370 333978
rect 439438 333922 439494 333978
rect 439562 333922 439618 333978
rect 439686 333922 439742 333978
rect 455308 334682 455364 334738
rect 455532 331802 455588 331858
rect 455308 330902 455364 330958
rect 455420 329822 455476 329878
rect 449238 328294 449294 328350
rect 449362 328294 449418 328350
rect 449238 328170 449294 328226
rect 449362 328170 449418 328226
rect 449238 328046 449294 328102
rect 449362 328046 449418 328102
rect 449238 327922 449294 327978
rect 449362 327922 449418 327978
rect 439314 316294 439370 316350
rect 439438 316294 439494 316350
rect 439562 316294 439618 316350
rect 439686 316294 439742 316350
rect 439314 316170 439370 316226
rect 439438 316170 439494 316226
rect 439562 316170 439618 316226
rect 439686 316170 439742 316226
rect 439314 316046 439370 316102
rect 439438 316046 439494 316102
rect 439562 316046 439618 316102
rect 439686 316046 439742 316102
rect 439314 315922 439370 315978
rect 439438 315922 439494 315978
rect 439562 315922 439618 315978
rect 439686 315922 439742 315978
rect 461132 339182 461188 339238
rect 460236 324962 460292 325018
rect 460236 322442 460292 322498
rect 464492 331082 464548 331138
rect 462812 330002 462868 330058
rect 462812 325862 462868 325918
rect 464492 323882 464548 323938
rect 466314 328294 466370 328350
rect 466438 328294 466494 328350
rect 466562 328294 466618 328350
rect 466686 328294 466742 328350
rect 466314 328170 466370 328226
rect 466438 328170 466494 328226
rect 466562 328170 466618 328226
rect 466686 328170 466742 328226
rect 466314 328046 466370 328102
rect 466438 328046 466494 328102
rect 466562 328046 466618 328102
rect 466686 328046 466742 328102
rect 466314 327922 466370 327978
rect 466438 327922 466494 327978
rect 466562 327922 466618 327978
rect 466686 327922 466742 327978
rect 461132 319022 461188 319078
rect 466314 310294 466370 310350
rect 466438 310294 466494 310350
rect 466562 310294 466618 310350
rect 466686 310294 466742 310350
rect 466314 310170 466370 310226
rect 466438 310170 466494 310226
rect 466562 310170 466618 310226
rect 466686 310170 466742 310226
rect 466314 310046 466370 310102
rect 466438 310046 466494 310102
rect 466562 310046 466618 310102
rect 466686 310046 466742 310102
rect 466314 309922 466370 309978
rect 466438 309922 466494 309978
rect 466562 309922 466618 309978
rect 466686 309922 466742 309978
rect 439314 298294 439370 298350
rect 439438 298294 439494 298350
rect 439562 298294 439618 298350
rect 439686 298294 439742 298350
rect 439314 298170 439370 298226
rect 439438 298170 439494 298226
rect 439562 298170 439618 298226
rect 439686 298170 439742 298226
rect 439314 298046 439370 298102
rect 439438 298046 439494 298102
rect 439562 298046 439618 298102
rect 439686 298046 439742 298102
rect 439314 297922 439370 297978
rect 439438 297922 439494 297978
rect 439562 297922 439618 297978
rect 439686 297922 439742 297978
rect 466314 292294 466370 292350
rect 466438 292294 466494 292350
rect 466562 292294 466618 292350
rect 466686 292294 466742 292350
rect 466314 292170 466370 292226
rect 466438 292170 466494 292226
rect 466562 292170 466618 292226
rect 466686 292170 466742 292226
rect 466314 292046 466370 292102
rect 466438 292046 466494 292102
rect 466562 292046 466618 292102
rect 466686 292046 466742 292102
rect 466314 291922 466370 291978
rect 466438 291922 466494 291978
rect 466562 291922 466618 291978
rect 466686 291922 466742 291978
rect 439314 280294 439370 280350
rect 439438 280294 439494 280350
rect 439562 280294 439618 280350
rect 439686 280294 439742 280350
rect 439314 280170 439370 280226
rect 439438 280170 439494 280226
rect 439562 280170 439618 280226
rect 439686 280170 439742 280226
rect 439314 280046 439370 280102
rect 439438 280046 439494 280102
rect 439562 280046 439618 280102
rect 439686 280046 439742 280102
rect 439314 279922 439370 279978
rect 439438 279922 439494 279978
rect 439562 279922 439618 279978
rect 439686 279922 439742 279978
rect 455420 277982 455476 278038
rect 455308 277116 455364 277138
rect 455308 277082 455364 277116
rect 449238 274294 449294 274350
rect 449362 274294 449418 274350
rect 449238 274170 449294 274226
rect 449362 274170 449418 274226
rect 449238 274046 449294 274102
rect 449362 274046 449418 274102
rect 449238 273922 449294 273978
rect 449362 273922 449418 273978
rect 455532 270962 455588 271018
rect 439314 262294 439370 262350
rect 439438 262294 439494 262350
rect 439562 262294 439618 262350
rect 439686 262294 439742 262350
rect 439314 262170 439370 262226
rect 439438 262170 439494 262226
rect 439562 262170 439618 262226
rect 439686 262170 439742 262226
rect 439314 262046 439370 262102
rect 439438 262046 439494 262102
rect 439562 262046 439618 262102
rect 439686 262046 439742 262102
rect 439314 261922 439370 261978
rect 439438 261922 439494 261978
rect 439562 261922 439618 261978
rect 439686 261922 439742 261978
rect 456876 258182 456932 258238
rect 449238 256294 449294 256350
rect 449362 256294 449418 256350
rect 449238 256170 449294 256226
rect 449362 256170 449418 256226
rect 449238 256046 449294 256102
rect 449362 256046 449418 256102
rect 449238 255922 449294 255978
rect 449362 255922 449418 255978
rect 457100 253502 457156 253558
rect 466314 274294 466370 274350
rect 466438 274294 466494 274350
rect 466562 274294 466618 274350
rect 466686 274294 466742 274350
rect 466314 274170 466370 274226
rect 466438 274170 466494 274226
rect 466562 274170 466618 274226
rect 466686 274170 466742 274226
rect 466314 274046 466370 274102
rect 466438 274046 466494 274102
rect 466562 274046 466618 274102
rect 466686 274046 466742 274102
rect 466314 273922 466370 273978
rect 466438 273922 466494 273978
rect 466562 273922 466618 273978
rect 466686 273922 466742 273978
rect 457212 251882 457268 251938
rect 464492 255302 464548 255358
rect 495878 406294 495934 406350
rect 496002 406294 496058 406350
rect 495878 406170 495934 406226
rect 496002 406170 496058 406226
rect 495878 406046 495934 406102
rect 496002 406046 496058 406102
rect 495878 405922 495934 405978
rect 496002 405922 496058 405978
rect 480518 400294 480574 400350
rect 480642 400294 480698 400350
rect 480518 400170 480574 400226
rect 480642 400170 480698 400226
rect 480518 400046 480574 400102
rect 480642 400046 480698 400102
rect 480518 399922 480574 399978
rect 480642 399922 480698 399978
rect 511238 472294 511294 472350
rect 511362 472294 511418 472350
rect 511238 472170 511294 472226
rect 511362 472170 511418 472226
rect 511238 472046 511294 472102
rect 511362 472046 511418 472102
rect 511238 471922 511294 471978
rect 511362 471922 511418 471978
rect 500754 460294 500810 460350
rect 500878 460294 500934 460350
rect 501002 460294 501058 460350
rect 501126 460294 501182 460350
rect 500754 460170 500810 460226
rect 500878 460170 500934 460226
rect 501002 460170 501058 460226
rect 501126 460170 501182 460226
rect 500754 460046 500810 460102
rect 500878 460046 500934 460102
rect 501002 460046 501058 460102
rect 501126 460046 501182 460102
rect 500754 459922 500810 459978
rect 500878 459922 500934 459978
rect 501002 459922 501058 459978
rect 501126 459922 501182 459978
rect 500754 442294 500810 442350
rect 500878 442294 500934 442350
rect 501002 442294 501058 442350
rect 501126 442294 501182 442350
rect 500754 442170 500810 442226
rect 500878 442170 500934 442226
rect 501002 442170 501058 442226
rect 501126 442170 501182 442226
rect 500754 442046 500810 442102
rect 500878 442046 500934 442102
rect 501002 442046 501058 442102
rect 501126 442046 501182 442102
rect 500754 441922 500810 441978
rect 500878 441922 500934 441978
rect 501002 441922 501058 441978
rect 501126 441922 501182 441978
rect 521052 466082 521108 466138
rect 527754 472294 527810 472350
rect 527878 472294 527934 472350
rect 528002 472294 528058 472350
rect 528126 472294 528182 472350
rect 527754 472170 527810 472226
rect 527878 472170 527934 472226
rect 528002 472170 528058 472226
rect 528126 472170 528182 472226
rect 527754 472046 527810 472102
rect 527878 472046 527934 472102
rect 528002 472046 528058 472102
rect 528126 472046 528182 472102
rect 527754 471922 527810 471978
rect 527878 471922 527934 471978
rect 528002 471922 528058 471978
rect 528126 471922 528182 471978
rect 527754 454294 527810 454350
rect 527878 454294 527934 454350
rect 528002 454294 528058 454350
rect 528126 454294 528182 454350
rect 527754 454170 527810 454226
rect 527878 454170 527934 454226
rect 528002 454170 528058 454226
rect 528126 454170 528182 454226
rect 527754 454046 527810 454102
rect 527878 454046 527934 454102
rect 528002 454046 528058 454102
rect 528126 454046 528182 454102
rect 527754 453922 527810 453978
rect 527878 453922 527934 453978
rect 528002 453922 528058 453978
rect 528126 453922 528182 453978
rect 527754 436294 527810 436350
rect 527878 436294 527934 436350
rect 528002 436294 528058 436350
rect 528126 436294 528182 436350
rect 527754 436170 527810 436226
rect 527878 436170 527934 436226
rect 528002 436170 528058 436226
rect 528126 436170 528182 436226
rect 527754 436046 527810 436102
rect 527878 436046 527934 436102
rect 528002 436046 528058 436102
rect 528126 436046 528182 436102
rect 527754 435922 527810 435978
rect 527878 435922 527934 435978
rect 528002 435922 528058 435978
rect 528126 435922 528182 435978
rect 500754 424294 500810 424350
rect 500878 424294 500934 424350
rect 501002 424294 501058 424350
rect 501126 424294 501182 424350
rect 500754 424170 500810 424226
rect 500878 424170 500934 424226
rect 501002 424170 501058 424226
rect 501126 424170 501182 424226
rect 500754 424046 500810 424102
rect 500878 424046 500934 424102
rect 501002 424046 501058 424102
rect 501126 424046 501182 424102
rect 500754 423922 500810 423978
rect 500878 423922 500934 423978
rect 501002 423922 501058 423978
rect 501126 423922 501182 423978
rect 511238 418294 511294 418350
rect 511362 418294 511418 418350
rect 511238 418170 511294 418226
rect 511362 418170 511418 418226
rect 511238 418046 511294 418102
rect 511362 418046 511418 418102
rect 511238 417922 511294 417978
rect 511362 417922 511418 417978
rect 527754 418294 527810 418350
rect 527878 418294 527934 418350
rect 528002 418294 528058 418350
rect 528126 418294 528182 418350
rect 527754 418170 527810 418226
rect 527878 418170 527934 418226
rect 528002 418170 528058 418226
rect 528126 418170 528182 418226
rect 527754 418046 527810 418102
rect 527878 418046 527934 418102
rect 528002 418046 528058 418102
rect 528126 418046 528182 418102
rect 527754 417922 527810 417978
rect 527878 417922 527934 417978
rect 528002 417922 528058 417978
rect 528126 417922 528182 417978
rect 523292 414962 523348 415018
rect 518252 413522 518308 413578
rect 518252 403982 518308 404038
rect 497034 400294 497090 400350
rect 497158 400294 497214 400350
rect 497282 400294 497338 400350
rect 497406 400294 497462 400350
rect 497034 400170 497090 400226
rect 497158 400170 497214 400226
rect 497282 400170 497338 400226
rect 497406 400170 497462 400226
rect 497034 400046 497090 400102
rect 497158 400046 497214 400102
rect 497282 400046 497338 400102
rect 497406 400046 497462 400102
rect 497034 399922 497090 399978
rect 497158 399922 497214 399978
rect 497282 399922 497338 399978
rect 497406 399922 497462 399978
rect 495836 388333 495892 388389
rect 495940 388333 495996 388389
rect 496044 388333 496100 388389
rect 497034 382294 497090 382350
rect 497158 382294 497214 382350
rect 497282 382294 497338 382350
rect 497406 382294 497462 382350
rect 497034 382170 497090 382226
rect 497158 382170 497214 382226
rect 497282 382170 497338 382226
rect 497406 382170 497462 382226
rect 497034 382046 497090 382102
rect 497158 382046 497214 382102
rect 497282 382046 497338 382102
rect 497406 382046 497462 382102
rect 497034 381922 497090 381978
rect 497158 381922 497214 381978
rect 497282 381922 497338 381978
rect 497406 381922 497462 381978
rect 470034 370294 470090 370350
rect 470158 370294 470214 370350
rect 470282 370294 470338 370350
rect 470406 370294 470462 370350
rect 470034 370170 470090 370226
rect 470158 370170 470214 370226
rect 470282 370170 470338 370226
rect 470406 370170 470462 370226
rect 470034 370046 470090 370102
rect 470158 370046 470214 370102
rect 470282 370046 470338 370102
rect 470406 370046 470462 370102
rect 470034 369922 470090 369978
rect 470158 369922 470214 369978
rect 470282 369922 470338 369978
rect 470406 369922 470462 369978
rect 497034 364294 497090 364350
rect 497158 364294 497214 364350
rect 497282 364294 497338 364350
rect 497406 364294 497462 364350
rect 497034 364170 497090 364226
rect 497158 364170 497214 364226
rect 497282 364170 497338 364226
rect 497406 364170 497462 364226
rect 497034 364046 497090 364102
rect 497158 364046 497214 364102
rect 497282 364046 497338 364102
rect 497406 364046 497462 364102
rect 497034 363922 497090 363978
rect 497158 363922 497214 363978
rect 497282 363922 497338 363978
rect 497406 363922 497462 363978
rect 470034 352294 470090 352350
rect 470158 352294 470214 352350
rect 470282 352294 470338 352350
rect 470406 352294 470462 352350
rect 470034 352170 470090 352226
rect 470158 352170 470214 352226
rect 470282 352170 470338 352226
rect 470406 352170 470462 352226
rect 470034 352046 470090 352102
rect 470158 352046 470214 352102
rect 470282 352046 470338 352102
rect 470406 352046 470462 352102
rect 470034 351922 470090 351978
rect 470158 351922 470214 351978
rect 470282 351922 470338 351978
rect 470406 351922 470462 351978
rect 495878 352294 495934 352350
rect 496002 352294 496058 352350
rect 495878 352170 495934 352226
rect 496002 352170 496058 352226
rect 495878 352046 495934 352102
rect 496002 352046 496058 352102
rect 495878 351922 495934 351978
rect 496002 351922 496058 351978
rect 473228 348542 473284 348598
rect 480518 346294 480574 346350
rect 480642 346294 480698 346350
rect 480518 346170 480574 346226
rect 480642 346170 480698 346226
rect 480518 346046 480574 346102
rect 480642 346046 480698 346102
rect 480518 345922 480574 345978
rect 480642 345922 480698 345978
rect 497034 346294 497090 346350
rect 497158 346294 497214 346350
rect 497282 346294 497338 346350
rect 497406 346294 497462 346350
rect 497034 346170 497090 346226
rect 497158 346170 497214 346226
rect 497282 346170 497338 346226
rect 497406 346170 497462 346226
rect 497034 346046 497090 346102
rect 497158 346046 497214 346102
rect 497282 346046 497338 346102
rect 497406 346046 497462 346102
rect 497034 345922 497090 345978
rect 497158 345922 497214 345978
rect 497282 345922 497338 345978
rect 497406 345922 497462 345978
rect 476028 341702 476084 341758
rect 473676 341162 473732 341218
rect 470034 334294 470090 334350
rect 470158 334294 470214 334350
rect 470282 334294 470338 334350
rect 470406 334294 470462 334350
rect 470034 334170 470090 334226
rect 470158 334170 470214 334226
rect 470282 334170 470338 334226
rect 470406 334170 470462 334226
rect 470034 334046 470090 334102
rect 470158 334046 470214 334102
rect 470282 334046 470338 334102
rect 470406 334046 470462 334102
rect 470034 333922 470090 333978
rect 470158 333922 470214 333978
rect 470282 333922 470338 333978
rect 470406 333922 470462 333978
rect 517244 403262 517300 403318
rect 511238 400294 511294 400350
rect 511362 400294 511418 400350
rect 511238 400170 511294 400226
rect 511362 400170 511418 400226
rect 511238 400046 511294 400102
rect 511362 400046 511418 400102
rect 511238 399922 511294 399978
rect 511362 399922 511418 399978
rect 500754 388294 500810 388350
rect 500878 388294 500934 388350
rect 501002 388294 501058 388350
rect 501126 388294 501182 388350
rect 500754 388170 500810 388226
rect 500878 388170 500934 388226
rect 501002 388170 501058 388226
rect 501126 388170 501182 388226
rect 500754 388046 500810 388102
rect 500878 388046 500934 388102
rect 501002 388046 501058 388102
rect 501126 388046 501182 388102
rect 500754 387922 500810 387978
rect 500878 387922 500934 387978
rect 501002 387922 501058 387978
rect 501126 387922 501182 387978
rect 523292 403082 523348 403138
rect 531474 598116 531530 598172
rect 531598 598116 531654 598172
rect 531722 598116 531778 598172
rect 531846 598116 531902 598172
rect 531474 597992 531530 598048
rect 531598 597992 531654 598048
rect 531722 597992 531778 598048
rect 531846 597992 531902 598048
rect 531474 597868 531530 597924
rect 531598 597868 531654 597924
rect 531722 597868 531778 597924
rect 531846 597868 531902 597924
rect 531474 597744 531530 597800
rect 531598 597744 531654 597800
rect 531722 597744 531778 597800
rect 531846 597744 531902 597800
rect 531474 586294 531530 586350
rect 531598 586294 531654 586350
rect 531722 586294 531778 586350
rect 531846 586294 531902 586350
rect 531474 586170 531530 586226
rect 531598 586170 531654 586226
rect 531722 586170 531778 586226
rect 531846 586170 531902 586226
rect 531474 586046 531530 586102
rect 531598 586046 531654 586102
rect 531722 586046 531778 586102
rect 531846 586046 531902 586102
rect 531474 585922 531530 585978
rect 531598 585922 531654 585978
rect 531722 585922 531778 585978
rect 531846 585922 531902 585978
rect 531474 568294 531530 568350
rect 531598 568294 531654 568350
rect 531722 568294 531778 568350
rect 531846 568294 531902 568350
rect 531474 568170 531530 568226
rect 531598 568170 531654 568226
rect 531722 568170 531778 568226
rect 531846 568170 531902 568226
rect 531474 568046 531530 568102
rect 531598 568046 531654 568102
rect 531722 568046 531778 568102
rect 531846 568046 531902 568102
rect 531474 567922 531530 567978
rect 531598 567922 531654 567978
rect 531722 567922 531778 567978
rect 531846 567922 531902 567978
rect 558474 597156 558530 597212
rect 558598 597156 558654 597212
rect 558722 597156 558778 597212
rect 558846 597156 558902 597212
rect 558474 597032 558530 597088
rect 558598 597032 558654 597088
rect 558722 597032 558778 597088
rect 558846 597032 558902 597088
rect 558474 596908 558530 596964
rect 558598 596908 558654 596964
rect 558722 596908 558778 596964
rect 558846 596908 558902 596964
rect 558474 596784 558530 596840
rect 558598 596784 558654 596840
rect 558722 596784 558778 596840
rect 558846 596784 558902 596840
rect 558474 580294 558530 580350
rect 558598 580294 558654 580350
rect 558722 580294 558778 580350
rect 558846 580294 558902 580350
rect 558474 580170 558530 580226
rect 558598 580170 558654 580226
rect 558722 580170 558778 580226
rect 558846 580170 558902 580226
rect 558474 580046 558530 580102
rect 558598 580046 558654 580102
rect 558722 580046 558778 580102
rect 558846 580046 558902 580102
rect 558474 579922 558530 579978
rect 558598 579922 558654 579978
rect 558722 579922 558778 579978
rect 558846 579922 558902 579978
rect 542518 562294 542574 562350
rect 542642 562294 542698 562350
rect 542518 562170 542574 562226
rect 542642 562170 542698 562226
rect 542518 562046 542574 562102
rect 542642 562046 542698 562102
rect 542518 561922 542574 561978
rect 542642 561922 542698 561978
rect 558474 562294 558530 562350
rect 558598 562294 558654 562350
rect 558722 562294 558778 562350
rect 558846 562294 558902 562350
rect 558474 562170 558530 562226
rect 558598 562170 558654 562226
rect 558722 562170 558778 562226
rect 558846 562170 558902 562226
rect 558474 562046 558530 562102
rect 558598 562046 558654 562102
rect 558722 562046 558778 562102
rect 558846 562046 558902 562102
rect 558474 561922 558530 561978
rect 558598 561922 558654 561978
rect 558722 561922 558778 561978
rect 558846 561922 558902 561978
rect 531474 550294 531530 550350
rect 531598 550294 531654 550350
rect 531722 550294 531778 550350
rect 531846 550294 531902 550350
rect 531474 550170 531530 550226
rect 531598 550170 531654 550226
rect 531722 550170 531778 550226
rect 531846 550170 531902 550226
rect 531474 550046 531530 550102
rect 531598 550046 531654 550102
rect 531722 550046 531778 550102
rect 531846 550046 531902 550102
rect 531474 549922 531530 549978
rect 531598 549922 531654 549978
rect 531722 549922 531778 549978
rect 531846 549922 531902 549978
rect 531474 532294 531530 532350
rect 531598 532294 531654 532350
rect 531722 532294 531778 532350
rect 531846 532294 531902 532350
rect 531474 532170 531530 532226
rect 531598 532170 531654 532226
rect 531722 532170 531778 532226
rect 531846 532170 531902 532226
rect 531474 532046 531530 532102
rect 531598 532046 531654 532102
rect 531722 532046 531778 532102
rect 531846 532046 531902 532102
rect 531474 531922 531530 531978
rect 531598 531922 531654 531978
rect 531722 531922 531778 531978
rect 531846 531922 531902 531978
rect 531474 514294 531530 514350
rect 531598 514294 531654 514350
rect 531722 514294 531778 514350
rect 531846 514294 531902 514350
rect 531474 514170 531530 514226
rect 531598 514170 531654 514226
rect 531722 514170 531778 514226
rect 531846 514170 531902 514226
rect 531474 514046 531530 514102
rect 531598 514046 531654 514102
rect 531722 514046 531778 514102
rect 531846 514046 531902 514102
rect 531474 513922 531530 513978
rect 531598 513922 531654 513978
rect 531722 513922 531778 513978
rect 531846 513922 531902 513978
rect 562194 598116 562250 598172
rect 562318 598116 562374 598172
rect 562442 598116 562498 598172
rect 562566 598116 562622 598172
rect 562194 597992 562250 598048
rect 562318 597992 562374 598048
rect 562442 597992 562498 598048
rect 562566 597992 562622 598048
rect 562194 597868 562250 597924
rect 562318 597868 562374 597924
rect 562442 597868 562498 597924
rect 562566 597868 562622 597924
rect 562194 597744 562250 597800
rect 562318 597744 562374 597800
rect 562442 597744 562498 597800
rect 562566 597744 562622 597800
rect 562194 586294 562250 586350
rect 562318 586294 562374 586350
rect 562442 586294 562498 586350
rect 562566 586294 562622 586350
rect 562194 586170 562250 586226
rect 562318 586170 562374 586226
rect 562442 586170 562498 586226
rect 562566 586170 562622 586226
rect 562194 586046 562250 586102
rect 562318 586046 562374 586102
rect 562442 586046 562498 586102
rect 562566 586046 562622 586102
rect 562194 585922 562250 585978
rect 562318 585922 562374 585978
rect 562442 585922 562498 585978
rect 562566 585922 562622 585978
rect 562194 568294 562250 568350
rect 562318 568294 562374 568350
rect 562442 568294 562498 568350
rect 562566 568294 562622 568350
rect 562194 568170 562250 568226
rect 562318 568170 562374 568226
rect 562442 568170 562498 568226
rect 562566 568170 562622 568226
rect 562194 568046 562250 568102
rect 562318 568046 562374 568102
rect 562442 568046 562498 568102
rect 562566 568046 562622 568102
rect 562194 567922 562250 567978
rect 562318 567922 562374 567978
rect 562442 567922 562498 567978
rect 562566 567922 562622 567978
rect 557878 550294 557934 550350
rect 558002 550294 558058 550350
rect 557878 550170 557934 550226
rect 558002 550170 558058 550226
rect 557878 550046 557934 550102
rect 558002 550046 558058 550102
rect 557878 549922 557934 549978
rect 558002 549922 558058 549978
rect 589194 597156 589250 597212
rect 589318 597156 589374 597212
rect 589442 597156 589498 597212
rect 589566 597156 589622 597212
rect 589194 597032 589250 597088
rect 589318 597032 589374 597088
rect 589442 597032 589498 597088
rect 589566 597032 589622 597088
rect 589194 596908 589250 596964
rect 589318 596908 589374 596964
rect 589442 596908 589498 596964
rect 589566 596908 589622 596964
rect 589194 596784 589250 596840
rect 589318 596784 589374 596840
rect 589442 596784 589498 596840
rect 589566 596784 589622 596840
rect 589194 580294 589250 580350
rect 589318 580294 589374 580350
rect 589442 580294 589498 580350
rect 589566 580294 589622 580350
rect 589194 580170 589250 580226
rect 589318 580170 589374 580226
rect 589442 580170 589498 580226
rect 589566 580170 589622 580226
rect 589194 580046 589250 580102
rect 589318 580046 589374 580102
rect 589442 580046 589498 580102
rect 589566 580046 589622 580102
rect 589194 579922 589250 579978
rect 589318 579922 589374 579978
rect 589442 579922 589498 579978
rect 589566 579922 589622 579978
rect 585452 566882 585508 566938
rect 573238 562294 573294 562350
rect 573362 562294 573418 562350
rect 573238 562170 573294 562226
rect 573362 562170 573418 562226
rect 573238 562046 573294 562102
rect 573362 562046 573418 562102
rect 573238 561922 573294 561978
rect 573362 561922 573418 561978
rect 562194 550294 562250 550350
rect 562318 550294 562374 550350
rect 562442 550294 562498 550350
rect 562566 550294 562622 550350
rect 562194 550170 562250 550226
rect 562318 550170 562374 550226
rect 562442 550170 562498 550226
rect 562566 550170 562622 550226
rect 562194 550046 562250 550102
rect 562318 550046 562374 550102
rect 562442 550046 562498 550102
rect 562566 550046 562622 550102
rect 562194 549922 562250 549978
rect 562318 549922 562374 549978
rect 562442 549922 562498 549978
rect 562566 549922 562622 549978
rect 542518 544294 542574 544350
rect 542642 544294 542698 544350
rect 542518 544170 542574 544226
rect 542642 544170 542698 544226
rect 542518 544046 542574 544102
rect 542642 544046 542698 544102
rect 542518 543922 542574 543978
rect 542642 543922 542698 543978
rect 558474 544294 558530 544350
rect 558598 544294 558654 544350
rect 558722 544294 558778 544350
rect 558846 544294 558902 544350
rect 558474 544170 558530 544226
rect 558598 544170 558654 544226
rect 558722 544170 558778 544226
rect 558846 544170 558902 544226
rect 558474 544046 558530 544102
rect 558598 544046 558654 544102
rect 558722 544046 558778 544102
rect 558846 544046 558902 544102
rect 558474 543922 558530 543978
rect 558598 543922 558654 543978
rect 558722 543922 558778 543978
rect 558846 543922 558902 543978
rect 557878 532294 557934 532350
rect 558002 532294 558058 532350
rect 557878 532170 557934 532226
rect 558002 532170 558058 532226
rect 557878 532046 557934 532102
rect 558002 532046 558058 532102
rect 557878 531922 557934 531978
rect 558002 531922 558058 531978
rect 558474 526294 558530 526350
rect 558598 526294 558654 526350
rect 558722 526294 558778 526350
rect 558846 526294 558902 526350
rect 558474 526170 558530 526226
rect 558598 526170 558654 526226
rect 558722 526170 558778 526226
rect 558846 526170 558902 526226
rect 558474 526046 558530 526102
rect 558598 526046 558654 526102
rect 558722 526046 558778 526102
rect 558846 526046 558902 526102
rect 558474 525922 558530 525978
rect 558598 525922 558654 525978
rect 558722 525922 558778 525978
rect 558846 525922 558902 525978
rect 558474 508294 558530 508350
rect 558598 508294 558654 508350
rect 558722 508294 558778 508350
rect 558846 508294 558902 508350
rect 558474 508170 558530 508226
rect 558598 508170 558654 508226
rect 558722 508170 558778 508226
rect 558846 508170 558902 508226
rect 558474 508046 558530 508102
rect 558598 508046 558654 508102
rect 558722 508046 558778 508102
rect 558846 508046 558902 508102
rect 558474 507922 558530 507978
rect 558598 507922 558654 507978
rect 558722 507922 558778 507978
rect 558846 507922 558902 507978
rect 531474 496294 531530 496350
rect 531598 496294 531654 496350
rect 531722 496294 531778 496350
rect 531846 496294 531902 496350
rect 531474 496170 531530 496226
rect 531598 496170 531654 496226
rect 531722 496170 531778 496226
rect 531846 496170 531902 496226
rect 531474 496046 531530 496102
rect 531598 496046 531654 496102
rect 531722 496046 531778 496102
rect 531846 496046 531902 496102
rect 531474 495922 531530 495978
rect 531598 495922 531654 495978
rect 531722 495922 531778 495978
rect 531846 495922 531902 495978
rect 542518 490294 542574 490350
rect 542642 490294 542698 490350
rect 542518 490170 542574 490226
rect 542642 490170 542698 490226
rect 542518 490046 542574 490102
rect 542642 490046 542698 490102
rect 542518 489922 542574 489978
rect 542642 489922 542698 489978
rect 558474 490294 558530 490350
rect 558598 490294 558654 490350
rect 558722 490294 558778 490350
rect 558846 490294 558902 490350
rect 558474 490170 558530 490226
rect 558598 490170 558654 490226
rect 558722 490170 558778 490226
rect 558846 490170 558902 490226
rect 558474 490046 558530 490102
rect 558598 490046 558654 490102
rect 558722 490046 558778 490102
rect 558846 490046 558902 490102
rect 558474 489922 558530 489978
rect 558598 489922 558654 489978
rect 558722 489922 558778 489978
rect 558846 489922 558902 489978
rect 534268 484652 534324 484678
rect 534268 484622 534324 484652
rect 573238 544294 573294 544350
rect 573362 544294 573418 544350
rect 573238 544170 573294 544226
rect 573362 544170 573418 544226
rect 573238 544046 573294 544102
rect 573362 544046 573418 544102
rect 573238 543922 573294 543978
rect 573362 543922 573418 543978
rect 562194 532294 562250 532350
rect 562318 532294 562374 532350
rect 562442 532294 562498 532350
rect 562566 532294 562622 532350
rect 562194 532170 562250 532226
rect 562318 532170 562374 532226
rect 562442 532170 562498 532226
rect 562566 532170 562622 532226
rect 562194 532046 562250 532102
rect 562318 532046 562374 532102
rect 562442 532046 562498 532102
rect 562566 532046 562622 532102
rect 562194 531922 562250 531978
rect 562318 531922 562374 531978
rect 562442 531922 562498 531978
rect 562566 531922 562622 531978
rect 562194 514294 562250 514350
rect 562318 514294 562374 514350
rect 562442 514294 562498 514350
rect 562566 514294 562622 514350
rect 562194 514170 562250 514226
rect 562318 514170 562374 514226
rect 562442 514170 562498 514226
rect 562566 514170 562622 514226
rect 562194 514046 562250 514102
rect 562318 514046 562374 514102
rect 562442 514046 562498 514102
rect 562566 514046 562622 514102
rect 562194 513922 562250 513978
rect 562318 513922 562374 513978
rect 562442 513922 562498 513978
rect 562566 513922 562622 513978
rect 562194 496294 562250 496350
rect 562318 496294 562374 496350
rect 562442 496294 562498 496350
rect 562566 496294 562622 496350
rect 562194 496170 562250 496226
rect 562318 496170 562374 496226
rect 562442 496170 562498 496226
rect 562566 496170 562622 496226
rect 562194 496046 562250 496102
rect 562318 496046 562374 496102
rect 562442 496046 562498 496102
rect 562566 496046 562622 496102
rect 562194 495922 562250 495978
rect 562318 495922 562374 495978
rect 562442 495922 562498 495978
rect 562566 495922 562622 495978
rect 531474 478294 531530 478350
rect 531598 478294 531654 478350
rect 531722 478294 531778 478350
rect 531846 478294 531902 478350
rect 531474 478170 531530 478226
rect 531598 478170 531654 478226
rect 531722 478170 531778 478226
rect 531846 478170 531902 478226
rect 531474 478046 531530 478102
rect 531598 478046 531654 478102
rect 531722 478046 531778 478102
rect 531846 478046 531902 478102
rect 531474 477922 531530 477978
rect 531598 477922 531654 477978
rect 531722 477922 531778 477978
rect 531846 477922 531902 477978
rect 531474 460294 531530 460350
rect 531598 460294 531654 460350
rect 531722 460294 531778 460350
rect 531846 460294 531902 460350
rect 531474 460170 531530 460226
rect 531598 460170 531654 460226
rect 531722 460170 531778 460226
rect 531846 460170 531902 460226
rect 531474 460046 531530 460102
rect 531598 460046 531654 460102
rect 531722 460046 531778 460102
rect 531846 460046 531902 460102
rect 531474 459922 531530 459978
rect 531598 459922 531654 459978
rect 531722 459922 531778 459978
rect 531846 459922 531902 459978
rect 554316 480482 554372 480538
rect 557878 478294 557934 478350
rect 558002 478294 558058 478350
rect 557878 478170 557934 478226
rect 558002 478170 558058 478226
rect 557878 478046 557934 478102
rect 558002 478046 558058 478102
rect 557878 477922 557934 477978
rect 558002 477922 558058 477978
rect 573238 490294 573294 490350
rect 573362 490294 573418 490350
rect 573238 490170 573294 490226
rect 573362 490170 573418 490226
rect 573238 490046 573294 490102
rect 573362 490046 573418 490102
rect 573238 489922 573294 489978
rect 573362 489922 573418 489978
rect 579628 480482 579684 480538
rect 562194 478294 562250 478350
rect 562318 478294 562374 478350
rect 562442 478294 562498 478350
rect 562566 478294 562622 478350
rect 562194 478170 562250 478226
rect 562318 478170 562374 478226
rect 562442 478170 562498 478226
rect 562566 478170 562622 478226
rect 562194 478046 562250 478102
rect 562318 478046 562374 478102
rect 562442 478046 562498 478102
rect 562566 478046 562622 478102
rect 562194 477922 562250 477978
rect 562318 477922 562374 477978
rect 562442 477922 562498 477978
rect 562566 477922 562622 477978
rect 554316 473642 554372 473698
rect 542518 472294 542574 472350
rect 542642 472294 542698 472350
rect 542518 472170 542574 472226
rect 542642 472170 542698 472226
rect 542518 472046 542574 472102
rect 542642 472046 542698 472102
rect 542518 471922 542574 471978
rect 542642 471922 542698 471978
rect 554092 470402 554148 470458
rect 554092 468422 554148 468478
rect 557878 460294 557934 460350
rect 558002 460294 558058 460350
rect 557878 460170 557934 460226
rect 558002 460170 558058 460226
rect 557878 460046 557934 460102
rect 558002 460046 558058 460102
rect 557878 459922 557934 459978
rect 558002 459922 558058 459978
rect 558474 454294 558530 454350
rect 558598 454294 558654 454350
rect 558722 454294 558778 454350
rect 558846 454294 558902 454350
rect 558474 454170 558530 454226
rect 558598 454170 558654 454226
rect 558722 454170 558778 454226
rect 558846 454170 558902 454226
rect 558474 454046 558530 454102
rect 558598 454046 558654 454102
rect 558722 454046 558778 454102
rect 558846 454046 558902 454102
rect 558474 453922 558530 453978
rect 558598 453922 558654 453978
rect 558722 453922 558778 453978
rect 558846 453922 558902 453978
rect 531474 442294 531530 442350
rect 531598 442294 531654 442350
rect 531722 442294 531778 442350
rect 531846 442294 531902 442350
rect 531474 442170 531530 442226
rect 531598 442170 531654 442226
rect 531722 442170 531778 442226
rect 531846 442170 531902 442226
rect 531474 442046 531530 442102
rect 531598 442046 531654 442102
rect 531722 442046 531778 442102
rect 531846 442046 531902 442102
rect 531474 441922 531530 441978
rect 531598 441922 531654 441978
rect 531722 441922 531778 441978
rect 531846 441922 531902 441978
rect 531474 424294 531530 424350
rect 531598 424294 531654 424350
rect 531722 424294 531778 424350
rect 531846 424294 531902 424350
rect 531474 424170 531530 424226
rect 531598 424170 531654 424226
rect 531722 424170 531778 424226
rect 531846 424170 531902 424226
rect 531474 424046 531530 424102
rect 531598 424046 531654 424102
rect 531722 424046 531778 424102
rect 531846 424046 531902 424102
rect 531474 423922 531530 423978
rect 531598 423922 531654 423978
rect 531722 423922 531778 423978
rect 531846 423922 531902 423978
rect 527754 400294 527810 400350
rect 527878 400294 527934 400350
rect 528002 400294 528058 400350
rect 528126 400294 528182 400350
rect 527754 400170 527810 400226
rect 527878 400170 527934 400226
rect 528002 400170 528058 400226
rect 528126 400170 528182 400226
rect 527754 400046 527810 400102
rect 527878 400046 527934 400102
rect 528002 400046 528058 400102
rect 528126 400046 528182 400102
rect 527754 399922 527810 399978
rect 527878 399922 527934 399978
rect 528002 399922 528058 399978
rect 528126 399922 528182 399978
rect 527754 382294 527810 382350
rect 527878 382294 527934 382350
rect 528002 382294 528058 382350
rect 528126 382294 528182 382350
rect 527754 382170 527810 382226
rect 527878 382170 527934 382226
rect 528002 382170 528058 382226
rect 528126 382170 528182 382226
rect 527754 382046 527810 382102
rect 527878 382046 527934 382102
rect 528002 382046 528058 382102
rect 528126 382046 528182 382102
rect 527754 381922 527810 381978
rect 527878 381922 527934 381978
rect 528002 381922 528058 381978
rect 528126 381922 528182 381978
rect 500754 370294 500810 370350
rect 500878 370294 500934 370350
rect 501002 370294 501058 370350
rect 501126 370294 501182 370350
rect 500754 370170 500810 370226
rect 500878 370170 500934 370226
rect 501002 370170 501058 370226
rect 501126 370170 501182 370226
rect 500754 370046 500810 370102
rect 500878 370046 500934 370102
rect 501002 370046 501058 370102
rect 501126 370046 501182 370102
rect 500754 369922 500810 369978
rect 500878 369922 500934 369978
rect 501002 369922 501058 369978
rect 501126 369922 501182 369978
rect 558474 436294 558530 436350
rect 558598 436294 558654 436350
rect 558722 436294 558778 436350
rect 558846 436294 558902 436350
rect 558474 436170 558530 436226
rect 558598 436170 558654 436226
rect 558722 436170 558778 436226
rect 558846 436170 558902 436226
rect 558474 436046 558530 436102
rect 558598 436046 558654 436102
rect 558722 436046 558778 436102
rect 558846 436046 558902 436102
rect 558474 435922 558530 435978
rect 558598 435922 558654 435978
rect 558722 435922 558778 435978
rect 558846 435922 558902 435978
rect 542518 418294 542574 418350
rect 542642 418294 542698 418350
rect 542518 418170 542574 418226
rect 542642 418170 542698 418226
rect 542518 418046 542574 418102
rect 542642 418046 542698 418102
rect 542518 417922 542574 417978
rect 542642 417922 542698 417978
rect 558474 418294 558530 418350
rect 558598 418294 558654 418350
rect 558722 418294 558778 418350
rect 558846 418294 558902 418350
rect 558474 418170 558530 418226
rect 558598 418170 558654 418226
rect 558722 418170 558778 418226
rect 558846 418170 558902 418226
rect 558474 418046 558530 418102
rect 558598 418046 558654 418102
rect 558722 418046 558778 418102
rect 558846 418046 558902 418102
rect 558474 417922 558530 417978
rect 558598 417922 558654 417978
rect 558722 417922 558778 417978
rect 558846 417922 558902 417978
rect 534380 409922 534436 409978
rect 534268 409562 534324 409618
rect 531474 406294 531530 406350
rect 531598 406294 531654 406350
rect 531722 406294 531778 406350
rect 531846 406294 531902 406350
rect 531474 406170 531530 406226
rect 531598 406170 531654 406226
rect 531722 406170 531778 406226
rect 531846 406170 531902 406226
rect 531474 406046 531530 406102
rect 531598 406046 531654 406102
rect 531722 406046 531778 406102
rect 531846 406046 531902 406102
rect 531474 405922 531530 405978
rect 531598 405922 531654 405978
rect 531722 405922 531778 405978
rect 531846 405922 531902 405978
rect 531474 388294 531530 388350
rect 531598 388294 531654 388350
rect 531722 388294 531778 388350
rect 531846 388294 531902 388350
rect 531474 388170 531530 388226
rect 531598 388170 531654 388226
rect 531722 388170 531778 388226
rect 531846 388170 531902 388226
rect 531474 388046 531530 388102
rect 531598 388046 531654 388102
rect 531722 388046 531778 388102
rect 531846 388046 531902 388102
rect 531474 387922 531530 387978
rect 531598 387922 531654 387978
rect 531722 387922 531778 387978
rect 531846 387922 531902 387978
rect 527754 364294 527810 364350
rect 527878 364294 527934 364350
rect 528002 364294 528058 364350
rect 528126 364294 528182 364350
rect 527754 364170 527810 364226
rect 527878 364170 527934 364226
rect 528002 364170 528058 364226
rect 528126 364170 528182 364226
rect 527754 364046 527810 364102
rect 527878 364046 527934 364102
rect 528002 364046 528058 364102
rect 528126 364046 528182 364102
rect 527754 363922 527810 363978
rect 527878 363922 527934 363978
rect 528002 363922 528058 363978
rect 528126 363922 528182 363978
rect 500754 352294 500810 352350
rect 500878 352294 500934 352350
rect 501002 352294 501058 352350
rect 501126 352294 501182 352350
rect 500754 352170 500810 352226
rect 500878 352170 500934 352226
rect 501002 352170 501058 352226
rect 501126 352170 501182 352226
rect 500754 352046 500810 352102
rect 500878 352046 500934 352102
rect 501002 352046 501058 352102
rect 501126 352046 501182 352102
rect 500754 351922 500810 351978
rect 500878 351922 500934 351978
rect 501002 351922 501058 351978
rect 501126 351922 501182 351978
rect 495878 334294 495934 334350
rect 496002 334294 496058 334350
rect 495878 334170 495934 334226
rect 496002 334170 496058 334226
rect 495878 334046 495934 334102
rect 496002 334046 496058 334102
rect 495878 333922 495934 333978
rect 496002 333922 496058 333978
rect 511238 346294 511294 346350
rect 511362 346294 511418 346350
rect 511238 346170 511294 346226
rect 511362 346170 511418 346226
rect 511238 346046 511294 346102
rect 511362 346046 511418 346102
rect 511238 345922 511294 345978
rect 511362 345922 511418 345978
rect 523292 349442 523348 349498
rect 521052 343502 521108 343558
rect 520940 340082 520996 340138
rect 517468 338822 517524 338878
rect 500754 334294 500810 334350
rect 500878 334294 500934 334350
rect 501002 334294 501058 334350
rect 501126 334294 501182 334350
rect 500754 334170 500810 334226
rect 500878 334170 500934 334226
rect 501002 334170 501058 334226
rect 501126 334170 501182 334226
rect 500754 334046 500810 334102
rect 500878 334046 500934 334102
rect 501002 334046 501058 334102
rect 501126 334046 501182 334102
rect 500754 333922 500810 333978
rect 500878 333922 500934 333978
rect 501002 333922 501058 333978
rect 501126 333922 501182 333978
rect 480518 328294 480574 328350
rect 480642 328294 480698 328350
rect 480518 328170 480574 328226
rect 480642 328170 480698 328226
rect 480518 328046 480574 328102
rect 480642 328046 480698 328102
rect 480518 327922 480574 327978
rect 480642 327922 480698 327978
rect 497034 328294 497090 328350
rect 497158 328294 497214 328350
rect 497282 328294 497338 328350
rect 497406 328294 497462 328350
rect 497034 328170 497090 328226
rect 497158 328170 497214 328226
rect 497282 328170 497338 328226
rect 497406 328170 497462 328226
rect 497034 328046 497090 328102
rect 497158 328046 497214 328102
rect 497282 328046 497338 328102
rect 497406 328046 497462 328102
rect 497034 327922 497090 327978
rect 497158 327922 497214 327978
rect 497282 327922 497338 327978
rect 497406 327922 497462 327978
rect 470034 316294 470090 316350
rect 470158 316294 470214 316350
rect 470282 316294 470338 316350
rect 470406 316294 470462 316350
rect 470034 316170 470090 316226
rect 470158 316170 470214 316226
rect 470282 316170 470338 316226
rect 470406 316170 470462 316226
rect 470034 316046 470090 316102
rect 470158 316046 470214 316102
rect 470282 316046 470338 316102
rect 470406 316046 470462 316102
rect 470034 315922 470090 315978
rect 470158 315922 470214 315978
rect 470282 315922 470338 315978
rect 470406 315922 470462 315978
rect 470034 298294 470090 298350
rect 470158 298294 470214 298350
rect 470282 298294 470338 298350
rect 470406 298294 470462 298350
rect 470034 298170 470090 298226
rect 470158 298170 470214 298226
rect 470282 298170 470338 298226
rect 470406 298170 470462 298226
rect 470034 298046 470090 298102
rect 470158 298046 470214 298102
rect 470282 298046 470338 298102
rect 470406 298046 470462 298102
rect 470034 297922 470090 297978
rect 470158 297922 470214 297978
rect 470282 297922 470338 297978
rect 470406 297922 470462 297978
rect 497034 310294 497090 310350
rect 497158 310294 497214 310350
rect 497282 310294 497338 310350
rect 497406 310294 497462 310350
rect 497034 310170 497090 310226
rect 497158 310170 497214 310226
rect 497282 310170 497338 310226
rect 497406 310170 497462 310226
rect 497034 310046 497090 310102
rect 497158 310046 497214 310102
rect 497282 310046 497338 310102
rect 497406 310046 497462 310102
rect 497034 309922 497090 309978
rect 497158 309922 497214 309978
rect 497282 309922 497338 309978
rect 497406 309922 497462 309978
rect 497034 292294 497090 292350
rect 497158 292294 497214 292350
rect 497282 292294 497338 292350
rect 497406 292294 497462 292350
rect 497034 292170 497090 292226
rect 497158 292170 497214 292226
rect 497282 292170 497338 292226
rect 497406 292170 497462 292226
rect 497034 292046 497090 292102
rect 497158 292046 497214 292102
rect 497282 292046 497338 292102
rect 497406 292046 497462 292102
rect 497034 291922 497090 291978
rect 497158 291922 497214 291978
rect 497282 291922 497338 291978
rect 497406 291922 497462 291978
rect 470034 280294 470090 280350
rect 470158 280294 470214 280350
rect 470282 280294 470338 280350
rect 470406 280294 470462 280350
rect 470034 280170 470090 280226
rect 470158 280170 470214 280226
rect 470282 280170 470338 280226
rect 470406 280170 470462 280226
rect 470034 280046 470090 280102
rect 470158 280046 470214 280102
rect 470282 280046 470338 280102
rect 470406 280046 470462 280102
rect 470034 279922 470090 279978
rect 470158 279922 470214 279978
rect 470282 279922 470338 279978
rect 470406 279922 470462 279978
rect 472108 268982 472164 269038
rect 472108 267362 472164 267418
rect 495878 280294 495934 280350
rect 496002 280294 496058 280350
rect 495878 280170 495934 280226
rect 496002 280170 496058 280226
rect 495878 280046 495934 280102
rect 496002 280046 496058 280102
rect 495878 279922 495934 279978
rect 496002 279922 496058 279978
rect 480518 274294 480574 274350
rect 480642 274294 480698 274350
rect 480518 274170 480574 274226
rect 480642 274170 480698 274226
rect 480518 274046 480574 274102
rect 480642 274046 480698 274102
rect 480518 273922 480574 273978
rect 480642 273922 480698 273978
rect 497034 274294 497090 274350
rect 497158 274294 497214 274350
rect 497282 274294 497338 274350
rect 497406 274294 497462 274350
rect 497034 274170 497090 274226
rect 497158 274170 497214 274226
rect 497282 274170 497338 274226
rect 497406 274170 497462 274226
rect 497034 274046 497090 274102
rect 497158 274046 497214 274102
rect 497282 274046 497338 274102
rect 497406 274046 497462 274102
rect 497034 273922 497090 273978
rect 497158 273922 497214 273978
rect 497282 273922 497338 273978
rect 497406 273922 497462 273978
rect 473676 269522 473732 269578
rect 511238 328294 511294 328350
rect 511362 328294 511418 328350
rect 511238 328170 511294 328226
rect 511362 328170 511418 328226
rect 511238 328046 511294 328102
rect 511362 328046 511418 328102
rect 511238 327922 511294 327978
rect 511362 327922 511418 327978
rect 500754 316294 500810 316350
rect 500878 316294 500934 316350
rect 501002 316294 501058 316350
rect 501126 316294 501182 316350
rect 500754 316170 500810 316226
rect 500878 316170 500934 316226
rect 501002 316170 501058 316226
rect 501126 316170 501182 316226
rect 500754 316046 500810 316102
rect 500878 316046 500934 316102
rect 501002 316046 501058 316102
rect 501126 316046 501182 316102
rect 500754 315922 500810 315978
rect 500878 315922 500934 315978
rect 501002 315922 501058 315978
rect 501126 315922 501182 315978
rect 527754 346294 527810 346350
rect 527878 346294 527934 346350
rect 528002 346294 528058 346350
rect 528126 346294 528182 346350
rect 527754 346170 527810 346226
rect 527878 346170 527934 346226
rect 528002 346170 528058 346226
rect 528126 346170 528182 346226
rect 527754 346046 527810 346102
rect 527878 346046 527934 346102
rect 528002 346046 528058 346102
rect 528126 346046 528182 346102
rect 527754 345922 527810 345978
rect 527878 345922 527934 345978
rect 528002 345922 528058 345978
rect 528126 345922 528182 345978
rect 523292 324062 523348 324118
rect 527754 328294 527810 328350
rect 527878 328294 527934 328350
rect 528002 328294 528058 328350
rect 528126 328294 528182 328350
rect 527754 328170 527810 328226
rect 527878 328170 527934 328226
rect 528002 328170 528058 328226
rect 528126 328170 528182 328226
rect 527754 328046 527810 328102
rect 527878 328046 527934 328102
rect 528002 328046 528058 328102
rect 528126 328046 528182 328102
rect 527754 327922 527810 327978
rect 527878 327922 527934 327978
rect 528002 327922 528058 327978
rect 528126 327922 528182 327978
rect 500754 298294 500810 298350
rect 500878 298294 500934 298350
rect 501002 298294 501058 298350
rect 501126 298294 501182 298350
rect 500754 298170 500810 298226
rect 500878 298170 500934 298226
rect 501002 298170 501058 298226
rect 501126 298170 501182 298226
rect 500754 298046 500810 298102
rect 500878 298046 500934 298102
rect 501002 298046 501058 298102
rect 501126 298046 501182 298102
rect 500754 297922 500810 297978
rect 500878 297922 500934 297978
rect 501002 297922 501058 297978
rect 501126 297922 501182 297978
rect 527754 310294 527810 310350
rect 527878 310294 527934 310350
rect 528002 310294 528058 310350
rect 528126 310294 528182 310350
rect 527754 310170 527810 310226
rect 527878 310170 527934 310226
rect 528002 310170 528058 310226
rect 528126 310170 528182 310226
rect 527754 310046 527810 310102
rect 527878 310046 527934 310102
rect 528002 310046 528058 310102
rect 528126 310046 528182 310102
rect 527754 309922 527810 309978
rect 527878 309922 527934 309978
rect 528002 309922 528058 309978
rect 528126 309922 528182 309978
rect 500754 280294 500810 280350
rect 500878 280294 500934 280350
rect 501002 280294 501058 280350
rect 501126 280294 501182 280350
rect 500754 280170 500810 280226
rect 500878 280170 500934 280226
rect 501002 280170 501058 280226
rect 501126 280170 501182 280226
rect 500754 280046 500810 280102
rect 500878 280046 500934 280102
rect 501002 280046 501058 280102
rect 501126 280046 501182 280102
rect 500754 279922 500810 279978
rect 500878 279922 500934 279978
rect 501002 279922 501058 279978
rect 501126 279922 501182 279978
rect 511238 274294 511294 274350
rect 511362 274294 511418 274350
rect 511238 274170 511294 274226
rect 511362 274170 511418 274226
rect 511238 274046 511294 274102
rect 511362 274046 511418 274102
rect 511238 273922 511294 273978
rect 511362 273922 511418 273978
rect 517468 267182 517524 267238
rect 470034 262294 470090 262350
rect 470158 262294 470214 262350
rect 470282 262294 470338 262350
rect 470406 262294 470462 262350
rect 470034 262170 470090 262226
rect 470158 262170 470214 262226
rect 470282 262170 470338 262226
rect 470406 262170 470462 262226
rect 468636 258542 468692 258598
rect 470034 262046 470090 262102
rect 470158 262046 470214 262102
rect 470282 262046 470338 262102
rect 470406 262046 470462 262102
rect 470034 261922 470090 261978
rect 470158 261922 470214 261978
rect 470282 261922 470338 261978
rect 470406 261922 470462 261978
rect 466314 256294 466370 256350
rect 466438 256294 466494 256350
rect 466562 256294 466618 256350
rect 466686 256294 466742 256350
rect 466314 256170 466370 256226
rect 466438 256170 466494 256226
rect 466562 256170 466618 256226
rect 466686 256170 466742 256226
rect 466314 256046 466370 256102
rect 466438 256046 466494 256102
rect 466562 256046 466618 256102
rect 466686 256046 466742 256102
rect 466314 255922 466370 255978
rect 466438 255922 466494 255978
rect 466562 255922 466618 255978
rect 466686 255922 466742 255978
rect 461132 255122 461188 255178
rect 458892 250262 458948 250318
rect 439314 244294 439370 244350
rect 439438 244294 439494 244350
rect 439562 244294 439618 244350
rect 439686 244294 439742 244350
rect 439314 244170 439370 244226
rect 439438 244170 439494 244226
rect 439562 244170 439618 244226
rect 439686 244170 439742 244226
rect 439314 244046 439370 244102
rect 439438 244046 439494 244102
rect 439562 244046 439618 244102
rect 439686 244046 439742 244102
rect 439314 243922 439370 243978
rect 439438 243922 439494 243978
rect 439562 243922 439618 243978
rect 439686 243922 439742 243978
rect 466314 238294 466370 238350
rect 466438 238294 466494 238350
rect 466562 238294 466618 238350
rect 466686 238294 466742 238350
rect 466314 238170 466370 238226
rect 466438 238170 466494 238226
rect 466562 238170 466618 238226
rect 466686 238170 466742 238226
rect 466314 238046 466370 238102
rect 466438 238046 466494 238102
rect 466562 238046 466618 238102
rect 466686 238046 466742 238102
rect 466314 237922 466370 237978
rect 466438 237922 466494 237978
rect 466562 237922 466618 237978
rect 466686 237922 466742 237978
rect 439314 226294 439370 226350
rect 439438 226294 439494 226350
rect 439562 226294 439618 226350
rect 439686 226294 439742 226350
rect 439314 226170 439370 226226
rect 439438 226170 439494 226226
rect 439562 226170 439618 226226
rect 439686 226170 439742 226226
rect 439314 226046 439370 226102
rect 439438 226046 439494 226102
rect 439562 226046 439618 226102
rect 439686 226046 439742 226102
rect 439314 225922 439370 225978
rect 439438 225922 439494 225978
rect 439562 225922 439618 225978
rect 439686 225922 439742 225978
rect 439314 208294 439370 208350
rect 439438 208294 439494 208350
rect 439562 208294 439618 208350
rect 439686 208294 439742 208350
rect 439314 208170 439370 208226
rect 439438 208170 439494 208226
rect 439562 208170 439618 208226
rect 439686 208170 439742 208226
rect 439314 208046 439370 208102
rect 439438 208046 439494 208102
rect 439562 208046 439618 208102
rect 439686 208046 439742 208102
rect 439314 207922 439370 207978
rect 439438 207922 439494 207978
rect 439562 207922 439618 207978
rect 439686 207922 439742 207978
rect 449238 202294 449294 202350
rect 449362 202294 449418 202350
rect 449238 202170 449294 202226
rect 449362 202170 449418 202226
rect 449238 202046 449294 202102
rect 449362 202046 449418 202102
rect 449238 201922 449294 201978
rect 449362 201922 449418 201978
rect 455308 198422 455364 198478
rect 456092 196802 456148 196858
rect 455308 193922 455364 193978
rect 439314 190294 439370 190350
rect 439438 190294 439494 190350
rect 439562 190294 439618 190350
rect 439686 190294 439742 190350
rect 439314 190170 439370 190226
rect 439438 190170 439494 190226
rect 439562 190170 439618 190226
rect 439686 190170 439742 190226
rect 439314 190046 439370 190102
rect 439438 190046 439494 190102
rect 439562 190046 439618 190102
rect 439686 190046 439742 190102
rect 439314 189922 439370 189978
rect 439438 189922 439494 189978
rect 439562 189922 439618 189978
rect 439686 189922 439742 189978
rect 455420 192122 455476 192178
rect 455308 186396 455364 186418
rect 455308 186362 455364 186396
rect 466314 220294 466370 220350
rect 466438 220294 466494 220350
rect 466562 220294 466618 220350
rect 466686 220294 466742 220350
rect 466314 220170 466370 220226
rect 466438 220170 466494 220226
rect 466562 220170 466618 220226
rect 466686 220170 466742 220226
rect 466314 220046 466370 220102
rect 466438 220046 466494 220102
rect 466562 220046 466618 220102
rect 466686 220046 466742 220102
rect 466314 219922 466370 219978
rect 466438 219922 466494 219978
rect 466562 219922 466618 219978
rect 466686 219922 466742 219978
rect 466314 202294 466370 202350
rect 466438 202294 466494 202350
rect 466562 202294 466618 202350
rect 466686 202294 466742 202350
rect 466314 202170 466370 202226
rect 466438 202170 466494 202226
rect 466562 202170 466618 202226
rect 466686 202170 466742 202226
rect 466314 202046 466370 202102
rect 466438 202046 466494 202102
rect 466562 202046 466618 202102
rect 466686 202046 466742 202102
rect 466314 201922 466370 201978
rect 466438 201922 466494 201978
rect 466562 201922 466618 201978
rect 466686 201922 466742 201978
rect 463596 196622 463652 196678
rect 449238 184294 449294 184350
rect 449362 184294 449418 184350
rect 449238 184170 449294 184226
rect 449362 184170 449418 184226
rect 449238 184046 449294 184102
rect 449362 184046 449418 184102
rect 449238 183922 449294 183978
rect 449362 183922 449418 183978
rect 495878 262294 495934 262350
rect 496002 262294 496058 262350
rect 495878 262170 495934 262226
rect 496002 262170 496058 262226
rect 495878 262046 495934 262102
rect 496002 262046 496058 262102
rect 495878 261922 495934 261978
rect 496002 261922 496058 261978
rect 472108 258722 472164 258778
rect 480518 256294 480574 256350
rect 480642 256294 480698 256350
rect 480518 256170 480574 256226
rect 480642 256170 480698 256226
rect 480518 256046 480574 256102
rect 480642 256046 480698 256102
rect 480518 255922 480574 255978
rect 480642 255922 480698 255978
rect 497034 256294 497090 256350
rect 497158 256294 497214 256350
rect 497282 256294 497338 256350
rect 497406 256294 497462 256350
rect 497034 256170 497090 256226
rect 497158 256170 497214 256226
rect 497282 256170 497338 256226
rect 497406 256170 497462 256226
rect 497034 256046 497090 256102
rect 497158 256046 497214 256102
rect 497282 256046 497338 256102
rect 497406 256046 497462 256102
rect 497034 255922 497090 255978
rect 497158 255922 497214 255978
rect 497282 255922 497338 255978
rect 497406 255922 497462 255978
rect 470034 244294 470090 244350
rect 470158 244294 470214 244350
rect 470282 244294 470338 244350
rect 470406 244294 470462 244350
rect 470034 244170 470090 244226
rect 470158 244170 470214 244226
rect 470282 244170 470338 244226
rect 470406 244170 470462 244226
rect 470034 244046 470090 244102
rect 470158 244046 470214 244102
rect 470282 244046 470338 244102
rect 470406 244046 470462 244102
rect 470034 243922 470090 243978
rect 470158 243922 470214 243978
rect 470282 243922 470338 243978
rect 470406 243922 470462 243978
rect 470034 226294 470090 226350
rect 470158 226294 470214 226350
rect 470282 226294 470338 226350
rect 470406 226294 470462 226350
rect 470034 226170 470090 226226
rect 470158 226170 470214 226226
rect 470282 226170 470338 226226
rect 470406 226170 470462 226226
rect 470034 226046 470090 226102
rect 470158 226046 470214 226102
rect 470282 226046 470338 226102
rect 470406 226046 470462 226102
rect 470034 225922 470090 225978
rect 470158 225922 470214 225978
rect 470282 225922 470338 225978
rect 470406 225922 470462 225978
rect 497034 238294 497090 238350
rect 497158 238294 497214 238350
rect 497282 238294 497338 238350
rect 497406 238294 497462 238350
rect 497034 238170 497090 238226
rect 497158 238170 497214 238226
rect 497282 238170 497338 238226
rect 497406 238170 497462 238226
rect 497034 238046 497090 238102
rect 497158 238046 497214 238102
rect 497282 238046 497338 238102
rect 497406 238046 497462 238102
rect 497034 237922 497090 237978
rect 497158 237922 497214 237978
rect 497282 237922 497338 237978
rect 497406 237922 497462 237978
rect 497034 220294 497090 220350
rect 497158 220294 497214 220350
rect 497282 220294 497338 220350
rect 497406 220294 497462 220350
rect 497034 220170 497090 220226
rect 497158 220170 497214 220226
rect 497282 220170 497338 220226
rect 497406 220170 497462 220226
rect 497034 220046 497090 220102
rect 497158 220046 497214 220102
rect 497282 220046 497338 220102
rect 497406 220046 497462 220102
rect 497034 219922 497090 219978
rect 497158 219922 497214 219978
rect 497282 219922 497338 219978
rect 497406 219922 497462 219978
rect 470034 208294 470090 208350
rect 470158 208294 470214 208350
rect 470282 208294 470338 208350
rect 470406 208294 470462 208350
rect 470034 208170 470090 208226
rect 470158 208170 470214 208226
rect 470282 208170 470338 208226
rect 470406 208170 470462 208226
rect 470034 208046 470090 208102
rect 470158 208046 470214 208102
rect 470282 208046 470338 208102
rect 470406 208046 470462 208102
rect 470034 207922 470090 207978
rect 470158 207922 470214 207978
rect 470282 207922 470338 207978
rect 470406 207922 470462 207978
rect 467852 200042 467908 200098
rect 466314 184294 466370 184350
rect 466438 184294 466494 184350
rect 466562 184294 466618 184350
rect 466686 184294 466742 184350
rect 466314 184170 466370 184226
rect 466438 184170 466494 184226
rect 466562 184170 466618 184226
rect 466686 184170 466742 184226
rect 466314 184046 466370 184102
rect 466438 184046 466494 184102
rect 466562 184046 466618 184102
rect 466686 184046 466742 184102
rect 466314 183922 466370 183978
rect 466438 183922 466494 183978
rect 466562 183922 466618 183978
rect 466686 183922 466742 183978
rect 439314 172294 439370 172350
rect 439438 172294 439494 172350
rect 439562 172294 439618 172350
rect 439686 172294 439742 172350
rect 439314 172170 439370 172226
rect 439438 172170 439494 172226
rect 439562 172170 439618 172226
rect 439686 172170 439742 172226
rect 439314 172046 439370 172102
rect 439438 172046 439494 172102
rect 439562 172046 439618 172102
rect 439686 172046 439742 172102
rect 439314 171922 439370 171978
rect 439438 171922 439494 171978
rect 439562 171922 439618 171978
rect 439686 171922 439742 171978
rect 439314 154294 439370 154350
rect 439438 154294 439494 154350
rect 439562 154294 439618 154350
rect 439686 154294 439742 154350
rect 439314 154170 439370 154226
rect 439438 154170 439494 154226
rect 439562 154170 439618 154226
rect 439686 154170 439742 154226
rect 439314 154046 439370 154102
rect 439438 154046 439494 154102
rect 439562 154046 439618 154102
rect 439686 154046 439742 154102
rect 439314 153922 439370 153978
rect 439438 153922 439494 153978
rect 439562 153922 439618 153978
rect 439686 153922 439742 153978
rect 439314 136294 439370 136350
rect 439438 136294 439494 136350
rect 439562 136294 439618 136350
rect 439686 136294 439742 136350
rect 439314 136170 439370 136226
rect 439438 136170 439494 136226
rect 439562 136170 439618 136226
rect 439686 136170 439742 136226
rect 439314 136046 439370 136102
rect 439438 136046 439494 136102
rect 439562 136046 439618 136102
rect 439686 136046 439742 136102
rect 439314 135922 439370 135978
rect 439438 135922 439494 135978
rect 439562 135922 439618 135978
rect 439686 135922 439742 135978
rect 433878 118294 433934 118350
rect 434002 118294 434058 118350
rect 433878 118170 433934 118226
rect 434002 118170 434058 118226
rect 433878 118046 433934 118102
rect 434002 118046 434058 118102
rect 433878 117922 433934 117978
rect 434002 117922 434058 117978
rect 449238 130294 449294 130350
rect 449362 130294 449418 130350
rect 449238 130170 449294 130226
rect 449362 130170 449418 130226
rect 449238 130046 449294 130102
rect 449362 130046 449418 130102
rect 449238 129922 449294 129978
rect 449362 129922 449418 129978
rect 455420 125702 455476 125758
rect 455308 123956 455364 123958
rect 455308 123902 455364 123956
rect 455308 120482 455364 120538
rect 439314 118294 439370 118350
rect 439438 118294 439494 118350
rect 439562 118294 439618 118350
rect 439686 118294 439742 118350
rect 439314 118170 439370 118226
rect 439438 118170 439494 118226
rect 439562 118170 439618 118226
rect 439686 118170 439742 118226
rect 439314 118046 439370 118102
rect 439438 118046 439494 118102
rect 439562 118046 439618 118102
rect 439686 118046 439742 118102
rect 439314 117922 439370 117978
rect 439438 117922 439494 117978
rect 439562 117922 439618 117978
rect 439686 117922 439742 117978
rect 418518 112294 418574 112350
rect 418642 112294 418698 112350
rect 418518 112170 418574 112226
rect 418642 112170 418698 112226
rect 418518 112046 418574 112102
rect 418642 112046 418698 112102
rect 418518 111922 418574 111978
rect 418642 111922 418698 111978
rect 435594 112294 435650 112350
rect 435718 112294 435774 112350
rect 435842 112294 435898 112350
rect 435966 112294 436022 112350
rect 435594 112170 435650 112226
rect 435718 112170 435774 112226
rect 435842 112170 435898 112226
rect 435966 112170 436022 112226
rect 435594 112046 435650 112102
rect 435718 112046 435774 112102
rect 435842 112046 435898 112102
rect 435966 112046 436022 112102
rect 435594 111922 435650 111978
rect 435718 111922 435774 111978
rect 435842 111922 435898 111978
rect 435966 111922 436022 111978
rect 408594 100294 408650 100350
rect 408718 100294 408774 100350
rect 408842 100294 408898 100350
rect 408966 100294 409022 100350
rect 408594 100170 408650 100226
rect 408718 100170 408774 100226
rect 408842 100170 408898 100226
rect 408966 100170 409022 100226
rect 408594 100046 408650 100102
rect 408718 100046 408774 100102
rect 408842 100046 408898 100102
rect 408966 100046 409022 100102
rect 408594 99922 408650 99978
rect 408718 99922 408774 99978
rect 408842 99922 408898 99978
rect 408966 99922 409022 99978
rect 408594 82294 408650 82350
rect 408718 82294 408774 82350
rect 408842 82294 408898 82350
rect 408966 82294 409022 82350
rect 408594 82170 408650 82226
rect 408718 82170 408774 82226
rect 408842 82170 408898 82226
rect 408966 82170 409022 82226
rect 408594 82046 408650 82102
rect 408718 82046 408774 82102
rect 408842 82046 408898 82102
rect 408966 82046 409022 82102
rect 408594 81922 408650 81978
rect 408718 81922 408774 81978
rect 408842 81922 408898 81978
rect 408966 81922 409022 81978
rect 408594 64294 408650 64350
rect 408718 64294 408774 64350
rect 408842 64294 408898 64350
rect 408966 64294 409022 64350
rect 408594 64170 408650 64226
rect 408718 64170 408774 64226
rect 408842 64170 408898 64226
rect 408966 64170 409022 64226
rect 408594 64046 408650 64102
rect 408718 64046 408774 64102
rect 408842 64046 408898 64102
rect 408966 64046 409022 64102
rect 408594 63922 408650 63978
rect 408718 63922 408774 63978
rect 408842 63922 408898 63978
rect 408966 63922 409022 63978
rect 435594 94294 435650 94350
rect 435718 94294 435774 94350
rect 435842 94294 435898 94350
rect 435966 94294 436022 94350
rect 435594 94170 435650 94226
rect 435718 94170 435774 94226
rect 435842 94170 435898 94226
rect 435966 94170 436022 94226
rect 435594 94046 435650 94102
rect 435718 94046 435774 94102
rect 435842 94046 435898 94102
rect 435966 94046 436022 94102
rect 435594 93922 435650 93978
rect 435718 93922 435774 93978
rect 435842 93922 435898 93978
rect 435966 93922 436022 93978
rect 435594 76294 435650 76350
rect 435718 76294 435774 76350
rect 435842 76294 435898 76350
rect 435966 76294 436022 76350
rect 435594 76170 435650 76226
rect 435718 76170 435774 76226
rect 435842 76170 435898 76226
rect 435966 76170 436022 76226
rect 435594 76046 435650 76102
rect 435718 76046 435774 76102
rect 435842 76046 435898 76102
rect 435966 76046 436022 76102
rect 435594 75922 435650 75978
rect 435718 75922 435774 75978
rect 435842 75922 435898 75978
rect 435966 75922 436022 75978
rect 433878 64294 433934 64350
rect 434002 64294 434058 64350
rect 433878 64170 433934 64226
rect 434002 64170 434058 64226
rect 433878 64046 433934 64102
rect 434002 64046 434058 64102
rect 433878 63922 433934 63978
rect 434002 63922 434058 63978
rect 418518 58294 418574 58350
rect 418642 58294 418698 58350
rect 418518 58170 418574 58226
rect 418642 58170 418698 58226
rect 418518 58046 418574 58102
rect 418642 58046 418698 58102
rect 418518 57922 418574 57978
rect 418642 57922 418698 57978
rect 435594 58294 435650 58350
rect 435718 58294 435774 58350
rect 435842 58294 435898 58350
rect 435966 58294 436022 58350
rect 435594 58170 435650 58226
rect 435718 58170 435774 58226
rect 435842 58170 435898 58226
rect 435966 58170 436022 58226
rect 435594 58046 435650 58102
rect 435718 58046 435774 58102
rect 435842 58046 435898 58102
rect 435966 58046 436022 58102
rect 435594 57922 435650 57978
rect 435718 57922 435774 57978
rect 435842 57922 435898 57978
rect 435966 57922 436022 57978
rect 414652 56252 414708 56278
rect 414652 56222 414708 56252
rect 456988 133442 457044 133498
rect 466314 166294 466370 166350
rect 466438 166294 466494 166350
rect 466562 166294 466618 166350
rect 466686 166294 466742 166350
rect 466314 166170 466370 166226
rect 466438 166170 466494 166226
rect 466562 166170 466618 166226
rect 466686 166170 466742 166226
rect 466314 166046 466370 166102
rect 466438 166046 466494 166102
rect 466562 166046 466618 166102
rect 466686 166046 466742 166102
rect 466314 165922 466370 165978
rect 466438 165922 466494 165978
rect 466562 165922 466618 165978
rect 466686 165922 466742 165978
rect 466314 148294 466370 148350
rect 466438 148294 466494 148350
rect 466562 148294 466618 148350
rect 466686 148294 466742 148350
rect 466314 148170 466370 148226
rect 466438 148170 466494 148226
rect 466562 148170 466618 148226
rect 466686 148170 466742 148226
rect 466314 148046 466370 148102
rect 466438 148046 466494 148102
rect 466562 148046 466618 148102
rect 466686 148046 466742 148102
rect 466314 147922 466370 147978
rect 466438 147922 466494 147978
rect 466562 147922 466618 147978
rect 466686 147922 466742 147978
rect 466314 130294 466370 130350
rect 466438 130294 466494 130350
rect 466562 130294 466618 130350
rect 466686 130294 466742 130350
rect 466314 130170 466370 130226
rect 466438 130170 466494 130226
rect 466562 130170 466618 130226
rect 466686 130170 466742 130226
rect 466314 130046 466370 130102
rect 466438 130046 466494 130102
rect 466562 130046 466618 130102
rect 466686 130046 466742 130102
rect 466314 129922 466370 129978
rect 466438 129922 466494 129978
rect 466562 129922 466618 129978
rect 466686 129922 466742 129978
rect 449238 112294 449294 112350
rect 449362 112294 449418 112350
rect 449238 112170 449294 112226
rect 449362 112170 449418 112226
rect 449238 112046 449294 112102
rect 449362 112046 449418 112102
rect 449238 111922 449294 111978
rect 449362 111922 449418 111978
rect 466314 112294 466370 112350
rect 466438 112294 466494 112350
rect 466562 112294 466618 112350
rect 466686 112294 466742 112350
rect 466314 112170 466370 112226
rect 466438 112170 466494 112226
rect 466562 112170 466618 112226
rect 466686 112170 466742 112226
rect 466314 112046 466370 112102
rect 466438 112046 466494 112102
rect 466562 112046 466618 112102
rect 466686 112046 466742 112102
rect 466314 111922 466370 111978
rect 466438 111922 466494 111978
rect 466562 111922 466618 111978
rect 466686 111922 466742 111978
rect 439314 100294 439370 100350
rect 439438 100294 439494 100350
rect 439562 100294 439618 100350
rect 439686 100294 439742 100350
rect 439314 100170 439370 100226
rect 439438 100170 439494 100226
rect 439562 100170 439618 100226
rect 439686 100170 439742 100226
rect 439314 100046 439370 100102
rect 439438 100046 439494 100102
rect 439562 100046 439618 100102
rect 439686 100046 439742 100102
rect 439314 99922 439370 99978
rect 439438 99922 439494 99978
rect 439562 99922 439618 99978
rect 439686 99922 439742 99978
rect 439314 82294 439370 82350
rect 439438 82294 439494 82350
rect 439562 82294 439618 82350
rect 439686 82294 439742 82350
rect 439314 82170 439370 82226
rect 439438 82170 439494 82226
rect 439562 82170 439618 82226
rect 439686 82170 439742 82226
rect 439314 82046 439370 82102
rect 439438 82046 439494 82102
rect 439562 82046 439618 82102
rect 439686 82046 439742 82102
rect 439314 81922 439370 81978
rect 439438 81922 439494 81978
rect 439562 81922 439618 81978
rect 439686 81922 439742 81978
rect 439314 64294 439370 64350
rect 439438 64294 439494 64350
rect 439562 64294 439618 64350
rect 439686 64294 439742 64350
rect 439314 64170 439370 64226
rect 439438 64170 439494 64226
rect 439562 64170 439618 64226
rect 439686 64170 439742 64226
rect 439314 64046 439370 64102
rect 439438 64046 439494 64102
rect 439562 64046 439618 64102
rect 439686 64046 439742 64102
rect 439314 63922 439370 63978
rect 439438 63922 439494 63978
rect 439562 63922 439618 63978
rect 439686 63922 439742 63978
rect 408594 46294 408650 46350
rect 408718 46294 408774 46350
rect 408842 46294 408898 46350
rect 408966 46294 409022 46350
rect 408594 46170 408650 46226
rect 408718 46170 408774 46226
rect 408842 46170 408898 46226
rect 408966 46170 409022 46226
rect 408594 46046 408650 46102
rect 408718 46046 408774 46102
rect 408842 46046 408898 46102
rect 408966 46046 409022 46102
rect 408594 45922 408650 45978
rect 408718 45922 408774 45978
rect 408842 45922 408898 45978
rect 408966 45922 409022 45978
rect 433878 46294 433934 46350
rect 434002 46294 434058 46350
rect 433878 46170 433934 46226
rect 434002 46170 434058 46226
rect 433878 46046 433934 46102
rect 434002 46046 434058 46102
rect 433878 45922 433934 45978
rect 434002 45922 434058 45978
rect 449238 58294 449294 58350
rect 449362 58294 449418 58350
rect 449238 58170 449294 58226
rect 449362 58170 449418 58226
rect 449238 58046 449294 58102
rect 449362 58046 449418 58102
rect 449238 57922 449294 57978
rect 449362 57922 449418 57978
rect 466314 94294 466370 94350
rect 466438 94294 466494 94350
rect 466562 94294 466618 94350
rect 466686 94294 466742 94350
rect 466314 94170 466370 94226
rect 466438 94170 466494 94226
rect 466562 94170 466618 94226
rect 466686 94170 466742 94226
rect 466314 94046 466370 94102
rect 466438 94046 466494 94102
rect 466562 94046 466618 94102
rect 466686 94046 466742 94102
rect 466314 93922 466370 93978
rect 466438 93922 466494 93978
rect 466562 93922 466618 93978
rect 466686 93922 466742 93978
rect 466314 76294 466370 76350
rect 466438 76294 466494 76350
rect 466562 76294 466618 76350
rect 466686 76294 466742 76350
rect 466314 76170 466370 76226
rect 466438 76170 466494 76226
rect 466562 76170 466618 76226
rect 466686 76170 466742 76226
rect 466314 76046 466370 76102
rect 466438 76046 466494 76102
rect 466562 76046 466618 76102
rect 466686 76046 466742 76102
rect 466314 75922 466370 75978
rect 466438 75922 466494 75978
rect 466562 75922 466618 75978
rect 466686 75922 466742 75978
rect 466314 58294 466370 58350
rect 466438 58294 466494 58350
rect 466562 58294 466618 58350
rect 466686 58294 466742 58350
rect 466314 58170 466370 58226
rect 466438 58170 466494 58226
rect 466562 58170 466618 58226
rect 466686 58170 466742 58226
rect 466314 58046 466370 58102
rect 466438 58046 466494 58102
rect 466562 58046 466618 58102
rect 466686 58046 466742 58102
rect 466314 57922 466370 57978
rect 466438 57922 466494 57978
rect 466562 57922 466618 57978
rect 466686 57922 466742 57978
rect 439314 46294 439370 46350
rect 439438 46294 439494 46350
rect 439562 46294 439618 46350
rect 439686 46294 439742 46350
rect 439314 46170 439370 46226
rect 439438 46170 439494 46226
rect 439562 46170 439618 46226
rect 439686 46170 439742 46226
rect 439314 46046 439370 46102
rect 439438 46046 439494 46102
rect 439562 46046 439618 46102
rect 439686 46046 439742 46102
rect 439314 45922 439370 45978
rect 439438 45922 439494 45978
rect 439562 45922 439618 45978
rect 439686 45922 439742 45978
rect 418518 40294 418574 40350
rect 418642 40294 418698 40350
rect 418518 40170 418574 40226
rect 418642 40170 418698 40226
rect 418518 40046 418574 40102
rect 418642 40046 418698 40102
rect 418518 39922 418574 39978
rect 418642 39922 418698 39978
rect 435594 40294 435650 40350
rect 435718 40294 435774 40350
rect 435842 40294 435898 40350
rect 435966 40294 436022 40350
rect 435594 40170 435650 40226
rect 435718 40170 435774 40226
rect 435842 40170 435898 40226
rect 435966 40170 436022 40226
rect 435594 40046 435650 40102
rect 435718 40046 435774 40102
rect 435842 40046 435898 40102
rect 435966 40046 436022 40102
rect 435594 39922 435650 39978
rect 435718 39922 435774 39978
rect 435842 39922 435898 39978
rect 435966 39922 436022 39978
rect 408594 28294 408650 28350
rect 408718 28294 408774 28350
rect 408842 28294 408898 28350
rect 408966 28294 409022 28350
rect 408594 28170 408650 28226
rect 408718 28170 408774 28226
rect 408842 28170 408898 28226
rect 408966 28170 409022 28226
rect 408594 28046 408650 28102
rect 408718 28046 408774 28102
rect 408842 28046 408898 28102
rect 408966 28046 409022 28102
rect 408594 27922 408650 27978
rect 408718 27922 408774 27978
rect 408842 27922 408898 27978
rect 408966 27922 409022 27978
rect 408594 10294 408650 10350
rect 408718 10294 408774 10350
rect 408842 10294 408898 10350
rect 408966 10294 409022 10350
rect 408594 10170 408650 10226
rect 408718 10170 408774 10226
rect 408842 10170 408898 10226
rect 408966 10170 409022 10226
rect 408594 10046 408650 10102
rect 408718 10046 408774 10102
rect 408842 10046 408898 10102
rect 408966 10046 409022 10102
rect 408594 9922 408650 9978
rect 408718 9922 408774 9978
rect 408842 9922 408898 9978
rect 408966 9922 409022 9978
rect 408594 -1176 408650 -1120
rect 408718 -1176 408774 -1120
rect 408842 -1176 408898 -1120
rect 408966 -1176 409022 -1120
rect 408594 -1300 408650 -1244
rect 408718 -1300 408774 -1244
rect 408842 -1300 408898 -1244
rect 408966 -1300 409022 -1244
rect 408594 -1424 408650 -1368
rect 408718 -1424 408774 -1368
rect 408842 -1424 408898 -1368
rect 408966 -1424 409022 -1368
rect 408594 -1548 408650 -1492
rect 408718 -1548 408774 -1492
rect 408842 -1548 408898 -1492
rect 408966 -1548 409022 -1492
rect 435594 22294 435650 22350
rect 435718 22294 435774 22350
rect 435842 22294 435898 22350
rect 435966 22294 436022 22350
rect 435594 22170 435650 22226
rect 435718 22170 435774 22226
rect 435842 22170 435898 22226
rect 435966 22170 436022 22226
rect 435594 22046 435650 22102
rect 435718 22046 435774 22102
rect 435842 22046 435898 22102
rect 435966 22046 436022 22102
rect 435594 21922 435650 21978
rect 435718 21922 435774 21978
rect 435842 21922 435898 21978
rect 435966 21922 436022 21978
rect 435594 4294 435650 4350
rect 435718 4294 435774 4350
rect 435842 4294 435898 4350
rect 435966 4294 436022 4350
rect 435594 4170 435650 4226
rect 435718 4170 435774 4226
rect 435842 4170 435898 4226
rect 435966 4170 436022 4226
rect 435594 4046 435650 4102
rect 435718 4046 435774 4102
rect 435842 4046 435898 4102
rect 435966 4046 436022 4102
rect 435594 3922 435650 3978
rect 435718 3922 435774 3978
rect 435842 3922 435898 3978
rect 435966 3922 436022 3978
rect 435594 -216 435650 -160
rect 435718 -216 435774 -160
rect 435842 -216 435898 -160
rect 435966 -216 436022 -160
rect 435594 -340 435650 -284
rect 435718 -340 435774 -284
rect 435842 -340 435898 -284
rect 435966 -340 436022 -284
rect 435594 -464 435650 -408
rect 435718 -464 435774 -408
rect 435842 -464 435898 -408
rect 435966 -464 436022 -408
rect 435594 -588 435650 -532
rect 435718 -588 435774 -532
rect 435842 -588 435898 -532
rect 435966 -588 436022 -532
rect 449238 40294 449294 40350
rect 449362 40294 449418 40350
rect 449238 40170 449294 40226
rect 449362 40170 449418 40226
rect 449238 40046 449294 40102
rect 449362 40046 449418 40102
rect 449238 39922 449294 39978
rect 449362 39922 449418 39978
rect 466314 40294 466370 40350
rect 466438 40294 466494 40350
rect 466562 40294 466618 40350
rect 466686 40294 466742 40350
rect 466314 40170 466370 40226
rect 466438 40170 466494 40226
rect 466562 40170 466618 40226
rect 466686 40170 466742 40226
rect 466314 40046 466370 40102
rect 466438 40046 466494 40102
rect 466562 40046 466618 40102
rect 466686 40046 466742 40102
rect 466314 39922 466370 39978
rect 466438 39922 466494 39978
rect 466562 39922 466618 39978
rect 466686 39922 466742 39978
rect 439314 28294 439370 28350
rect 439438 28294 439494 28350
rect 439562 28294 439618 28350
rect 439686 28294 439742 28350
rect 439314 28170 439370 28226
rect 439438 28170 439494 28226
rect 439562 28170 439618 28226
rect 439686 28170 439742 28226
rect 439314 28046 439370 28102
rect 439438 28046 439494 28102
rect 439562 28046 439618 28102
rect 439686 28046 439742 28102
rect 439314 27922 439370 27978
rect 439438 27922 439494 27978
rect 439562 27922 439618 27978
rect 439686 27922 439742 27978
rect 439314 10294 439370 10350
rect 439438 10294 439494 10350
rect 439562 10294 439618 10350
rect 439686 10294 439742 10350
rect 439314 10170 439370 10226
rect 439438 10170 439494 10226
rect 439562 10170 439618 10226
rect 439686 10170 439742 10226
rect 439314 10046 439370 10102
rect 439438 10046 439494 10102
rect 439562 10046 439618 10102
rect 439686 10046 439742 10102
rect 439314 9922 439370 9978
rect 439438 9922 439494 9978
rect 439562 9922 439618 9978
rect 439686 9922 439742 9978
rect 439314 -1176 439370 -1120
rect 439438 -1176 439494 -1120
rect 439562 -1176 439618 -1120
rect 439686 -1176 439742 -1120
rect 439314 -1300 439370 -1244
rect 439438 -1300 439494 -1244
rect 439562 -1300 439618 -1244
rect 439686 -1300 439742 -1244
rect 439314 -1424 439370 -1368
rect 439438 -1424 439494 -1368
rect 439562 -1424 439618 -1368
rect 439686 -1424 439742 -1368
rect 439314 -1548 439370 -1492
rect 439438 -1548 439494 -1492
rect 439562 -1548 439618 -1492
rect 439686 -1548 439742 -1492
rect 466314 22294 466370 22350
rect 466438 22294 466494 22350
rect 466562 22294 466618 22350
rect 466686 22294 466742 22350
rect 466314 22170 466370 22226
rect 466438 22170 466494 22226
rect 466562 22170 466618 22226
rect 466686 22170 466742 22226
rect 466314 22046 466370 22102
rect 466438 22046 466494 22102
rect 466562 22046 466618 22102
rect 466686 22046 466742 22102
rect 466314 21922 466370 21978
rect 466438 21922 466494 21978
rect 466562 21922 466618 21978
rect 466686 21922 466742 21978
rect 466314 4294 466370 4350
rect 466438 4294 466494 4350
rect 466562 4294 466618 4350
rect 466686 4294 466742 4350
rect 466314 4170 466370 4226
rect 466438 4170 466494 4226
rect 466562 4170 466618 4226
rect 466686 4170 466742 4226
rect 466314 4046 466370 4102
rect 466438 4046 466494 4102
rect 466562 4046 466618 4102
rect 466686 4046 466742 4102
rect 466314 3922 466370 3978
rect 466438 3922 466494 3978
rect 466562 3922 466618 3978
rect 466686 3922 466742 3978
rect 466314 -216 466370 -160
rect 466438 -216 466494 -160
rect 466562 -216 466618 -160
rect 466686 -216 466742 -160
rect 466314 -340 466370 -284
rect 466438 -340 466494 -284
rect 466562 -340 466618 -284
rect 466686 -340 466742 -284
rect 466314 -464 466370 -408
rect 466438 -464 466494 -408
rect 466562 -464 466618 -408
rect 466686 -464 466742 -408
rect 466314 -588 466370 -532
rect 466438 -588 466494 -532
rect 466562 -588 466618 -532
rect 466686 -588 466742 -532
rect 495878 208294 495934 208350
rect 496002 208294 496058 208350
rect 495878 208170 495934 208226
rect 496002 208170 496058 208226
rect 495878 208046 495934 208102
rect 496002 208046 496058 208102
rect 495878 207922 495934 207978
rect 496002 207922 496058 207978
rect 480518 202294 480574 202350
rect 480642 202294 480698 202350
rect 480518 202170 480574 202226
rect 480642 202170 480698 202226
rect 480518 202046 480574 202102
rect 480642 202046 480698 202102
rect 480518 201922 480574 201978
rect 480642 201922 480698 201978
rect 497034 202294 497090 202350
rect 497158 202294 497214 202350
rect 497282 202294 497338 202350
rect 497406 202294 497462 202350
rect 497034 202170 497090 202226
rect 497158 202170 497214 202226
rect 497282 202170 497338 202226
rect 497406 202170 497462 202226
rect 497034 202046 497090 202102
rect 497158 202046 497214 202102
rect 497282 202046 497338 202102
rect 497406 202046 497462 202102
rect 497034 201922 497090 201978
rect 497158 201922 497214 201978
rect 497282 201922 497338 201978
rect 497406 201922 497462 201978
rect 473676 198242 473732 198298
rect 472108 195722 472164 195778
rect 470034 190294 470090 190350
rect 470158 190294 470214 190350
rect 470282 190294 470338 190350
rect 470406 190294 470462 190350
rect 470034 190170 470090 190226
rect 470158 190170 470214 190226
rect 470282 190170 470338 190226
rect 470406 190170 470462 190226
rect 470034 190046 470090 190102
rect 470158 190046 470214 190102
rect 470282 190046 470338 190102
rect 470406 190046 470462 190102
rect 470034 189922 470090 189978
rect 470158 189922 470214 189978
rect 470282 189922 470338 189978
rect 470406 189922 470462 189978
rect 495878 190294 495934 190350
rect 496002 190294 496058 190350
rect 495878 190170 495934 190226
rect 496002 190170 496058 190226
rect 495878 190046 495934 190102
rect 496002 190046 496058 190102
rect 495878 189922 495934 189978
rect 496002 189922 496058 189978
rect 472108 189602 472164 189658
rect 472108 187982 472164 188038
rect 480518 184294 480574 184350
rect 480642 184294 480698 184350
rect 480518 184170 480574 184226
rect 480642 184170 480698 184226
rect 480518 184046 480574 184102
rect 480642 184046 480698 184102
rect 480518 183922 480574 183978
rect 480642 183922 480698 183978
rect 497034 184294 497090 184350
rect 497158 184294 497214 184350
rect 497282 184294 497338 184350
rect 497406 184294 497462 184350
rect 497034 184170 497090 184226
rect 497158 184170 497214 184226
rect 497282 184170 497338 184226
rect 497406 184170 497462 184226
rect 497034 184046 497090 184102
rect 497158 184046 497214 184102
rect 497282 184046 497338 184102
rect 497406 184046 497462 184102
rect 497034 183922 497090 183978
rect 497158 183922 497214 183978
rect 497282 183922 497338 183978
rect 497406 183922 497462 183978
rect 470034 172294 470090 172350
rect 470158 172294 470214 172350
rect 470282 172294 470338 172350
rect 470406 172294 470462 172350
rect 470034 172170 470090 172226
rect 470158 172170 470214 172226
rect 470282 172170 470338 172226
rect 470406 172170 470462 172226
rect 470034 172046 470090 172102
rect 470158 172046 470214 172102
rect 470282 172046 470338 172102
rect 470406 172046 470462 172102
rect 470034 171922 470090 171978
rect 470158 171922 470214 171978
rect 470282 171922 470338 171978
rect 470406 171922 470462 171978
rect 470034 154294 470090 154350
rect 470158 154294 470214 154350
rect 470282 154294 470338 154350
rect 470406 154294 470462 154350
rect 470034 154170 470090 154226
rect 470158 154170 470214 154226
rect 470282 154170 470338 154226
rect 470406 154170 470462 154226
rect 470034 154046 470090 154102
rect 470158 154046 470214 154102
rect 470282 154046 470338 154102
rect 470406 154046 470462 154102
rect 470034 153922 470090 153978
rect 470158 153922 470214 153978
rect 470282 153922 470338 153978
rect 470406 153922 470462 153978
rect 497034 166294 497090 166350
rect 497158 166294 497214 166350
rect 497282 166294 497338 166350
rect 497406 166294 497462 166350
rect 497034 166170 497090 166226
rect 497158 166170 497214 166226
rect 497282 166170 497338 166226
rect 497406 166170 497462 166226
rect 497034 166046 497090 166102
rect 497158 166046 497214 166102
rect 497282 166046 497338 166102
rect 497406 166046 497462 166102
rect 497034 165922 497090 165978
rect 497158 165922 497214 165978
rect 497282 165922 497338 165978
rect 497406 165922 497462 165978
rect 470034 136294 470090 136350
rect 470158 136294 470214 136350
rect 470282 136294 470338 136350
rect 470406 136294 470462 136350
rect 470034 136170 470090 136226
rect 470158 136170 470214 136226
rect 470282 136170 470338 136226
rect 470406 136170 470462 136226
rect 470034 136046 470090 136102
rect 470158 136046 470214 136102
rect 470282 136046 470338 136102
rect 470406 136046 470462 136102
rect 470034 135922 470090 135978
rect 470158 135922 470214 135978
rect 470282 135922 470338 135978
rect 470406 135922 470462 135978
rect 470034 118294 470090 118350
rect 470158 118294 470214 118350
rect 470282 118294 470338 118350
rect 470406 118294 470462 118350
rect 470034 118170 470090 118226
rect 470158 118170 470214 118226
rect 470282 118170 470338 118226
rect 470406 118170 470462 118226
rect 470034 118046 470090 118102
rect 470158 118046 470214 118102
rect 470282 118046 470338 118102
rect 470406 118046 470462 118102
rect 470034 117922 470090 117978
rect 470158 117922 470214 117978
rect 470282 117922 470338 117978
rect 470406 117922 470462 117978
rect 497034 148294 497090 148350
rect 497158 148294 497214 148350
rect 497282 148294 497338 148350
rect 497406 148294 497462 148350
rect 497034 148170 497090 148226
rect 497158 148170 497214 148226
rect 497282 148170 497338 148226
rect 497406 148170 497462 148226
rect 497034 148046 497090 148102
rect 497158 148046 497214 148102
rect 497282 148046 497338 148102
rect 497406 148046 497462 148102
rect 497034 147922 497090 147978
rect 497158 147922 497214 147978
rect 497282 147922 497338 147978
rect 497406 147922 497462 147978
rect 495878 136294 495934 136350
rect 496002 136294 496058 136350
rect 495878 136170 495934 136226
rect 496002 136170 496058 136226
rect 495878 136046 495934 136102
rect 496002 136046 496058 136102
rect 495878 135922 495934 135978
rect 496002 135922 496058 135978
rect 480518 130294 480574 130350
rect 480642 130294 480698 130350
rect 480518 130170 480574 130226
rect 480642 130170 480698 130226
rect 480518 130046 480574 130102
rect 480642 130046 480698 130102
rect 480518 129922 480574 129978
rect 480642 129922 480698 129978
rect 497034 130294 497090 130350
rect 497158 130294 497214 130350
rect 497282 130294 497338 130350
rect 497406 130294 497462 130350
rect 497034 130170 497090 130226
rect 497158 130170 497214 130226
rect 497282 130170 497338 130226
rect 497406 130170 497462 130226
rect 497034 130046 497090 130102
rect 497158 130046 497214 130102
rect 497282 130046 497338 130102
rect 497406 130046 497462 130102
rect 497034 129922 497090 129978
rect 497158 129922 497214 129978
rect 497282 129922 497338 129978
rect 497406 129922 497462 129978
rect 473676 128402 473732 128458
rect 476028 127862 476084 127918
rect 500754 262294 500810 262350
rect 500878 262294 500934 262350
rect 501002 262294 501058 262350
rect 501126 262294 501182 262350
rect 500754 262170 500810 262226
rect 500878 262170 500934 262226
rect 501002 262170 501058 262226
rect 501126 262170 501182 262226
rect 500754 262046 500810 262102
rect 500878 262046 500934 262102
rect 501002 262046 501058 262102
rect 501126 262046 501182 262102
rect 500754 261922 500810 261978
rect 500878 261922 500934 261978
rect 501002 261922 501058 261978
rect 501126 261922 501182 261978
rect 527754 292294 527810 292350
rect 527878 292294 527934 292350
rect 528002 292294 528058 292350
rect 528126 292294 528182 292350
rect 527754 292170 527810 292226
rect 527878 292170 527934 292226
rect 528002 292170 528058 292226
rect 528126 292170 528182 292226
rect 527754 292046 527810 292102
rect 527878 292046 527934 292102
rect 528002 292046 528058 292102
rect 528126 292046 528182 292102
rect 527754 291922 527810 291978
rect 527878 291922 527934 291978
rect 528002 291922 528058 291978
rect 528126 291922 528182 291978
rect 527754 274294 527810 274350
rect 527878 274294 527934 274350
rect 528002 274294 528058 274350
rect 528126 274294 528182 274350
rect 527754 274170 527810 274226
rect 527878 274170 527934 274226
rect 528002 274170 528058 274226
rect 528126 274170 528182 274226
rect 527754 274046 527810 274102
rect 527878 274046 527934 274102
rect 528002 274046 528058 274102
rect 528126 274046 528182 274102
rect 527754 273922 527810 273978
rect 527878 273922 527934 273978
rect 528002 273922 528058 273978
rect 528126 273922 528182 273978
rect 517468 258182 517524 258238
rect 511238 256294 511294 256350
rect 511362 256294 511418 256350
rect 511238 256170 511294 256226
rect 511362 256170 511418 256226
rect 511238 256046 511294 256102
rect 511362 256046 511418 256102
rect 511238 255922 511294 255978
rect 511362 255922 511418 255978
rect 527754 256294 527810 256350
rect 527878 256294 527934 256350
rect 528002 256294 528058 256350
rect 528126 256294 528182 256350
rect 527754 256170 527810 256226
rect 527878 256170 527934 256226
rect 528002 256170 528058 256226
rect 528126 256170 528182 256226
rect 527754 256046 527810 256102
rect 527878 256046 527934 256102
rect 528002 256046 528058 256102
rect 528126 256046 528182 256102
rect 527754 255922 527810 255978
rect 527878 255922 527934 255978
rect 528002 255922 528058 255978
rect 528126 255922 528182 255978
rect 500754 244294 500810 244350
rect 500878 244294 500934 244350
rect 501002 244294 501058 244350
rect 501126 244294 501182 244350
rect 500754 244170 500810 244226
rect 500878 244170 500934 244226
rect 501002 244170 501058 244226
rect 501126 244170 501182 244226
rect 500754 244046 500810 244102
rect 500878 244046 500934 244102
rect 501002 244046 501058 244102
rect 501126 244046 501182 244102
rect 500754 243922 500810 243978
rect 500878 243922 500934 243978
rect 501002 243922 501058 243978
rect 501126 243922 501182 243978
rect 527754 238294 527810 238350
rect 527878 238294 527934 238350
rect 528002 238294 528058 238350
rect 528126 238294 528182 238350
rect 527754 238170 527810 238226
rect 527878 238170 527934 238226
rect 528002 238170 528058 238226
rect 528126 238170 528182 238226
rect 527754 238046 527810 238102
rect 527878 238046 527934 238102
rect 528002 238046 528058 238102
rect 528126 238046 528182 238102
rect 527754 237922 527810 237978
rect 527878 237922 527934 237978
rect 528002 237922 528058 237978
rect 528126 237922 528182 237978
rect 500754 226294 500810 226350
rect 500878 226294 500934 226350
rect 501002 226294 501058 226350
rect 501126 226294 501182 226350
rect 500754 226170 500810 226226
rect 500878 226170 500934 226226
rect 501002 226170 501058 226226
rect 501126 226170 501182 226226
rect 500754 226046 500810 226102
rect 500878 226046 500934 226102
rect 501002 226046 501058 226102
rect 501126 226046 501182 226102
rect 500754 225922 500810 225978
rect 500878 225922 500934 225978
rect 501002 225922 501058 225978
rect 501126 225922 501182 225978
rect 500754 208294 500810 208350
rect 500878 208294 500934 208350
rect 501002 208294 501058 208350
rect 501126 208294 501182 208350
rect 500754 208170 500810 208226
rect 500878 208170 500934 208226
rect 501002 208170 501058 208226
rect 501126 208170 501182 208226
rect 500754 208046 500810 208102
rect 500878 208046 500934 208102
rect 501002 208046 501058 208102
rect 501126 208046 501182 208102
rect 500754 207922 500810 207978
rect 500878 207922 500934 207978
rect 501002 207922 501058 207978
rect 501126 207922 501182 207978
rect 511238 202294 511294 202350
rect 511362 202294 511418 202350
rect 511238 202170 511294 202226
rect 511362 202170 511418 202226
rect 511238 202046 511294 202102
rect 511362 202046 511418 202102
rect 511238 201922 511294 201978
rect 511362 201922 511418 201978
rect 500754 190294 500810 190350
rect 500878 190294 500934 190350
rect 501002 190294 501058 190350
rect 501126 190294 501182 190350
rect 500754 190170 500810 190226
rect 500878 190170 500934 190226
rect 501002 190170 501058 190226
rect 501126 190170 501182 190226
rect 500754 190046 500810 190102
rect 500878 190046 500934 190102
rect 501002 190046 501058 190102
rect 501126 190046 501182 190102
rect 500754 189922 500810 189978
rect 500878 189922 500934 189978
rect 501002 189922 501058 189978
rect 501126 189922 501182 189978
rect 511238 184294 511294 184350
rect 511362 184294 511418 184350
rect 511238 184170 511294 184226
rect 511362 184170 511418 184226
rect 511238 184046 511294 184102
rect 511362 184046 511418 184102
rect 511238 183922 511294 183978
rect 511362 183922 511418 183978
rect 519148 200762 519204 200818
rect 527754 220294 527810 220350
rect 527878 220294 527934 220350
rect 528002 220294 528058 220350
rect 528126 220294 528182 220350
rect 527754 220170 527810 220226
rect 527878 220170 527934 220226
rect 528002 220170 528058 220226
rect 528126 220170 528182 220226
rect 527754 220046 527810 220102
rect 527878 220046 527934 220102
rect 528002 220046 528058 220102
rect 528126 220046 528182 220102
rect 527754 219922 527810 219978
rect 527878 219922 527934 219978
rect 528002 219922 528058 219978
rect 528126 219922 528182 219978
rect 526652 205082 526708 205138
rect 524972 203282 525028 203338
rect 526652 192302 526708 192358
rect 527754 202294 527810 202350
rect 527878 202294 527934 202350
rect 528002 202294 528058 202350
rect 528126 202294 528182 202350
rect 527754 202170 527810 202226
rect 527878 202170 527934 202226
rect 528002 202170 528058 202226
rect 528126 202170 528182 202226
rect 527754 202046 527810 202102
rect 527878 202046 527934 202102
rect 528002 202046 528058 202102
rect 528126 202046 528182 202102
rect 527754 201922 527810 201978
rect 527878 201922 527934 201978
rect 528002 201922 528058 201978
rect 528126 201922 528182 201978
rect 527754 184294 527810 184350
rect 527878 184294 527934 184350
rect 528002 184294 528058 184350
rect 528126 184294 528182 184350
rect 527754 184170 527810 184226
rect 527878 184170 527934 184226
rect 528002 184170 528058 184226
rect 528126 184170 528182 184226
rect 527754 184046 527810 184102
rect 527878 184046 527934 184102
rect 528002 184046 528058 184102
rect 528126 184046 528182 184102
rect 527754 183922 527810 183978
rect 527878 183922 527934 183978
rect 528002 183922 528058 183978
rect 528126 183922 528182 183978
rect 500754 172294 500810 172350
rect 500878 172294 500934 172350
rect 501002 172294 501058 172350
rect 501126 172294 501182 172350
rect 500754 172170 500810 172226
rect 500878 172170 500934 172226
rect 501002 172170 501058 172226
rect 501126 172170 501182 172226
rect 500754 172046 500810 172102
rect 500878 172046 500934 172102
rect 501002 172046 501058 172102
rect 501126 172046 501182 172102
rect 500754 171922 500810 171978
rect 500878 171922 500934 171978
rect 501002 171922 501058 171978
rect 501126 171922 501182 171978
rect 500754 154294 500810 154350
rect 500878 154294 500934 154350
rect 501002 154294 501058 154350
rect 501126 154294 501182 154350
rect 500754 154170 500810 154226
rect 500878 154170 500934 154226
rect 501002 154170 501058 154226
rect 501126 154170 501182 154226
rect 500754 154046 500810 154102
rect 500878 154046 500934 154102
rect 501002 154046 501058 154102
rect 501126 154046 501182 154102
rect 500754 153922 500810 153978
rect 500878 153922 500934 153978
rect 501002 153922 501058 153978
rect 501126 153922 501182 153978
rect 500754 136294 500810 136350
rect 500878 136294 500934 136350
rect 501002 136294 501058 136350
rect 501126 136294 501182 136350
rect 500754 136170 500810 136226
rect 500878 136170 500934 136226
rect 501002 136170 501058 136226
rect 501126 136170 501182 136226
rect 500754 136046 500810 136102
rect 500878 136046 500934 136102
rect 501002 136046 501058 136102
rect 501126 136046 501182 136102
rect 500754 135922 500810 135978
rect 500878 135922 500934 135978
rect 501002 135922 501058 135978
rect 501126 135922 501182 135978
rect 495878 118294 495934 118350
rect 496002 118294 496058 118350
rect 495878 118170 495934 118226
rect 496002 118170 496058 118226
rect 495878 118046 495934 118102
rect 496002 118046 496058 118102
rect 495878 117922 495934 117978
rect 496002 117922 496058 117978
rect 511238 130294 511294 130350
rect 511362 130294 511418 130350
rect 511238 130170 511294 130226
rect 511362 130170 511418 130226
rect 511238 130046 511294 130102
rect 511362 130046 511418 130102
rect 511238 129922 511294 129978
rect 511362 129922 511418 129978
rect 500754 118294 500810 118350
rect 500878 118294 500934 118350
rect 501002 118294 501058 118350
rect 501126 118294 501182 118350
rect 500754 118170 500810 118226
rect 500878 118170 500934 118226
rect 501002 118170 501058 118226
rect 501126 118170 501182 118226
rect 500754 118046 500810 118102
rect 500878 118046 500934 118102
rect 501002 118046 501058 118102
rect 501126 118046 501182 118102
rect 500754 117922 500810 117978
rect 500878 117922 500934 117978
rect 501002 117922 501058 117978
rect 501126 117922 501182 117978
rect 480518 112294 480574 112350
rect 480642 112294 480698 112350
rect 480518 112170 480574 112226
rect 480642 112170 480698 112226
rect 480518 112046 480574 112102
rect 480642 112046 480698 112102
rect 480518 111922 480574 111978
rect 480642 111922 480698 111978
rect 497034 112294 497090 112350
rect 497158 112294 497214 112350
rect 497282 112294 497338 112350
rect 497406 112294 497462 112350
rect 497034 112170 497090 112226
rect 497158 112170 497214 112226
rect 497282 112170 497338 112226
rect 497406 112170 497462 112226
rect 497034 112046 497090 112102
rect 497158 112046 497214 112102
rect 497282 112046 497338 112102
rect 497406 112046 497462 112102
rect 497034 111922 497090 111978
rect 497158 111922 497214 111978
rect 497282 111922 497338 111978
rect 497406 111922 497462 111978
rect 470034 100294 470090 100350
rect 470158 100294 470214 100350
rect 470282 100294 470338 100350
rect 470406 100294 470462 100350
rect 470034 100170 470090 100226
rect 470158 100170 470214 100226
rect 470282 100170 470338 100226
rect 470406 100170 470462 100226
rect 470034 100046 470090 100102
rect 470158 100046 470214 100102
rect 470282 100046 470338 100102
rect 470406 100046 470462 100102
rect 470034 99922 470090 99978
rect 470158 99922 470214 99978
rect 470282 99922 470338 99978
rect 470406 99922 470462 99978
rect 497034 94294 497090 94350
rect 497158 94294 497214 94350
rect 497282 94294 497338 94350
rect 497406 94294 497462 94350
rect 497034 94170 497090 94226
rect 497158 94170 497214 94226
rect 497282 94170 497338 94226
rect 497406 94170 497462 94226
rect 497034 94046 497090 94102
rect 497158 94046 497214 94102
rect 497282 94046 497338 94102
rect 497406 94046 497462 94102
rect 497034 93922 497090 93978
rect 497158 93922 497214 93978
rect 497282 93922 497338 93978
rect 497406 93922 497462 93978
rect 470034 82294 470090 82350
rect 470158 82294 470214 82350
rect 470282 82294 470338 82350
rect 470406 82294 470462 82350
rect 470034 82170 470090 82226
rect 470158 82170 470214 82226
rect 470282 82170 470338 82226
rect 470406 82170 470462 82226
rect 470034 82046 470090 82102
rect 470158 82046 470214 82102
rect 470282 82046 470338 82102
rect 470406 82046 470462 82102
rect 470034 81922 470090 81978
rect 470158 81922 470214 81978
rect 470282 81922 470338 81978
rect 470406 81922 470462 81978
rect 470034 64294 470090 64350
rect 470158 64294 470214 64350
rect 470282 64294 470338 64350
rect 470406 64294 470462 64350
rect 470034 64170 470090 64226
rect 470158 64170 470214 64226
rect 470282 64170 470338 64226
rect 470406 64170 470462 64226
rect 470034 64046 470090 64102
rect 470158 64046 470214 64102
rect 470282 64046 470338 64102
rect 470406 64046 470462 64102
rect 470034 63922 470090 63978
rect 470158 63922 470214 63978
rect 470282 63922 470338 63978
rect 470406 63922 470462 63978
rect 470034 46294 470090 46350
rect 470158 46294 470214 46350
rect 470282 46294 470338 46350
rect 470406 46294 470462 46350
rect 470034 46170 470090 46226
rect 470158 46170 470214 46226
rect 470282 46170 470338 46226
rect 470406 46170 470462 46226
rect 470034 46046 470090 46102
rect 470158 46046 470214 46102
rect 470282 46046 470338 46102
rect 470406 46046 470462 46102
rect 470034 45922 470090 45978
rect 470158 45922 470214 45978
rect 470282 45922 470338 45978
rect 470406 45922 470462 45978
rect 497034 76294 497090 76350
rect 497158 76294 497214 76350
rect 497282 76294 497338 76350
rect 497406 76294 497462 76350
rect 497034 76170 497090 76226
rect 497158 76170 497214 76226
rect 497282 76170 497338 76226
rect 497406 76170 497462 76226
rect 497034 76046 497090 76102
rect 497158 76046 497214 76102
rect 497282 76046 497338 76102
rect 497406 76046 497462 76102
rect 497034 75922 497090 75978
rect 497158 75922 497214 75978
rect 497282 75922 497338 75978
rect 497406 75922 497462 75978
rect 495878 64294 495934 64350
rect 496002 64294 496058 64350
rect 495878 64170 495934 64226
rect 496002 64170 496058 64226
rect 495878 64046 495934 64102
rect 496002 64046 496058 64102
rect 495878 63922 495934 63978
rect 496002 63922 496058 63978
rect 480518 58294 480574 58350
rect 480642 58294 480698 58350
rect 480518 58170 480574 58226
rect 480642 58170 480698 58226
rect 480518 58046 480574 58102
rect 480642 58046 480698 58102
rect 480518 57922 480574 57978
rect 480642 57922 480698 57978
rect 497034 58294 497090 58350
rect 497158 58294 497214 58350
rect 497282 58294 497338 58350
rect 497406 58294 497462 58350
rect 497034 58170 497090 58226
rect 497158 58170 497214 58226
rect 497282 58170 497338 58226
rect 497406 58170 497462 58226
rect 497034 58046 497090 58102
rect 497158 58046 497214 58102
rect 497282 58046 497338 58102
rect 497406 58046 497462 58102
rect 497034 57922 497090 57978
rect 497158 57922 497214 57978
rect 497282 57922 497338 57978
rect 497406 57922 497462 57978
rect 473676 56222 473732 56278
rect 495878 46294 495934 46350
rect 496002 46294 496058 46350
rect 495878 46170 495934 46226
rect 496002 46170 496058 46226
rect 495878 46046 495934 46102
rect 496002 46046 496058 46102
rect 495878 45922 495934 45978
rect 496002 45922 496058 45978
rect 480518 40294 480574 40350
rect 480642 40294 480698 40350
rect 480518 40170 480574 40226
rect 480642 40170 480698 40226
rect 480518 40046 480574 40102
rect 480642 40046 480698 40102
rect 480518 39922 480574 39978
rect 480642 39922 480698 39978
rect 497034 40294 497090 40350
rect 497158 40294 497214 40350
rect 497282 40294 497338 40350
rect 497406 40294 497462 40350
rect 497034 40170 497090 40226
rect 497158 40170 497214 40226
rect 497282 40170 497338 40226
rect 497406 40170 497462 40226
rect 497034 40046 497090 40102
rect 497158 40046 497214 40102
rect 497282 40046 497338 40102
rect 497406 40046 497462 40102
rect 497034 39922 497090 39978
rect 497158 39922 497214 39978
rect 497282 39922 497338 39978
rect 497406 39922 497462 39978
rect 470034 28294 470090 28350
rect 470158 28294 470214 28350
rect 470282 28294 470338 28350
rect 470406 28294 470462 28350
rect 470034 28170 470090 28226
rect 470158 28170 470214 28226
rect 470282 28170 470338 28226
rect 470406 28170 470462 28226
rect 470034 28046 470090 28102
rect 470158 28046 470214 28102
rect 470282 28046 470338 28102
rect 470406 28046 470462 28102
rect 470034 27922 470090 27978
rect 470158 27922 470214 27978
rect 470282 27922 470338 27978
rect 470406 27922 470462 27978
rect 470034 10294 470090 10350
rect 470158 10294 470214 10350
rect 470282 10294 470338 10350
rect 470406 10294 470462 10350
rect 470034 10170 470090 10226
rect 470158 10170 470214 10226
rect 470282 10170 470338 10226
rect 470406 10170 470462 10226
rect 470034 10046 470090 10102
rect 470158 10046 470214 10102
rect 470282 10046 470338 10102
rect 470406 10046 470462 10102
rect 470034 9922 470090 9978
rect 470158 9922 470214 9978
rect 470282 9922 470338 9978
rect 470406 9922 470462 9978
rect 470034 -1176 470090 -1120
rect 470158 -1176 470214 -1120
rect 470282 -1176 470338 -1120
rect 470406 -1176 470462 -1120
rect 470034 -1300 470090 -1244
rect 470158 -1300 470214 -1244
rect 470282 -1300 470338 -1244
rect 470406 -1300 470462 -1244
rect 470034 -1424 470090 -1368
rect 470158 -1424 470214 -1368
rect 470282 -1424 470338 -1368
rect 470406 -1424 470462 -1368
rect 470034 -1548 470090 -1492
rect 470158 -1548 470214 -1492
rect 470282 -1548 470338 -1492
rect 470406 -1548 470462 -1492
rect 497034 22294 497090 22350
rect 497158 22294 497214 22350
rect 497282 22294 497338 22350
rect 497406 22294 497462 22350
rect 497034 22170 497090 22226
rect 497158 22170 497214 22226
rect 497282 22170 497338 22226
rect 497406 22170 497462 22226
rect 497034 22046 497090 22102
rect 497158 22046 497214 22102
rect 497282 22046 497338 22102
rect 497406 22046 497462 22102
rect 497034 21922 497090 21978
rect 497158 21922 497214 21978
rect 497282 21922 497338 21978
rect 497406 21922 497462 21978
rect 497034 4294 497090 4350
rect 497158 4294 497214 4350
rect 497282 4294 497338 4350
rect 497406 4294 497462 4350
rect 497034 4170 497090 4226
rect 497158 4170 497214 4226
rect 497282 4170 497338 4226
rect 497406 4170 497462 4226
rect 497034 4046 497090 4102
rect 497158 4046 497214 4102
rect 497282 4046 497338 4102
rect 497406 4046 497462 4102
rect 497034 3922 497090 3978
rect 497158 3922 497214 3978
rect 497282 3922 497338 3978
rect 497406 3922 497462 3978
rect 497034 -216 497090 -160
rect 497158 -216 497214 -160
rect 497282 -216 497338 -160
rect 497406 -216 497462 -160
rect 497034 -340 497090 -284
rect 497158 -340 497214 -284
rect 497282 -340 497338 -284
rect 497406 -340 497462 -284
rect 497034 -464 497090 -408
rect 497158 -464 497214 -408
rect 497282 -464 497338 -408
rect 497406 -464 497462 -408
rect 497034 -588 497090 -532
rect 497158 -588 497214 -532
rect 497282 -588 497338 -532
rect 497406 -588 497462 -532
rect 527754 166294 527810 166350
rect 527878 166294 527934 166350
rect 528002 166294 528058 166350
rect 528126 166294 528182 166350
rect 527754 166170 527810 166226
rect 527878 166170 527934 166226
rect 528002 166170 528058 166226
rect 528126 166170 528182 166226
rect 527754 166046 527810 166102
rect 527878 166046 527934 166102
rect 528002 166046 528058 166102
rect 528126 166046 528182 166102
rect 527754 165922 527810 165978
rect 527878 165922 527934 165978
rect 528002 165922 528058 165978
rect 528126 165922 528182 165978
rect 527754 148294 527810 148350
rect 527878 148294 527934 148350
rect 528002 148294 528058 148350
rect 528126 148294 528182 148350
rect 527754 148170 527810 148226
rect 527878 148170 527934 148226
rect 528002 148170 528058 148226
rect 528126 148170 528182 148226
rect 527754 148046 527810 148102
rect 527878 148046 527934 148102
rect 528002 148046 528058 148102
rect 528126 148046 528182 148102
rect 527754 147922 527810 147978
rect 527878 147922 527934 147978
rect 528002 147922 528058 147978
rect 528126 147922 528182 147978
rect 527754 130294 527810 130350
rect 527878 130294 527934 130350
rect 528002 130294 528058 130350
rect 528126 130294 528182 130350
rect 527754 130170 527810 130226
rect 527878 130170 527934 130226
rect 528002 130170 528058 130226
rect 528126 130170 528182 130226
rect 527754 130046 527810 130102
rect 527878 130046 527934 130102
rect 528002 130046 528058 130102
rect 528126 130046 528182 130102
rect 527754 129922 527810 129978
rect 527878 129922 527934 129978
rect 528002 129922 528058 129978
rect 528126 129922 528182 129978
rect 511238 112294 511294 112350
rect 511362 112294 511418 112350
rect 511238 112170 511294 112226
rect 511362 112170 511418 112226
rect 511238 112046 511294 112102
rect 511362 112046 511418 112102
rect 511238 111922 511294 111978
rect 511362 111922 511418 111978
rect 534268 402902 534324 402958
rect 557878 406294 557934 406350
rect 558002 406294 558058 406350
rect 557878 406170 557934 406226
rect 558002 406170 558058 406226
rect 557878 406046 557934 406102
rect 558002 406046 558058 406102
rect 557878 405922 557934 405978
rect 558002 405922 558058 405978
rect 542518 400294 542574 400350
rect 542642 400294 542698 400350
rect 542518 400170 542574 400226
rect 542642 400170 542698 400226
rect 542518 400046 542574 400102
rect 542642 400046 542698 400102
rect 542518 399922 542574 399978
rect 542642 399922 542698 399978
rect 558474 400294 558530 400350
rect 558598 400294 558654 400350
rect 558722 400294 558778 400350
rect 558846 400294 558902 400350
rect 558474 400170 558530 400226
rect 558598 400170 558654 400226
rect 558722 400170 558778 400226
rect 558846 400170 558902 400226
rect 558474 400046 558530 400102
rect 558598 400046 558654 400102
rect 558722 400046 558778 400102
rect 558846 400046 558902 400102
rect 558474 399922 558530 399978
rect 558598 399922 558654 399978
rect 558722 399922 558778 399978
rect 558846 399922 558902 399978
rect 557836 388333 557892 388389
rect 557940 388333 557996 388389
rect 558044 388333 558100 388389
rect 558474 382294 558530 382350
rect 558598 382294 558654 382350
rect 558722 382294 558778 382350
rect 558846 382294 558902 382350
rect 558474 382170 558530 382226
rect 558598 382170 558654 382226
rect 558722 382170 558778 382226
rect 558846 382170 558902 382226
rect 558474 382046 558530 382102
rect 558598 382046 558654 382102
rect 558722 382046 558778 382102
rect 558846 382046 558902 382102
rect 558474 381922 558530 381978
rect 558598 381922 558654 381978
rect 558722 381922 558778 381978
rect 558846 381922 558902 381978
rect 531474 370294 531530 370350
rect 531598 370294 531654 370350
rect 531722 370294 531778 370350
rect 531846 370294 531902 370350
rect 531474 370170 531530 370226
rect 531598 370170 531654 370226
rect 531722 370170 531778 370226
rect 531846 370170 531902 370226
rect 531474 370046 531530 370102
rect 531598 370046 531654 370102
rect 531722 370046 531778 370102
rect 531846 370046 531902 370102
rect 531474 369922 531530 369978
rect 531598 369922 531654 369978
rect 531722 369922 531778 369978
rect 531846 369922 531902 369978
rect 558474 364294 558530 364350
rect 558598 364294 558654 364350
rect 558722 364294 558778 364350
rect 558846 364294 558902 364350
rect 558474 364170 558530 364226
rect 558598 364170 558654 364226
rect 558722 364170 558778 364226
rect 558846 364170 558902 364226
rect 558474 364046 558530 364102
rect 558598 364046 558654 364102
rect 558722 364046 558778 364102
rect 558846 364046 558902 364102
rect 558474 363922 558530 363978
rect 558598 363922 558654 363978
rect 558722 363922 558778 363978
rect 558846 363922 558902 363978
rect 531474 352294 531530 352350
rect 531598 352294 531654 352350
rect 531722 352294 531778 352350
rect 531846 352294 531902 352350
rect 531474 352170 531530 352226
rect 531598 352170 531654 352226
rect 531722 352170 531778 352226
rect 531846 352170 531902 352226
rect 531474 352046 531530 352102
rect 531598 352046 531654 352102
rect 531722 352046 531778 352102
rect 531846 352046 531902 352102
rect 531474 351922 531530 351978
rect 531598 351922 531654 351978
rect 531722 351922 531778 351978
rect 531846 351922 531902 351978
rect 534268 341882 534324 341938
rect 531474 334294 531530 334350
rect 531598 334294 531654 334350
rect 531722 334294 531778 334350
rect 531846 334294 531902 334350
rect 557878 352294 557934 352350
rect 558002 352294 558058 352350
rect 557878 352170 557934 352226
rect 558002 352170 558058 352226
rect 557878 352046 557934 352102
rect 558002 352046 558058 352102
rect 557878 351922 557934 351978
rect 558002 351922 558058 351978
rect 542518 346294 542574 346350
rect 542642 346294 542698 346350
rect 542518 346170 542574 346226
rect 542642 346170 542698 346226
rect 542518 346046 542574 346102
rect 542642 346046 542698 346102
rect 542518 345922 542574 345978
rect 542642 345922 542698 345978
rect 558474 346294 558530 346350
rect 558598 346294 558654 346350
rect 558722 346294 558778 346350
rect 558846 346294 558902 346350
rect 558474 346170 558530 346226
rect 558598 346170 558654 346226
rect 558722 346170 558778 346226
rect 558846 346170 558902 346226
rect 558474 346046 558530 346102
rect 558598 346046 558654 346102
rect 558722 346046 558778 346102
rect 558846 346046 558902 346102
rect 558474 345922 558530 345978
rect 558598 345922 558654 345978
rect 558722 345922 558778 345978
rect 558846 345922 558902 345978
rect 557878 334294 557934 334350
rect 558002 334294 558058 334350
rect 531474 334170 531530 334226
rect 531598 334170 531654 334226
rect 531722 334170 531778 334226
rect 531846 334170 531902 334226
rect 531474 334046 531530 334102
rect 531598 334046 531654 334102
rect 531722 334046 531778 334102
rect 531846 334046 531902 334102
rect 531474 333922 531530 333978
rect 531598 333922 531654 333978
rect 531722 333922 531778 333978
rect 531846 333922 531902 333978
rect 557878 334170 557934 334226
rect 558002 334170 558058 334226
rect 557878 334046 557934 334102
rect 558002 334046 558058 334102
rect 557878 333922 557934 333978
rect 558002 333922 558058 333978
rect 534268 330002 534324 330058
rect 542518 328294 542574 328350
rect 542642 328294 542698 328350
rect 542518 328170 542574 328226
rect 542642 328170 542698 328226
rect 542518 328046 542574 328102
rect 542642 328046 542698 328102
rect 542518 327922 542574 327978
rect 542642 327922 542698 327978
rect 573238 472294 573294 472350
rect 573362 472294 573418 472350
rect 573238 472170 573294 472226
rect 573362 472170 573418 472226
rect 573238 472046 573294 472102
rect 573362 472046 573418 472102
rect 573238 471922 573294 471978
rect 573362 471922 573418 471978
rect 579292 469868 579348 469918
rect 579292 469862 579348 469868
rect 579404 468602 579460 468658
rect 579628 468602 579684 468658
rect 562194 460294 562250 460350
rect 562318 460294 562374 460350
rect 562442 460294 562498 460350
rect 562566 460294 562622 460350
rect 562194 460170 562250 460226
rect 562318 460170 562374 460226
rect 562442 460170 562498 460226
rect 562566 460170 562622 460226
rect 562194 460046 562250 460102
rect 562318 460046 562374 460102
rect 562442 460046 562498 460102
rect 562566 460046 562622 460102
rect 562194 459922 562250 459978
rect 562318 459922 562374 459978
rect 562442 459922 562498 459978
rect 562566 459922 562622 459978
rect 562194 442294 562250 442350
rect 562318 442294 562374 442350
rect 562442 442294 562498 442350
rect 562566 442294 562622 442350
rect 562194 442170 562250 442226
rect 562318 442170 562374 442226
rect 562442 442170 562498 442226
rect 562566 442170 562622 442226
rect 562194 442046 562250 442102
rect 562318 442046 562374 442102
rect 562442 442046 562498 442102
rect 562566 442046 562622 442102
rect 562194 441922 562250 441978
rect 562318 441922 562374 441978
rect 562442 441922 562498 441978
rect 562566 441922 562622 441978
rect 582988 470222 583044 470278
rect 562194 424294 562250 424350
rect 562318 424294 562374 424350
rect 562442 424294 562498 424350
rect 562566 424294 562622 424350
rect 562194 424170 562250 424226
rect 562318 424170 562374 424226
rect 562442 424170 562498 424226
rect 562566 424170 562622 424226
rect 562194 424046 562250 424102
rect 562318 424046 562374 424102
rect 562442 424046 562498 424102
rect 562566 424046 562622 424102
rect 562194 423922 562250 423978
rect 562318 423922 562374 423978
rect 562442 423922 562498 423978
rect 562566 423922 562622 423978
rect 573238 418294 573294 418350
rect 573362 418294 573418 418350
rect 573238 418170 573294 418226
rect 573362 418170 573418 418226
rect 573238 418046 573294 418102
rect 573362 418046 573418 418102
rect 573238 417922 573294 417978
rect 573362 417922 573418 417978
rect 579628 411722 579684 411778
rect 579292 410642 579348 410698
rect 579292 409388 579348 409438
rect 579292 409382 579348 409388
rect 579852 407042 579908 407098
rect 562194 406294 562250 406350
rect 562318 406294 562374 406350
rect 562442 406294 562498 406350
rect 562566 406294 562622 406350
rect 562194 406170 562250 406226
rect 562318 406170 562374 406226
rect 562442 406170 562498 406226
rect 562566 406170 562622 406226
rect 562194 406046 562250 406102
rect 562318 406046 562374 406102
rect 562442 406046 562498 406102
rect 562566 406046 562622 406102
rect 562194 405922 562250 405978
rect 562318 405922 562374 405978
rect 562442 405922 562498 405978
rect 562566 405922 562622 405978
rect 579740 403802 579796 403858
rect 579628 402556 579684 402598
rect 579628 402542 579684 402556
rect 573238 400294 573294 400350
rect 573362 400294 573418 400350
rect 573238 400170 573294 400226
rect 573362 400170 573418 400226
rect 573238 400046 573294 400102
rect 573362 400046 573418 400102
rect 573238 399922 573294 399978
rect 573362 399922 573418 399978
rect 579628 391076 579684 391078
rect 579628 391022 579684 391076
rect 562194 388294 562250 388350
rect 562318 388294 562374 388350
rect 562442 388294 562498 388350
rect 562566 388294 562622 388350
rect 562194 388170 562250 388226
rect 562318 388170 562374 388226
rect 562442 388170 562498 388226
rect 562566 388170 562622 388226
rect 562194 388046 562250 388102
rect 562318 388046 562374 388102
rect 562442 388046 562498 388102
rect 562566 388046 562622 388102
rect 562194 387922 562250 387978
rect 562318 387922 562374 387978
rect 562442 387922 562498 387978
rect 562566 387922 562622 387978
rect 562194 370294 562250 370350
rect 562318 370294 562374 370350
rect 562442 370294 562498 370350
rect 562566 370294 562622 370350
rect 562194 370170 562250 370226
rect 562318 370170 562374 370226
rect 562442 370170 562498 370226
rect 562566 370170 562622 370226
rect 562194 370046 562250 370102
rect 562318 370046 562374 370102
rect 562442 370046 562498 370102
rect 562566 370046 562622 370102
rect 562194 369922 562250 369978
rect 562318 369922 562374 369978
rect 562442 369922 562498 369978
rect 562566 369922 562622 369978
rect 562194 352294 562250 352350
rect 562318 352294 562374 352350
rect 562442 352294 562498 352350
rect 562566 352294 562622 352350
rect 562194 352170 562250 352226
rect 562318 352170 562374 352226
rect 562442 352170 562498 352226
rect 562566 352170 562622 352226
rect 562194 352046 562250 352102
rect 562318 352046 562374 352102
rect 562442 352046 562498 352102
rect 562566 352046 562622 352102
rect 562194 351922 562250 351978
rect 562318 351922 562374 351978
rect 562442 351922 562498 351978
rect 562566 351922 562622 351978
rect 573238 346294 573294 346350
rect 573362 346294 573418 346350
rect 573238 346170 573294 346226
rect 573362 346170 573418 346226
rect 573238 346046 573294 346102
rect 573362 346046 573418 346102
rect 573238 345922 573294 345978
rect 573362 345922 573418 345978
rect 558474 328294 558530 328350
rect 558598 328294 558654 328350
rect 558722 328294 558778 328350
rect 558846 328294 558902 328350
rect 558474 328170 558530 328226
rect 558598 328170 558654 328226
rect 558722 328170 558778 328226
rect 558846 328170 558902 328226
rect 558474 328046 558530 328102
rect 558598 328046 558654 328102
rect 558722 328046 558778 328102
rect 558846 328046 558902 328102
rect 558474 327922 558530 327978
rect 558598 327922 558654 327978
rect 558722 327922 558778 327978
rect 558846 327922 558902 327978
rect 535052 324962 535108 325018
rect 531474 316294 531530 316350
rect 531598 316294 531654 316350
rect 531722 316294 531778 316350
rect 531846 316294 531902 316350
rect 531474 316170 531530 316226
rect 531598 316170 531654 316226
rect 531722 316170 531778 316226
rect 531846 316170 531902 316226
rect 531474 316046 531530 316102
rect 531598 316046 531654 316102
rect 531722 316046 531778 316102
rect 531846 316046 531902 316102
rect 531474 315922 531530 315978
rect 531598 315922 531654 315978
rect 531722 315922 531778 315978
rect 531846 315922 531902 315978
rect 531474 298294 531530 298350
rect 531598 298294 531654 298350
rect 531722 298294 531778 298350
rect 531846 298294 531902 298350
rect 531474 298170 531530 298226
rect 531598 298170 531654 298226
rect 531722 298170 531778 298226
rect 531846 298170 531902 298226
rect 531474 298046 531530 298102
rect 531598 298046 531654 298102
rect 531722 298046 531778 298102
rect 531846 298046 531902 298102
rect 531474 297922 531530 297978
rect 531598 297922 531654 297978
rect 531722 297922 531778 297978
rect 531846 297922 531902 297978
rect 558474 310294 558530 310350
rect 558598 310294 558654 310350
rect 558722 310294 558778 310350
rect 558846 310294 558902 310350
rect 558474 310170 558530 310226
rect 558598 310170 558654 310226
rect 558722 310170 558778 310226
rect 558846 310170 558902 310226
rect 558474 310046 558530 310102
rect 558598 310046 558654 310102
rect 558722 310046 558778 310102
rect 558846 310046 558902 310102
rect 558474 309922 558530 309978
rect 558598 309922 558654 309978
rect 558722 309922 558778 309978
rect 558846 309922 558902 309978
rect 558474 292294 558530 292350
rect 558598 292294 558654 292350
rect 558722 292294 558778 292350
rect 558846 292294 558902 292350
rect 558474 292170 558530 292226
rect 558598 292170 558654 292226
rect 558722 292170 558778 292226
rect 558846 292170 558902 292226
rect 558474 292046 558530 292102
rect 558598 292046 558654 292102
rect 558722 292046 558778 292102
rect 558846 292046 558902 292102
rect 558474 291922 558530 291978
rect 558598 291922 558654 291978
rect 558722 291922 558778 291978
rect 558846 291922 558902 291978
rect 531474 280294 531530 280350
rect 531598 280294 531654 280350
rect 531722 280294 531778 280350
rect 531846 280294 531902 280350
rect 531474 280170 531530 280226
rect 531598 280170 531654 280226
rect 531722 280170 531778 280226
rect 531846 280170 531902 280226
rect 531474 280046 531530 280102
rect 531598 280046 531654 280102
rect 531722 280046 531778 280102
rect 531846 280046 531902 280102
rect 531474 279922 531530 279978
rect 531598 279922 531654 279978
rect 531722 279922 531778 279978
rect 531846 279922 531902 279978
rect 534268 269522 534324 269578
rect 534268 267902 534324 267958
rect 531474 262294 531530 262350
rect 531598 262294 531654 262350
rect 531722 262294 531778 262350
rect 531846 262294 531902 262350
rect 531474 262170 531530 262226
rect 531598 262170 531654 262226
rect 531722 262170 531778 262226
rect 531846 262170 531902 262226
rect 531474 262046 531530 262102
rect 531598 262046 531654 262102
rect 531722 262046 531778 262102
rect 531846 262046 531902 262102
rect 531474 261922 531530 261978
rect 531598 261922 531654 261978
rect 531722 261922 531778 261978
rect 531846 261922 531902 261978
rect 534268 260162 534324 260218
rect 557878 280294 557934 280350
rect 558002 280294 558058 280350
rect 557878 280170 557934 280226
rect 558002 280170 558058 280226
rect 557878 280046 557934 280102
rect 558002 280046 558058 280102
rect 557878 279922 557934 279978
rect 558002 279922 558058 279978
rect 542518 274294 542574 274350
rect 542642 274294 542698 274350
rect 542518 274170 542574 274226
rect 542642 274170 542698 274226
rect 542518 274046 542574 274102
rect 542642 274046 542698 274102
rect 542518 273922 542574 273978
rect 542642 273922 542698 273978
rect 558474 274294 558530 274350
rect 558598 274294 558654 274350
rect 558722 274294 558778 274350
rect 558846 274294 558902 274350
rect 558474 274170 558530 274226
rect 558598 274170 558654 274226
rect 558722 274170 558778 274226
rect 558846 274170 558902 274226
rect 558474 274046 558530 274102
rect 558598 274046 558654 274102
rect 558722 274046 558778 274102
rect 558846 274046 558902 274102
rect 558474 273922 558530 273978
rect 558598 273922 558654 273978
rect 558722 273922 558778 273978
rect 558846 273922 558902 273978
rect 557878 262294 557934 262350
rect 558002 262294 558058 262350
rect 557878 262170 557934 262226
rect 558002 262170 558058 262226
rect 557878 262046 557934 262102
rect 558002 262046 558058 262102
rect 557878 261922 557934 261978
rect 558002 261922 558058 261978
rect 542518 256294 542574 256350
rect 542642 256294 542698 256350
rect 542518 256170 542574 256226
rect 542642 256170 542698 256226
rect 542518 256046 542574 256102
rect 542642 256046 542698 256102
rect 542518 255922 542574 255978
rect 542642 255922 542698 255978
rect 558474 256294 558530 256350
rect 558598 256294 558654 256350
rect 558722 256294 558778 256350
rect 558846 256294 558902 256350
rect 558474 256170 558530 256226
rect 558598 256170 558654 256226
rect 558722 256170 558778 256226
rect 558846 256170 558902 256226
rect 558474 256046 558530 256102
rect 558598 256046 558654 256102
rect 558722 256046 558778 256102
rect 558846 256046 558902 256102
rect 558474 255922 558530 255978
rect 558598 255922 558654 255978
rect 558722 255922 558778 255978
rect 558846 255922 558902 255978
rect 531474 244294 531530 244350
rect 531598 244294 531654 244350
rect 531722 244294 531778 244350
rect 531846 244294 531902 244350
rect 531474 244170 531530 244226
rect 531598 244170 531654 244226
rect 531722 244170 531778 244226
rect 531846 244170 531902 244226
rect 531474 244046 531530 244102
rect 531598 244046 531654 244102
rect 531722 244046 531778 244102
rect 531846 244046 531902 244102
rect 531474 243922 531530 243978
rect 531598 243922 531654 243978
rect 531722 243922 531778 243978
rect 531846 243922 531902 243978
rect 531474 226294 531530 226350
rect 531598 226294 531654 226350
rect 531722 226294 531778 226350
rect 531846 226294 531902 226350
rect 531474 226170 531530 226226
rect 531598 226170 531654 226226
rect 531722 226170 531778 226226
rect 531846 226170 531902 226226
rect 531474 226046 531530 226102
rect 531598 226046 531654 226102
rect 531722 226046 531778 226102
rect 531846 226046 531902 226102
rect 531474 225922 531530 225978
rect 531598 225922 531654 225978
rect 531722 225922 531778 225978
rect 531846 225922 531902 225978
rect 558474 238294 558530 238350
rect 558598 238294 558654 238350
rect 558722 238294 558778 238350
rect 558846 238294 558902 238350
rect 558474 238170 558530 238226
rect 558598 238170 558654 238226
rect 558722 238170 558778 238226
rect 558846 238170 558902 238226
rect 558474 238046 558530 238102
rect 558598 238046 558654 238102
rect 558722 238046 558778 238102
rect 558846 238046 558902 238102
rect 558474 237922 558530 237978
rect 558598 237922 558654 237978
rect 558722 237922 558778 237978
rect 558846 237922 558902 237978
rect 558474 220294 558530 220350
rect 558598 220294 558654 220350
rect 558722 220294 558778 220350
rect 558846 220294 558902 220350
rect 558474 220170 558530 220226
rect 558598 220170 558654 220226
rect 558722 220170 558778 220226
rect 558846 220170 558902 220226
rect 558474 220046 558530 220102
rect 558598 220046 558654 220102
rect 558722 220046 558778 220102
rect 558846 220046 558902 220102
rect 558474 219922 558530 219978
rect 558598 219922 558654 219978
rect 558722 219922 558778 219978
rect 558846 219922 558902 219978
rect 531474 208294 531530 208350
rect 531598 208294 531654 208350
rect 531722 208294 531778 208350
rect 531846 208294 531902 208350
rect 531474 208170 531530 208226
rect 531598 208170 531654 208226
rect 531722 208170 531778 208226
rect 531846 208170 531902 208226
rect 531474 208046 531530 208102
rect 531598 208046 531654 208102
rect 531722 208046 531778 208102
rect 531846 208046 531902 208102
rect 531474 207922 531530 207978
rect 531598 207922 531654 207978
rect 531722 207922 531778 207978
rect 531846 207922 531902 207978
rect 534268 198242 534324 198298
rect 557878 208294 557934 208350
rect 558002 208294 558058 208350
rect 557878 208170 557934 208226
rect 558002 208170 558058 208226
rect 557878 208046 557934 208102
rect 558002 208046 558058 208102
rect 557878 207922 557934 207978
rect 558002 207922 558058 207978
rect 542518 202294 542574 202350
rect 542642 202294 542698 202350
rect 542518 202170 542574 202226
rect 542642 202170 542698 202226
rect 542518 202046 542574 202102
rect 542642 202046 542698 202102
rect 542518 201922 542574 201978
rect 542642 201922 542698 201978
rect 558474 202294 558530 202350
rect 558598 202294 558654 202350
rect 558722 202294 558778 202350
rect 558846 202294 558902 202350
rect 558474 202170 558530 202226
rect 558598 202170 558654 202226
rect 558722 202170 558778 202226
rect 558846 202170 558902 202226
rect 558474 202046 558530 202102
rect 558598 202046 558654 202102
rect 558722 202046 558778 202102
rect 558846 202046 558902 202102
rect 558474 201922 558530 201978
rect 558598 201922 558654 201978
rect 558722 201922 558778 201978
rect 558846 201922 558902 201978
rect 531474 190294 531530 190350
rect 531598 190294 531654 190350
rect 531722 190294 531778 190350
rect 531846 190294 531902 190350
rect 531474 190170 531530 190226
rect 531598 190170 531654 190226
rect 531722 190170 531778 190226
rect 531846 190170 531902 190226
rect 531474 190046 531530 190102
rect 531598 190046 531654 190102
rect 531722 190046 531778 190102
rect 531846 190046 531902 190102
rect 531474 189922 531530 189978
rect 531598 189922 531654 189978
rect 531722 189922 531778 189978
rect 531846 189922 531902 189978
rect 557878 190294 557934 190350
rect 558002 190294 558058 190350
rect 557878 190170 557934 190226
rect 558002 190170 558058 190226
rect 557878 190046 557934 190102
rect 558002 190046 558058 190102
rect 557878 189922 557934 189978
rect 558002 189922 558058 189978
rect 542518 184294 542574 184350
rect 542642 184294 542698 184350
rect 542518 184170 542574 184226
rect 542642 184170 542698 184226
rect 542518 184046 542574 184102
rect 542642 184046 542698 184102
rect 542518 183922 542574 183978
rect 542642 183922 542698 183978
rect 558474 184294 558530 184350
rect 558598 184294 558654 184350
rect 558722 184294 558778 184350
rect 558846 184294 558902 184350
rect 558474 184170 558530 184226
rect 558598 184170 558654 184226
rect 558722 184170 558778 184226
rect 558846 184170 558902 184226
rect 558474 184046 558530 184102
rect 558598 184046 558654 184102
rect 558722 184046 558778 184102
rect 558846 184046 558902 184102
rect 558474 183922 558530 183978
rect 558598 183922 558654 183978
rect 558722 183922 558778 183978
rect 558846 183922 558902 183978
rect 531474 172294 531530 172350
rect 531598 172294 531654 172350
rect 531722 172294 531778 172350
rect 531846 172294 531902 172350
rect 531474 172170 531530 172226
rect 531598 172170 531654 172226
rect 531722 172170 531778 172226
rect 531846 172170 531902 172226
rect 531474 172046 531530 172102
rect 531598 172046 531654 172102
rect 531722 172046 531778 172102
rect 531846 172046 531902 172102
rect 531474 171922 531530 171978
rect 531598 171922 531654 171978
rect 531722 171922 531778 171978
rect 531846 171922 531902 171978
rect 558474 166294 558530 166350
rect 558598 166294 558654 166350
rect 558722 166294 558778 166350
rect 558846 166294 558902 166350
rect 558474 166170 558530 166226
rect 558598 166170 558654 166226
rect 558722 166170 558778 166226
rect 558846 166170 558902 166226
rect 558474 166046 558530 166102
rect 558598 166046 558654 166102
rect 558722 166046 558778 166102
rect 558846 166046 558902 166102
rect 558474 165922 558530 165978
rect 558598 165922 558654 165978
rect 558722 165922 558778 165978
rect 558846 165922 558902 165978
rect 531474 154294 531530 154350
rect 531598 154294 531654 154350
rect 531722 154294 531778 154350
rect 531846 154294 531902 154350
rect 531474 154170 531530 154226
rect 531598 154170 531654 154226
rect 531722 154170 531778 154226
rect 531846 154170 531902 154226
rect 531474 154046 531530 154102
rect 531598 154046 531654 154102
rect 531722 154046 531778 154102
rect 531846 154046 531902 154102
rect 531474 153922 531530 153978
rect 531598 153922 531654 153978
rect 531722 153922 531778 153978
rect 531846 153922 531902 153978
rect 531474 136294 531530 136350
rect 531598 136294 531654 136350
rect 531722 136294 531778 136350
rect 531846 136294 531902 136350
rect 531474 136170 531530 136226
rect 531598 136170 531654 136226
rect 531722 136170 531778 136226
rect 531846 136170 531902 136226
rect 531474 136046 531530 136102
rect 531598 136046 531654 136102
rect 531722 136046 531778 136102
rect 531846 136046 531902 136102
rect 531474 135922 531530 135978
rect 531598 135922 531654 135978
rect 531722 135922 531778 135978
rect 531846 135922 531902 135978
rect 530796 127682 530852 127738
rect 527754 112294 527810 112350
rect 527878 112294 527934 112350
rect 528002 112294 528058 112350
rect 528126 112294 528182 112350
rect 527754 112170 527810 112226
rect 527878 112170 527934 112226
rect 528002 112170 528058 112226
rect 528126 112170 528182 112226
rect 527754 112046 527810 112102
rect 527878 112046 527934 112102
rect 528002 112046 528058 112102
rect 528126 112046 528182 112102
rect 527754 111922 527810 111978
rect 527878 111922 527934 111978
rect 528002 111922 528058 111978
rect 528126 111922 528182 111978
rect 500754 100294 500810 100350
rect 500878 100294 500934 100350
rect 501002 100294 501058 100350
rect 501126 100294 501182 100350
rect 500754 100170 500810 100226
rect 500878 100170 500934 100226
rect 501002 100170 501058 100226
rect 501126 100170 501182 100226
rect 500754 100046 500810 100102
rect 500878 100046 500934 100102
rect 501002 100046 501058 100102
rect 501126 100046 501182 100102
rect 500754 99922 500810 99978
rect 500878 99922 500934 99978
rect 501002 99922 501058 99978
rect 501126 99922 501182 99978
rect 500754 82294 500810 82350
rect 500878 82294 500934 82350
rect 501002 82294 501058 82350
rect 501126 82294 501182 82350
rect 500754 82170 500810 82226
rect 500878 82170 500934 82226
rect 501002 82170 501058 82226
rect 501126 82170 501182 82226
rect 500754 82046 500810 82102
rect 500878 82046 500934 82102
rect 501002 82046 501058 82102
rect 501126 82046 501182 82102
rect 500754 81922 500810 81978
rect 500878 81922 500934 81978
rect 501002 81922 501058 81978
rect 501126 81922 501182 81978
rect 500754 64294 500810 64350
rect 500878 64294 500934 64350
rect 501002 64294 501058 64350
rect 501126 64294 501182 64350
rect 500754 64170 500810 64226
rect 500878 64170 500934 64226
rect 501002 64170 501058 64226
rect 501126 64170 501182 64226
rect 500754 64046 500810 64102
rect 500878 64046 500934 64102
rect 501002 64046 501058 64102
rect 501126 64046 501182 64102
rect 500754 63922 500810 63978
rect 500878 63922 500934 63978
rect 501002 63922 501058 63978
rect 501126 63922 501182 63978
rect 511238 58294 511294 58350
rect 511362 58294 511418 58350
rect 511238 58170 511294 58226
rect 511362 58170 511418 58226
rect 511238 58046 511294 58102
rect 511362 58046 511418 58102
rect 511238 57922 511294 57978
rect 511362 57922 511418 57978
rect 500754 46294 500810 46350
rect 500878 46294 500934 46350
rect 501002 46294 501058 46350
rect 501126 46294 501182 46350
rect 500754 46170 500810 46226
rect 500878 46170 500934 46226
rect 501002 46170 501058 46226
rect 501126 46170 501182 46226
rect 500754 46046 500810 46102
rect 500878 46046 500934 46102
rect 501002 46046 501058 46102
rect 501126 46046 501182 46102
rect 500754 45922 500810 45978
rect 500878 45922 500934 45978
rect 501002 45922 501058 45978
rect 501126 45922 501182 45978
rect 531474 118294 531530 118350
rect 531598 118294 531654 118350
rect 531722 118294 531778 118350
rect 531846 118294 531902 118350
rect 531474 118170 531530 118226
rect 531598 118170 531654 118226
rect 531722 118170 531778 118226
rect 531846 118170 531902 118226
rect 531474 118046 531530 118102
rect 531598 118046 531654 118102
rect 531722 118046 531778 118102
rect 531846 118046 531902 118102
rect 531474 117922 531530 117978
rect 531598 117922 531654 117978
rect 531722 117922 531778 117978
rect 531846 117922 531902 117978
rect 527754 94294 527810 94350
rect 527878 94294 527934 94350
rect 528002 94294 528058 94350
rect 528126 94294 528182 94350
rect 527754 94170 527810 94226
rect 527878 94170 527934 94226
rect 528002 94170 528058 94226
rect 528126 94170 528182 94226
rect 527754 94046 527810 94102
rect 527878 94046 527934 94102
rect 528002 94046 528058 94102
rect 528126 94046 528182 94102
rect 527754 93922 527810 93978
rect 527878 93922 527934 93978
rect 528002 93922 528058 93978
rect 528126 93922 528182 93978
rect 527754 76294 527810 76350
rect 527878 76294 527934 76350
rect 528002 76294 528058 76350
rect 528126 76294 528182 76350
rect 527754 76170 527810 76226
rect 527878 76170 527934 76226
rect 528002 76170 528058 76226
rect 528126 76170 528182 76226
rect 527754 76046 527810 76102
rect 527878 76046 527934 76102
rect 528002 76046 528058 76102
rect 528126 76046 528182 76102
rect 527754 75922 527810 75978
rect 527878 75922 527934 75978
rect 528002 75922 528058 75978
rect 528126 75922 528182 75978
rect 527754 58294 527810 58350
rect 527878 58294 527934 58350
rect 528002 58294 528058 58350
rect 528126 58294 528182 58350
rect 527754 58170 527810 58226
rect 527878 58170 527934 58226
rect 528002 58170 528058 58226
rect 528126 58170 528182 58226
rect 527754 58046 527810 58102
rect 527878 58046 527934 58102
rect 528002 58046 528058 58102
rect 528126 58046 528182 58102
rect 527754 57922 527810 57978
rect 527878 57922 527934 57978
rect 528002 57922 528058 57978
rect 528126 57922 528182 57978
rect 511238 40294 511294 40350
rect 511362 40294 511418 40350
rect 511238 40170 511294 40226
rect 511362 40170 511418 40226
rect 511238 40046 511294 40102
rect 511362 40046 511418 40102
rect 511238 39922 511294 39978
rect 511362 39922 511418 39978
rect 558474 148294 558530 148350
rect 558598 148294 558654 148350
rect 558722 148294 558778 148350
rect 558846 148294 558902 148350
rect 558474 148170 558530 148226
rect 558598 148170 558654 148226
rect 558722 148170 558778 148226
rect 558846 148170 558902 148226
rect 558474 148046 558530 148102
rect 558598 148046 558654 148102
rect 558722 148046 558778 148102
rect 558846 148046 558902 148102
rect 558474 147922 558530 147978
rect 558598 147922 558654 147978
rect 558722 147922 558778 147978
rect 558846 147922 558902 147978
rect 557878 136294 557934 136350
rect 558002 136294 558058 136350
rect 557878 136170 557934 136226
rect 558002 136170 558058 136226
rect 557878 136046 557934 136102
rect 558002 136046 558058 136102
rect 557878 135922 557934 135978
rect 558002 135922 558058 135978
rect 542518 130294 542574 130350
rect 542642 130294 542698 130350
rect 542518 130170 542574 130226
rect 542642 130170 542698 130226
rect 542518 130046 542574 130102
rect 542642 130046 542698 130102
rect 542518 129922 542574 129978
rect 542642 129922 542698 129978
rect 558474 130294 558530 130350
rect 558598 130294 558654 130350
rect 558722 130294 558778 130350
rect 558846 130294 558902 130350
rect 558474 130170 558530 130226
rect 558598 130170 558654 130226
rect 558722 130170 558778 130226
rect 558846 130170 558902 130226
rect 558474 130046 558530 130102
rect 558598 130046 558654 130102
rect 558722 130046 558778 130102
rect 558846 130046 558902 130102
rect 558474 129922 558530 129978
rect 558598 129922 558654 129978
rect 558722 129922 558778 129978
rect 558846 129922 558902 129978
rect 557878 118294 557934 118350
rect 558002 118294 558058 118350
rect 557878 118170 557934 118226
rect 558002 118170 558058 118226
rect 557878 118046 557934 118102
rect 558002 118046 558058 118102
rect 557878 117922 557934 117978
rect 558002 117922 558058 117978
rect 542518 112294 542574 112350
rect 542642 112294 542698 112350
rect 542518 112170 542574 112226
rect 542642 112170 542698 112226
rect 542518 112046 542574 112102
rect 542642 112046 542698 112102
rect 542518 111922 542574 111978
rect 542642 111922 542698 111978
rect 558474 112294 558530 112350
rect 558598 112294 558654 112350
rect 558722 112294 558778 112350
rect 558846 112294 558902 112350
rect 558474 112170 558530 112226
rect 558598 112170 558654 112226
rect 558722 112170 558778 112226
rect 558846 112170 558902 112226
rect 558474 112046 558530 112102
rect 558598 112046 558654 112102
rect 558722 112046 558778 112102
rect 558846 112046 558902 112102
rect 558474 111922 558530 111978
rect 558598 111922 558654 111978
rect 558722 111922 558778 111978
rect 558846 111922 558902 111978
rect 531474 100294 531530 100350
rect 531598 100294 531654 100350
rect 531722 100294 531778 100350
rect 531846 100294 531902 100350
rect 531474 100170 531530 100226
rect 531598 100170 531654 100226
rect 531722 100170 531778 100226
rect 531846 100170 531902 100226
rect 531474 100046 531530 100102
rect 531598 100046 531654 100102
rect 531722 100046 531778 100102
rect 531846 100046 531902 100102
rect 531474 99922 531530 99978
rect 531598 99922 531654 99978
rect 531722 99922 531778 99978
rect 531846 99922 531902 99978
rect 531474 82294 531530 82350
rect 531598 82294 531654 82350
rect 531722 82294 531778 82350
rect 531846 82294 531902 82350
rect 531474 82170 531530 82226
rect 531598 82170 531654 82226
rect 531722 82170 531778 82226
rect 531846 82170 531902 82226
rect 531474 82046 531530 82102
rect 531598 82046 531654 82102
rect 531722 82046 531778 82102
rect 531846 82046 531902 82102
rect 531474 81922 531530 81978
rect 531598 81922 531654 81978
rect 531722 81922 531778 81978
rect 531846 81922 531902 81978
rect 531474 64294 531530 64350
rect 531598 64294 531654 64350
rect 531722 64294 531778 64350
rect 531846 64294 531902 64350
rect 531474 64170 531530 64226
rect 531598 64170 531654 64226
rect 531722 64170 531778 64226
rect 531846 64170 531902 64226
rect 531474 64046 531530 64102
rect 531598 64046 531654 64102
rect 531722 64046 531778 64102
rect 531846 64046 531902 64102
rect 531474 63922 531530 63978
rect 531598 63922 531654 63978
rect 531722 63922 531778 63978
rect 531846 63922 531902 63978
rect 527754 40294 527810 40350
rect 527878 40294 527934 40350
rect 528002 40294 528058 40350
rect 528126 40294 528182 40350
rect 527754 40170 527810 40226
rect 527878 40170 527934 40226
rect 528002 40170 528058 40226
rect 528126 40170 528182 40226
rect 527754 40046 527810 40102
rect 527878 40046 527934 40102
rect 528002 40046 528058 40102
rect 528126 40046 528182 40102
rect 527754 39922 527810 39978
rect 527878 39922 527934 39978
rect 528002 39922 528058 39978
rect 528126 39922 528182 39978
rect 500754 28294 500810 28350
rect 500878 28294 500934 28350
rect 501002 28294 501058 28350
rect 501126 28294 501182 28350
rect 500754 28170 500810 28226
rect 500878 28170 500934 28226
rect 501002 28170 501058 28226
rect 501126 28170 501182 28226
rect 500754 28046 500810 28102
rect 500878 28046 500934 28102
rect 501002 28046 501058 28102
rect 501126 28046 501182 28102
rect 500754 27922 500810 27978
rect 500878 27922 500934 27978
rect 501002 27922 501058 27978
rect 501126 27922 501182 27978
rect 500754 10294 500810 10350
rect 500878 10294 500934 10350
rect 501002 10294 501058 10350
rect 501126 10294 501182 10350
rect 500754 10170 500810 10226
rect 500878 10170 500934 10226
rect 501002 10170 501058 10226
rect 501126 10170 501182 10226
rect 500754 10046 500810 10102
rect 500878 10046 500934 10102
rect 501002 10046 501058 10102
rect 501126 10046 501182 10102
rect 500754 9922 500810 9978
rect 500878 9922 500934 9978
rect 501002 9922 501058 9978
rect 501126 9922 501182 9978
rect 500754 -1176 500810 -1120
rect 500878 -1176 500934 -1120
rect 501002 -1176 501058 -1120
rect 501126 -1176 501182 -1120
rect 500754 -1300 500810 -1244
rect 500878 -1300 500934 -1244
rect 501002 -1300 501058 -1244
rect 501126 -1300 501182 -1244
rect 500754 -1424 500810 -1368
rect 500878 -1424 500934 -1368
rect 501002 -1424 501058 -1368
rect 501126 -1424 501182 -1368
rect 500754 -1548 500810 -1492
rect 500878 -1548 500934 -1492
rect 501002 -1548 501058 -1492
rect 501126 -1548 501182 -1492
rect 527754 22294 527810 22350
rect 527878 22294 527934 22350
rect 528002 22294 528058 22350
rect 528126 22294 528182 22350
rect 527754 22170 527810 22226
rect 527878 22170 527934 22226
rect 528002 22170 528058 22226
rect 528126 22170 528182 22226
rect 527754 22046 527810 22102
rect 527878 22046 527934 22102
rect 528002 22046 528058 22102
rect 528126 22046 528182 22102
rect 527754 21922 527810 21978
rect 527878 21922 527934 21978
rect 528002 21922 528058 21978
rect 528126 21922 528182 21978
rect 527754 4294 527810 4350
rect 527878 4294 527934 4350
rect 528002 4294 528058 4350
rect 528126 4294 528182 4350
rect 527754 4170 527810 4226
rect 527878 4170 527934 4226
rect 528002 4170 528058 4226
rect 528126 4170 528182 4226
rect 527754 4046 527810 4102
rect 527878 4046 527934 4102
rect 528002 4046 528058 4102
rect 528126 4046 528182 4102
rect 527754 3922 527810 3978
rect 527878 3922 527934 3978
rect 528002 3922 528058 3978
rect 528126 3922 528182 3978
rect 527754 -216 527810 -160
rect 527878 -216 527934 -160
rect 528002 -216 528058 -160
rect 528126 -216 528182 -160
rect 527754 -340 527810 -284
rect 527878 -340 527934 -284
rect 528002 -340 528058 -284
rect 528126 -340 528182 -284
rect 527754 -464 527810 -408
rect 527878 -464 527934 -408
rect 528002 -464 528058 -408
rect 528126 -464 528182 -408
rect 527754 -588 527810 -532
rect 527878 -588 527934 -532
rect 528002 -588 528058 -532
rect 528126 -588 528182 -532
rect 534268 56222 534324 56278
rect 558474 94294 558530 94350
rect 558598 94294 558654 94350
rect 558722 94294 558778 94350
rect 558846 94294 558902 94350
rect 558474 94170 558530 94226
rect 558598 94170 558654 94226
rect 558722 94170 558778 94226
rect 558846 94170 558902 94226
rect 558474 94046 558530 94102
rect 558598 94046 558654 94102
rect 558722 94046 558778 94102
rect 558846 94046 558902 94102
rect 558474 93922 558530 93978
rect 558598 93922 558654 93978
rect 558722 93922 558778 93978
rect 558846 93922 558902 93978
rect 531474 46294 531530 46350
rect 531598 46294 531654 46350
rect 531722 46294 531778 46350
rect 531846 46294 531902 46350
rect 531474 46170 531530 46226
rect 531598 46170 531654 46226
rect 531722 46170 531778 46226
rect 531846 46170 531902 46226
rect 531474 46046 531530 46102
rect 531598 46046 531654 46102
rect 531722 46046 531778 46102
rect 531846 46046 531902 46102
rect 558474 76294 558530 76350
rect 558598 76294 558654 76350
rect 558722 76294 558778 76350
rect 558846 76294 558902 76350
rect 558474 76170 558530 76226
rect 558598 76170 558654 76226
rect 558722 76170 558778 76226
rect 558846 76170 558902 76226
rect 558474 76046 558530 76102
rect 558598 76046 558654 76102
rect 558722 76046 558778 76102
rect 558846 76046 558902 76102
rect 558474 75922 558530 75978
rect 558598 75922 558654 75978
rect 558722 75922 558778 75978
rect 558846 75922 558902 75978
rect 531474 45922 531530 45978
rect 531598 45922 531654 45978
rect 531722 45922 531778 45978
rect 531846 45922 531902 45978
rect 557878 64294 557934 64350
rect 558002 64294 558058 64350
rect 557878 64170 557934 64226
rect 558002 64170 558058 64226
rect 557878 64046 557934 64102
rect 558002 64046 558058 64102
rect 557878 63922 557934 63978
rect 558002 63922 558058 63978
rect 542518 58294 542574 58350
rect 542642 58294 542698 58350
rect 542518 58170 542574 58226
rect 542642 58170 542698 58226
rect 542518 58046 542574 58102
rect 542642 58046 542698 58102
rect 542518 57922 542574 57978
rect 542642 57922 542698 57978
rect 558474 58294 558530 58350
rect 558598 58294 558654 58350
rect 558722 58294 558778 58350
rect 558846 58294 558902 58350
rect 558474 58170 558530 58226
rect 558598 58170 558654 58226
rect 558722 58170 558778 58226
rect 558846 58170 558902 58226
rect 558474 58046 558530 58102
rect 558598 58046 558654 58102
rect 558722 58046 558778 58102
rect 558846 58046 558902 58102
rect 558474 57922 558530 57978
rect 558598 57922 558654 57978
rect 558722 57922 558778 57978
rect 558846 57922 558902 57978
rect 579628 331660 579684 331678
rect 579628 331622 579684 331660
rect 573238 328294 573294 328350
rect 573362 328294 573418 328350
rect 573238 328170 573294 328226
rect 573362 328170 573418 328226
rect 573238 328046 573294 328102
rect 573362 328046 573418 328102
rect 573238 327922 573294 327978
rect 573362 327922 573418 327978
rect 582988 326762 583044 326818
rect 562194 316294 562250 316350
rect 562318 316294 562374 316350
rect 562442 316294 562498 316350
rect 562566 316294 562622 316350
rect 562194 316170 562250 316226
rect 562318 316170 562374 316226
rect 562442 316170 562498 316226
rect 562566 316170 562622 316226
rect 562194 316046 562250 316102
rect 562318 316046 562374 316102
rect 562442 316046 562498 316102
rect 562566 316046 562622 316102
rect 562194 315922 562250 315978
rect 562318 315922 562374 315978
rect 562442 315922 562498 315978
rect 562566 315922 562622 315978
rect 562940 313982 562996 314038
rect 562194 298294 562250 298350
rect 562318 298294 562374 298350
rect 562442 298294 562498 298350
rect 562566 298294 562622 298350
rect 562194 298170 562250 298226
rect 562318 298170 562374 298226
rect 562442 298170 562498 298226
rect 562566 298170 562622 298226
rect 562194 298046 562250 298102
rect 562318 298046 562374 298102
rect 562442 298046 562498 298102
rect 562566 298046 562622 298102
rect 562194 297922 562250 297978
rect 562318 297922 562374 297978
rect 562442 297922 562498 297978
rect 562566 297922 562622 297978
rect 562194 280294 562250 280350
rect 562318 280294 562374 280350
rect 562442 280294 562498 280350
rect 562566 280294 562622 280350
rect 562194 280170 562250 280226
rect 562318 280170 562374 280226
rect 562442 280170 562498 280226
rect 562566 280170 562622 280226
rect 562194 280046 562250 280102
rect 562318 280046 562374 280102
rect 562442 280046 562498 280102
rect 562566 280046 562622 280102
rect 562194 279922 562250 279978
rect 562318 279922 562374 279978
rect 562442 279922 562498 279978
rect 562566 279922 562622 279978
rect 573238 274294 573294 274350
rect 573362 274294 573418 274350
rect 573238 274170 573294 274226
rect 573362 274170 573418 274226
rect 573238 274046 573294 274102
rect 573362 274046 573418 274102
rect 573238 273922 573294 273978
rect 573362 273922 573418 273978
rect 579292 267036 579348 267058
rect 579292 267002 579348 267036
rect 579068 266642 579124 266698
rect 562194 262294 562250 262350
rect 562318 262294 562374 262350
rect 562442 262294 562498 262350
rect 562566 262294 562622 262350
rect 562194 262170 562250 262226
rect 562318 262170 562374 262226
rect 562442 262170 562498 262226
rect 562566 262170 562622 262226
rect 562194 262046 562250 262102
rect 562318 262046 562374 262102
rect 562442 262046 562498 262102
rect 562566 262046 562622 262102
rect 562194 261922 562250 261978
rect 562318 261922 562374 261978
rect 562442 261922 562498 261978
rect 562566 261922 562622 261978
rect 579292 260882 579348 260938
rect 579628 260342 579684 260398
rect 582988 268802 583044 268858
rect 573238 256294 573294 256350
rect 573362 256294 573418 256350
rect 573238 256170 573294 256226
rect 573362 256170 573418 256226
rect 573238 256046 573294 256102
rect 573362 256046 573418 256102
rect 573238 255922 573294 255978
rect 573362 255922 573418 255978
rect 562194 244294 562250 244350
rect 562318 244294 562374 244350
rect 562442 244294 562498 244350
rect 562566 244294 562622 244350
rect 562194 244170 562250 244226
rect 562318 244170 562374 244226
rect 562442 244170 562498 244226
rect 562566 244170 562622 244226
rect 562194 244046 562250 244102
rect 562318 244046 562374 244102
rect 562442 244046 562498 244102
rect 562566 244046 562622 244102
rect 562194 243922 562250 243978
rect 562318 243922 562374 243978
rect 562442 243922 562498 243978
rect 562566 243922 562622 243978
rect 562194 226294 562250 226350
rect 562318 226294 562374 226350
rect 562442 226294 562498 226350
rect 562566 226294 562622 226350
rect 562194 226170 562250 226226
rect 562318 226170 562374 226226
rect 562442 226170 562498 226226
rect 562566 226170 562622 226226
rect 562194 226046 562250 226102
rect 562318 226046 562374 226102
rect 562442 226046 562498 226102
rect 562566 226046 562622 226102
rect 562194 225922 562250 225978
rect 562318 225922 562374 225978
rect 562442 225922 562498 225978
rect 562566 225922 562622 225978
rect 562194 208294 562250 208350
rect 562318 208294 562374 208350
rect 562442 208294 562498 208350
rect 562566 208294 562622 208350
rect 562194 208170 562250 208226
rect 562318 208170 562374 208226
rect 562442 208170 562498 208226
rect 562566 208170 562622 208226
rect 562194 208046 562250 208102
rect 562318 208046 562374 208102
rect 562442 208046 562498 208102
rect 562566 208046 562622 208102
rect 562194 207922 562250 207978
rect 562318 207922 562374 207978
rect 562442 207922 562498 207978
rect 562566 207922 562622 207978
rect 573238 202294 573294 202350
rect 573362 202294 573418 202350
rect 573238 202170 573294 202226
rect 573362 202170 573418 202226
rect 573238 202046 573294 202102
rect 573362 202046 573418 202102
rect 573238 201922 573294 201978
rect 573362 201922 573418 201978
rect 579740 192122 579796 192178
rect 562194 190294 562250 190350
rect 562318 190294 562374 190350
rect 562442 190294 562498 190350
rect 562566 190294 562622 190350
rect 562194 190170 562250 190226
rect 562318 190170 562374 190226
rect 562442 190170 562498 190226
rect 562566 190170 562622 190226
rect 562194 190046 562250 190102
rect 562318 190046 562374 190102
rect 562442 190046 562498 190102
rect 562566 190046 562622 190102
rect 562194 189922 562250 189978
rect 562318 189922 562374 189978
rect 562442 189922 562498 189978
rect 562566 189922 562622 189978
rect 573238 184294 573294 184350
rect 573362 184294 573418 184350
rect 573238 184170 573294 184226
rect 573362 184170 573418 184226
rect 573238 184046 573294 184102
rect 573362 184046 573418 184102
rect 573238 183922 573294 183978
rect 573362 183922 573418 183978
rect 562194 172294 562250 172350
rect 562318 172294 562374 172350
rect 562442 172294 562498 172350
rect 562566 172294 562622 172350
rect 562194 172170 562250 172226
rect 562318 172170 562374 172226
rect 562442 172170 562498 172226
rect 562566 172170 562622 172226
rect 562194 172046 562250 172102
rect 562318 172046 562374 172102
rect 562442 172046 562498 172102
rect 562566 172046 562622 172102
rect 562194 171922 562250 171978
rect 562318 171922 562374 171978
rect 562442 171922 562498 171978
rect 562566 171922 562622 171978
rect 562194 154294 562250 154350
rect 562318 154294 562374 154350
rect 562442 154294 562498 154350
rect 562566 154294 562622 154350
rect 562194 154170 562250 154226
rect 562318 154170 562374 154226
rect 562442 154170 562498 154226
rect 562566 154170 562622 154226
rect 562194 154046 562250 154102
rect 562318 154046 562374 154102
rect 562442 154046 562498 154102
rect 562566 154046 562622 154102
rect 562194 153922 562250 153978
rect 562318 153922 562374 153978
rect 562442 153922 562498 153978
rect 562566 153922 562622 153978
rect 562194 136294 562250 136350
rect 562318 136294 562374 136350
rect 562442 136294 562498 136350
rect 562566 136294 562622 136350
rect 562194 136170 562250 136226
rect 562318 136170 562374 136226
rect 562442 136170 562498 136226
rect 562566 136170 562622 136226
rect 562194 136046 562250 136102
rect 562318 136046 562374 136102
rect 562442 136046 562498 136102
rect 562566 136046 562622 136102
rect 562194 135922 562250 135978
rect 562318 135922 562374 135978
rect 562442 135922 562498 135978
rect 562566 135922 562622 135978
rect 573238 130294 573294 130350
rect 573362 130294 573418 130350
rect 573238 130170 573294 130226
rect 573362 130170 573418 130226
rect 573238 130046 573294 130102
rect 573362 130046 573418 130102
rect 573238 129922 573294 129978
rect 573362 129922 573418 129978
rect 562194 118294 562250 118350
rect 562318 118294 562374 118350
rect 562442 118294 562498 118350
rect 562566 118294 562622 118350
rect 562194 118170 562250 118226
rect 562318 118170 562374 118226
rect 562442 118170 562498 118226
rect 562566 118170 562622 118226
rect 562194 118046 562250 118102
rect 562318 118046 562374 118102
rect 562442 118046 562498 118102
rect 562566 118046 562622 118102
rect 562194 117922 562250 117978
rect 562318 117922 562374 117978
rect 562442 117922 562498 117978
rect 562566 117922 562622 117978
rect 573238 112294 573294 112350
rect 573362 112294 573418 112350
rect 573238 112170 573294 112226
rect 573362 112170 573418 112226
rect 573238 112046 573294 112102
rect 573362 112046 573418 112102
rect 573238 111922 573294 111978
rect 573362 111922 573418 111978
rect 562194 100294 562250 100350
rect 562318 100294 562374 100350
rect 562442 100294 562498 100350
rect 562566 100294 562622 100350
rect 562194 100170 562250 100226
rect 562318 100170 562374 100226
rect 562442 100170 562498 100226
rect 562566 100170 562622 100226
rect 562194 100046 562250 100102
rect 562318 100046 562374 100102
rect 562442 100046 562498 100102
rect 562566 100046 562622 100102
rect 562194 99922 562250 99978
rect 562318 99922 562374 99978
rect 562442 99922 562498 99978
rect 562566 99922 562622 99978
rect 562194 82294 562250 82350
rect 562318 82294 562374 82350
rect 562442 82294 562498 82350
rect 562566 82294 562622 82350
rect 562194 82170 562250 82226
rect 562318 82170 562374 82226
rect 562442 82170 562498 82226
rect 562566 82170 562622 82226
rect 562194 82046 562250 82102
rect 562318 82046 562374 82102
rect 562442 82046 562498 82102
rect 562566 82046 562622 82102
rect 562194 81922 562250 81978
rect 562318 81922 562374 81978
rect 562442 81922 562498 81978
rect 562566 81922 562622 81978
rect 562194 64294 562250 64350
rect 562318 64294 562374 64350
rect 562442 64294 562498 64350
rect 562566 64294 562622 64350
rect 562194 64170 562250 64226
rect 562318 64170 562374 64226
rect 562442 64170 562498 64226
rect 562566 64170 562622 64226
rect 562194 64046 562250 64102
rect 562318 64046 562374 64102
rect 562442 64046 562498 64102
rect 562566 64046 562622 64102
rect 562194 63922 562250 63978
rect 562318 63922 562374 63978
rect 562442 63922 562498 63978
rect 562566 63922 562622 63978
rect 557878 46294 557934 46350
rect 558002 46294 558058 46350
rect 557878 46170 557934 46226
rect 558002 46170 558058 46226
rect 557878 46046 557934 46102
rect 558002 46046 558058 46102
rect 557878 45922 557934 45978
rect 558002 45922 558058 45978
rect 573238 58294 573294 58350
rect 573362 58294 573418 58350
rect 573238 58170 573294 58226
rect 573362 58170 573418 58226
rect 573238 58046 573294 58102
rect 573362 58046 573418 58102
rect 573238 57922 573294 57978
rect 573362 57922 573418 57978
rect 562194 46294 562250 46350
rect 562318 46294 562374 46350
rect 562442 46294 562498 46350
rect 562566 46294 562622 46350
rect 562194 46170 562250 46226
rect 562318 46170 562374 46226
rect 562442 46170 562498 46226
rect 562566 46170 562622 46226
rect 562194 46046 562250 46102
rect 562318 46046 562374 46102
rect 562442 46046 562498 46102
rect 562566 46046 562622 46102
rect 562194 45922 562250 45978
rect 562318 45922 562374 45978
rect 562442 45922 562498 45978
rect 562566 45922 562622 45978
rect 542518 40294 542574 40350
rect 542642 40294 542698 40350
rect 542518 40170 542574 40226
rect 542642 40170 542698 40226
rect 542518 40046 542574 40102
rect 542642 40046 542698 40102
rect 542518 39922 542574 39978
rect 542642 39922 542698 39978
rect 558474 40294 558530 40350
rect 558598 40294 558654 40350
rect 558722 40294 558778 40350
rect 558846 40294 558902 40350
rect 558474 40170 558530 40226
rect 558598 40170 558654 40226
rect 558722 40170 558778 40226
rect 558846 40170 558902 40226
rect 558474 40046 558530 40102
rect 558598 40046 558654 40102
rect 558722 40046 558778 40102
rect 558846 40046 558902 40102
rect 558474 39922 558530 39978
rect 558598 39922 558654 39978
rect 558722 39922 558778 39978
rect 558846 39922 558902 39978
rect 531474 28294 531530 28350
rect 531598 28294 531654 28350
rect 531722 28294 531778 28350
rect 531846 28294 531902 28350
rect 531474 28170 531530 28226
rect 531598 28170 531654 28226
rect 531722 28170 531778 28226
rect 531846 28170 531902 28226
rect 531474 28046 531530 28102
rect 531598 28046 531654 28102
rect 531722 28046 531778 28102
rect 531846 28046 531902 28102
rect 531474 27922 531530 27978
rect 531598 27922 531654 27978
rect 531722 27922 531778 27978
rect 531846 27922 531902 27978
rect 531474 10294 531530 10350
rect 531598 10294 531654 10350
rect 531722 10294 531778 10350
rect 531846 10294 531902 10350
rect 531474 10170 531530 10226
rect 531598 10170 531654 10226
rect 531722 10170 531778 10226
rect 531846 10170 531902 10226
rect 531474 10046 531530 10102
rect 531598 10046 531654 10102
rect 531722 10046 531778 10102
rect 531846 10046 531902 10102
rect 531474 9922 531530 9978
rect 531598 9922 531654 9978
rect 531722 9922 531778 9978
rect 531846 9922 531902 9978
rect 531474 -1176 531530 -1120
rect 531598 -1176 531654 -1120
rect 531722 -1176 531778 -1120
rect 531846 -1176 531902 -1120
rect 531474 -1300 531530 -1244
rect 531598 -1300 531654 -1244
rect 531722 -1300 531778 -1244
rect 531846 -1300 531902 -1244
rect 531474 -1424 531530 -1368
rect 531598 -1424 531654 -1368
rect 531722 -1424 531778 -1368
rect 531846 -1424 531902 -1368
rect 531474 -1548 531530 -1492
rect 531598 -1548 531654 -1492
rect 531722 -1548 531778 -1492
rect 531846 -1548 531902 -1492
rect 558474 22294 558530 22350
rect 558598 22294 558654 22350
rect 558722 22294 558778 22350
rect 558846 22294 558902 22350
rect 558474 22170 558530 22226
rect 558598 22170 558654 22226
rect 558722 22170 558778 22226
rect 558846 22170 558902 22226
rect 558474 22046 558530 22102
rect 558598 22046 558654 22102
rect 558722 22046 558778 22102
rect 558846 22046 558902 22102
rect 558474 21922 558530 21978
rect 558598 21922 558654 21978
rect 558722 21922 558778 21978
rect 558846 21922 558902 21978
rect 558474 4294 558530 4350
rect 558598 4294 558654 4350
rect 558722 4294 558778 4350
rect 558846 4294 558902 4350
rect 558474 4170 558530 4226
rect 558598 4170 558654 4226
rect 558722 4170 558778 4226
rect 558846 4170 558902 4226
rect 558474 4046 558530 4102
rect 558598 4046 558654 4102
rect 558722 4046 558778 4102
rect 558846 4046 558902 4102
rect 558474 3922 558530 3978
rect 558598 3922 558654 3978
rect 558722 3922 558778 3978
rect 558846 3922 558902 3978
rect 558474 -216 558530 -160
rect 558598 -216 558654 -160
rect 558722 -216 558778 -160
rect 558846 -216 558902 -160
rect 558474 -340 558530 -284
rect 558598 -340 558654 -284
rect 558722 -340 558778 -284
rect 558846 -340 558902 -284
rect 558474 -464 558530 -408
rect 558598 -464 558654 -408
rect 558722 -464 558778 -408
rect 558846 -464 558902 -408
rect 558474 -588 558530 -532
rect 558598 -588 558654 -532
rect 558722 -588 558778 -532
rect 558846 -588 558902 -532
rect 573238 40294 573294 40350
rect 573362 40294 573418 40350
rect 573238 40170 573294 40226
rect 573362 40170 573418 40226
rect 573238 40046 573294 40102
rect 573362 40046 573418 40102
rect 573238 39922 573294 39978
rect 573362 39922 573418 39978
rect 589194 562294 589250 562350
rect 589318 562294 589374 562350
rect 589442 562294 589498 562350
rect 589566 562294 589622 562350
rect 589194 562170 589250 562226
rect 589318 562170 589374 562226
rect 589442 562170 589498 562226
rect 589566 562170 589622 562226
rect 589194 562046 589250 562102
rect 589318 562046 589374 562102
rect 589442 562046 589498 562102
rect 589566 562046 589622 562102
rect 589194 561922 589250 561978
rect 589318 561922 589374 561978
rect 589442 561922 589498 561978
rect 589566 561922 589622 561978
rect 589194 544294 589250 544350
rect 589318 544294 589374 544350
rect 589442 544294 589498 544350
rect 589566 544294 589622 544350
rect 589194 544170 589250 544226
rect 589318 544170 589374 544226
rect 589442 544170 589498 544226
rect 589566 544170 589622 544226
rect 589194 544046 589250 544102
rect 589318 544046 589374 544102
rect 589442 544046 589498 544102
rect 589566 544046 589622 544102
rect 589194 543922 589250 543978
rect 589318 543922 589374 543978
rect 589442 543922 589498 543978
rect 589566 543922 589622 543978
rect 589194 526294 589250 526350
rect 589318 526294 589374 526350
rect 589442 526294 589498 526350
rect 589566 526294 589622 526350
rect 589194 526170 589250 526226
rect 589318 526170 589374 526226
rect 589442 526170 589498 526226
rect 589566 526170 589622 526226
rect 589194 526046 589250 526102
rect 589318 526046 589374 526102
rect 589442 526046 589498 526102
rect 589566 526046 589622 526102
rect 589194 525922 589250 525978
rect 589318 525922 589374 525978
rect 589442 525922 589498 525978
rect 589566 525922 589622 525978
rect 589194 508294 589250 508350
rect 589318 508294 589374 508350
rect 589442 508294 589498 508350
rect 589566 508294 589622 508350
rect 589194 508170 589250 508226
rect 589318 508170 589374 508226
rect 589442 508170 589498 508226
rect 589566 508170 589622 508226
rect 589194 508046 589250 508102
rect 589318 508046 589374 508102
rect 589442 508046 589498 508102
rect 589566 508046 589622 508102
rect 589194 507922 589250 507978
rect 589318 507922 589374 507978
rect 589442 507922 589498 507978
rect 589566 507922 589622 507978
rect 589194 490294 589250 490350
rect 589318 490294 589374 490350
rect 589442 490294 589498 490350
rect 589566 490294 589622 490350
rect 589194 490170 589250 490226
rect 589318 490170 589374 490226
rect 589442 490170 589498 490226
rect 589566 490170 589622 490226
rect 589194 490046 589250 490102
rect 589318 490046 589374 490102
rect 589442 490046 589498 490102
rect 589566 490046 589622 490102
rect 589194 489922 589250 489978
rect 589318 489922 589374 489978
rect 589442 489922 589498 489978
rect 589566 489922 589622 489978
rect 589194 472294 589250 472350
rect 589318 472294 589374 472350
rect 589442 472294 589498 472350
rect 589566 472294 589622 472350
rect 589194 472170 589250 472226
rect 589318 472170 589374 472226
rect 589442 472170 589498 472226
rect 589566 472170 589622 472226
rect 589194 472046 589250 472102
rect 589318 472046 589374 472102
rect 589442 472046 589498 472102
rect 589566 472046 589622 472102
rect 589194 471922 589250 471978
rect 589318 471922 589374 471978
rect 589442 471922 589498 471978
rect 589566 471922 589622 471978
rect 589194 454294 589250 454350
rect 589318 454294 589374 454350
rect 589442 454294 589498 454350
rect 589566 454294 589622 454350
rect 589194 454170 589250 454226
rect 589318 454170 589374 454226
rect 589442 454170 589498 454226
rect 589566 454170 589622 454226
rect 589194 454046 589250 454102
rect 589318 454046 589374 454102
rect 589442 454046 589498 454102
rect 589566 454046 589622 454102
rect 589194 453922 589250 453978
rect 589318 453922 589374 453978
rect 589442 453922 589498 453978
rect 589566 453922 589622 453978
rect 589194 436294 589250 436350
rect 589318 436294 589374 436350
rect 589442 436294 589498 436350
rect 589566 436294 589622 436350
rect 589194 436170 589250 436226
rect 589318 436170 589374 436226
rect 589442 436170 589498 436226
rect 589566 436170 589622 436226
rect 589194 436046 589250 436102
rect 589318 436046 589374 436102
rect 589442 436046 589498 436102
rect 589566 436046 589622 436102
rect 589194 435922 589250 435978
rect 589318 435922 589374 435978
rect 589442 435922 589498 435978
rect 589566 435922 589622 435978
rect 589194 418294 589250 418350
rect 589318 418294 589374 418350
rect 589442 418294 589498 418350
rect 589566 418294 589622 418350
rect 589194 418170 589250 418226
rect 589318 418170 589374 418226
rect 589442 418170 589498 418226
rect 589566 418170 589622 418226
rect 589194 418046 589250 418102
rect 589318 418046 589374 418102
rect 589442 418046 589498 418102
rect 589566 418046 589622 418102
rect 589194 417922 589250 417978
rect 589318 417922 589374 417978
rect 589442 417922 589498 417978
rect 589566 417922 589622 417978
rect 589194 400294 589250 400350
rect 589318 400294 589374 400350
rect 589442 400294 589498 400350
rect 589566 400294 589622 400350
rect 589194 400170 589250 400226
rect 589318 400170 589374 400226
rect 589442 400170 589498 400226
rect 589566 400170 589622 400226
rect 589194 400046 589250 400102
rect 589318 400046 589374 400102
rect 589442 400046 589498 400102
rect 589566 400046 589622 400102
rect 589194 399922 589250 399978
rect 589318 399922 589374 399978
rect 589442 399922 589498 399978
rect 589566 399922 589622 399978
rect 589194 382294 589250 382350
rect 589318 382294 589374 382350
rect 589442 382294 589498 382350
rect 589566 382294 589622 382350
rect 589194 382170 589250 382226
rect 589318 382170 589374 382226
rect 589442 382170 589498 382226
rect 589566 382170 589622 382226
rect 589194 382046 589250 382102
rect 589318 382046 589374 382102
rect 589442 382046 589498 382102
rect 589566 382046 589622 382102
rect 589194 381922 589250 381978
rect 589318 381922 589374 381978
rect 589442 381922 589498 381978
rect 589566 381922 589622 381978
rect 589194 364294 589250 364350
rect 589318 364294 589374 364350
rect 589442 364294 589498 364350
rect 589566 364294 589622 364350
rect 589194 364170 589250 364226
rect 589318 364170 589374 364226
rect 589442 364170 589498 364226
rect 589566 364170 589622 364226
rect 589194 364046 589250 364102
rect 589318 364046 589374 364102
rect 589442 364046 589498 364102
rect 589566 364046 589622 364102
rect 589194 363922 589250 363978
rect 589318 363922 589374 363978
rect 589442 363922 589498 363978
rect 589566 363922 589622 363978
rect 589194 346294 589250 346350
rect 589318 346294 589374 346350
rect 589442 346294 589498 346350
rect 589566 346294 589622 346350
rect 589194 346170 589250 346226
rect 589318 346170 589374 346226
rect 589442 346170 589498 346226
rect 589566 346170 589622 346226
rect 589194 346046 589250 346102
rect 589318 346046 589374 346102
rect 589442 346046 589498 346102
rect 589566 346046 589622 346102
rect 589194 345922 589250 345978
rect 589318 345922 589374 345978
rect 589442 345922 589498 345978
rect 589566 345922 589622 345978
rect 589194 328294 589250 328350
rect 589318 328294 589374 328350
rect 589442 328294 589498 328350
rect 589566 328294 589622 328350
rect 589194 328170 589250 328226
rect 589318 328170 589374 328226
rect 589442 328170 589498 328226
rect 589566 328170 589622 328226
rect 589194 328046 589250 328102
rect 589318 328046 589374 328102
rect 589442 328046 589498 328102
rect 589566 328046 589622 328102
rect 589194 327922 589250 327978
rect 589318 327922 589374 327978
rect 589442 327922 589498 327978
rect 589566 327922 589622 327978
rect 589194 310294 589250 310350
rect 589318 310294 589374 310350
rect 589442 310294 589498 310350
rect 589566 310294 589622 310350
rect 589194 310170 589250 310226
rect 589318 310170 589374 310226
rect 589442 310170 589498 310226
rect 589566 310170 589622 310226
rect 589194 310046 589250 310102
rect 589318 310046 589374 310102
rect 589442 310046 589498 310102
rect 589566 310046 589622 310102
rect 589194 309922 589250 309978
rect 589318 309922 589374 309978
rect 589442 309922 589498 309978
rect 589566 309922 589622 309978
rect 589194 292294 589250 292350
rect 589318 292294 589374 292350
rect 589442 292294 589498 292350
rect 589566 292294 589622 292350
rect 589194 292170 589250 292226
rect 589318 292170 589374 292226
rect 589442 292170 589498 292226
rect 589566 292170 589622 292226
rect 589194 292046 589250 292102
rect 589318 292046 589374 292102
rect 589442 292046 589498 292102
rect 589566 292046 589622 292102
rect 589194 291922 589250 291978
rect 589318 291922 589374 291978
rect 589442 291922 589498 291978
rect 589566 291922 589622 291978
rect 589194 274294 589250 274350
rect 589318 274294 589374 274350
rect 589442 274294 589498 274350
rect 589566 274294 589622 274350
rect 589194 274170 589250 274226
rect 589318 274170 589374 274226
rect 589442 274170 589498 274226
rect 589566 274170 589622 274226
rect 589194 274046 589250 274102
rect 589318 274046 589374 274102
rect 589442 274046 589498 274102
rect 589566 274046 589622 274102
rect 589194 273922 589250 273978
rect 589318 273922 589374 273978
rect 589442 273922 589498 273978
rect 589566 273922 589622 273978
rect 589194 256294 589250 256350
rect 589318 256294 589374 256350
rect 589442 256294 589498 256350
rect 589566 256294 589622 256350
rect 589194 256170 589250 256226
rect 589318 256170 589374 256226
rect 589442 256170 589498 256226
rect 589566 256170 589622 256226
rect 589194 256046 589250 256102
rect 589318 256046 589374 256102
rect 589442 256046 589498 256102
rect 589566 256046 589622 256102
rect 589194 255922 589250 255978
rect 589318 255922 589374 255978
rect 589442 255922 589498 255978
rect 589566 255922 589622 255978
rect 589194 238294 589250 238350
rect 589318 238294 589374 238350
rect 589442 238294 589498 238350
rect 589566 238294 589622 238350
rect 589194 238170 589250 238226
rect 589318 238170 589374 238226
rect 589442 238170 589498 238226
rect 589566 238170 589622 238226
rect 589194 238046 589250 238102
rect 589318 238046 589374 238102
rect 589442 238046 589498 238102
rect 589566 238046 589622 238102
rect 589194 237922 589250 237978
rect 589318 237922 589374 237978
rect 589442 237922 589498 237978
rect 589566 237922 589622 237978
rect 589194 220294 589250 220350
rect 589318 220294 589374 220350
rect 589442 220294 589498 220350
rect 589566 220294 589622 220350
rect 589194 220170 589250 220226
rect 589318 220170 589374 220226
rect 589442 220170 589498 220226
rect 589566 220170 589622 220226
rect 589194 220046 589250 220102
rect 589318 220046 589374 220102
rect 589442 220046 589498 220102
rect 589566 220046 589622 220102
rect 589194 219922 589250 219978
rect 589318 219922 589374 219978
rect 589442 219922 589498 219978
rect 589566 219922 589622 219978
rect 589194 202294 589250 202350
rect 589318 202294 589374 202350
rect 589442 202294 589498 202350
rect 589566 202294 589622 202350
rect 589194 202170 589250 202226
rect 589318 202170 589374 202226
rect 589442 202170 589498 202226
rect 589566 202170 589622 202226
rect 589194 202046 589250 202102
rect 589318 202046 589374 202102
rect 589442 202046 589498 202102
rect 589566 202046 589622 202102
rect 589194 201922 589250 201978
rect 589318 201922 589374 201978
rect 589442 201922 589498 201978
rect 589566 201922 589622 201978
rect 589194 184294 589250 184350
rect 589318 184294 589374 184350
rect 589442 184294 589498 184350
rect 589566 184294 589622 184350
rect 589194 184170 589250 184226
rect 589318 184170 589374 184226
rect 589442 184170 589498 184226
rect 589566 184170 589622 184226
rect 589194 184046 589250 184102
rect 589318 184046 589374 184102
rect 589442 184046 589498 184102
rect 589566 184046 589622 184102
rect 589194 183922 589250 183978
rect 589318 183922 589374 183978
rect 589442 183922 589498 183978
rect 589566 183922 589622 183978
rect 589194 166294 589250 166350
rect 589318 166294 589374 166350
rect 589442 166294 589498 166350
rect 589566 166294 589622 166350
rect 589194 166170 589250 166226
rect 589318 166170 589374 166226
rect 589442 166170 589498 166226
rect 589566 166170 589622 166226
rect 589194 166046 589250 166102
rect 589318 166046 589374 166102
rect 589442 166046 589498 166102
rect 589566 166046 589622 166102
rect 589194 165922 589250 165978
rect 589318 165922 589374 165978
rect 589442 165922 589498 165978
rect 589566 165922 589622 165978
rect 589194 148294 589250 148350
rect 589318 148294 589374 148350
rect 589442 148294 589498 148350
rect 589566 148294 589622 148350
rect 589194 148170 589250 148226
rect 589318 148170 589374 148226
rect 589442 148170 589498 148226
rect 589566 148170 589622 148226
rect 589194 148046 589250 148102
rect 589318 148046 589374 148102
rect 589442 148046 589498 148102
rect 589566 148046 589622 148102
rect 589194 147922 589250 147978
rect 589318 147922 589374 147978
rect 589442 147922 589498 147978
rect 589566 147922 589622 147978
rect 589194 130294 589250 130350
rect 589318 130294 589374 130350
rect 589442 130294 589498 130350
rect 589566 130294 589622 130350
rect 589194 130170 589250 130226
rect 589318 130170 589374 130226
rect 589442 130170 589498 130226
rect 589566 130170 589622 130226
rect 589194 130046 589250 130102
rect 589318 130046 589374 130102
rect 589442 130046 589498 130102
rect 589566 130046 589622 130102
rect 589194 129922 589250 129978
rect 589318 129922 589374 129978
rect 589442 129922 589498 129978
rect 589566 129922 589622 129978
rect 589194 112294 589250 112350
rect 589318 112294 589374 112350
rect 589442 112294 589498 112350
rect 589566 112294 589622 112350
rect 589194 112170 589250 112226
rect 589318 112170 589374 112226
rect 589442 112170 589498 112226
rect 589566 112170 589622 112226
rect 589194 112046 589250 112102
rect 589318 112046 589374 112102
rect 589442 112046 589498 112102
rect 589566 112046 589622 112102
rect 589194 111922 589250 111978
rect 589318 111922 589374 111978
rect 589442 111922 589498 111978
rect 589566 111922 589622 111978
rect 589194 94294 589250 94350
rect 589318 94294 589374 94350
rect 589442 94294 589498 94350
rect 589566 94294 589622 94350
rect 589194 94170 589250 94226
rect 589318 94170 589374 94226
rect 589442 94170 589498 94226
rect 589566 94170 589622 94226
rect 589194 94046 589250 94102
rect 589318 94046 589374 94102
rect 589442 94046 589498 94102
rect 589566 94046 589622 94102
rect 589194 93922 589250 93978
rect 589318 93922 589374 93978
rect 589442 93922 589498 93978
rect 589566 93922 589622 93978
rect 589194 76294 589250 76350
rect 589318 76294 589374 76350
rect 589442 76294 589498 76350
rect 589566 76294 589622 76350
rect 589194 76170 589250 76226
rect 589318 76170 589374 76226
rect 589442 76170 589498 76226
rect 589566 76170 589622 76226
rect 589194 76046 589250 76102
rect 589318 76046 589374 76102
rect 589442 76046 589498 76102
rect 589566 76046 589622 76102
rect 589194 75922 589250 75978
rect 589318 75922 589374 75978
rect 589442 75922 589498 75978
rect 589566 75922 589622 75978
rect 589194 58294 589250 58350
rect 589318 58294 589374 58350
rect 589442 58294 589498 58350
rect 589566 58294 589622 58350
rect 589194 58170 589250 58226
rect 589318 58170 589374 58226
rect 589442 58170 589498 58226
rect 589566 58170 589622 58226
rect 589194 58046 589250 58102
rect 589318 58046 589374 58102
rect 589442 58046 589498 58102
rect 589566 58046 589622 58102
rect 589194 57922 589250 57978
rect 589318 57922 589374 57978
rect 589442 57922 589498 57978
rect 589566 57922 589622 57978
rect 589194 40294 589250 40350
rect 589318 40294 589374 40350
rect 589442 40294 589498 40350
rect 589566 40294 589622 40350
rect 589194 40170 589250 40226
rect 589318 40170 589374 40226
rect 589442 40170 589498 40226
rect 589566 40170 589622 40226
rect 589194 40046 589250 40102
rect 589318 40046 589374 40102
rect 589442 40046 589498 40102
rect 589566 40046 589622 40102
rect 589194 39922 589250 39978
rect 589318 39922 589374 39978
rect 589442 39922 589498 39978
rect 589566 39922 589622 39978
rect 562194 28294 562250 28350
rect 562318 28294 562374 28350
rect 562442 28294 562498 28350
rect 562566 28294 562622 28350
rect 562194 28170 562250 28226
rect 562318 28170 562374 28226
rect 562442 28170 562498 28226
rect 562566 28170 562622 28226
rect 562194 28046 562250 28102
rect 562318 28046 562374 28102
rect 562442 28046 562498 28102
rect 562566 28046 562622 28102
rect 562194 27922 562250 27978
rect 562318 27922 562374 27978
rect 562442 27922 562498 27978
rect 562566 27922 562622 27978
rect 562194 10294 562250 10350
rect 562318 10294 562374 10350
rect 562442 10294 562498 10350
rect 562566 10294 562622 10350
rect 562194 10170 562250 10226
rect 562318 10170 562374 10226
rect 562442 10170 562498 10226
rect 562566 10170 562622 10226
rect 562194 10046 562250 10102
rect 562318 10046 562374 10102
rect 562442 10046 562498 10102
rect 562566 10046 562622 10102
rect 562194 9922 562250 9978
rect 562318 9922 562374 9978
rect 562442 9922 562498 9978
rect 562566 9922 562622 9978
rect 562194 -1176 562250 -1120
rect 562318 -1176 562374 -1120
rect 562442 -1176 562498 -1120
rect 562566 -1176 562622 -1120
rect 562194 -1300 562250 -1244
rect 562318 -1300 562374 -1244
rect 562442 -1300 562498 -1244
rect 562566 -1300 562622 -1244
rect 562194 -1424 562250 -1368
rect 562318 -1424 562374 -1368
rect 562442 -1424 562498 -1368
rect 562566 -1424 562622 -1368
rect 562194 -1548 562250 -1492
rect 562318 -1548 562374 -1492
rect 562442 -1548 562498 -1492
rect 562566 -1548 562622 -1492
rect 589194 22294 589250 22350
rect 589318 22294 589374 22350
rect 589442 22294 589498 22350
rect 589566 22294 589622 22350
rect 589194 22170 589250 22226
rect 589318 22170 589374 22226
rect 589442 22170 589498 22226
rect 589566 22170 589622 22226
rect 589194 22046 589250 22102
rect 589318 22046 589374 22102
rect 589442 22046 589498 22102
rect 589566 22046 589622 22102
rect 589194 21922 589250 21978
rect 589318 21922 589374 21978
rect 589442 21922 589498 21978
rect 589566 21922 589622 21978
rect 589194 4294 589250 4350
rect 589318 4294 589374 4350
rect 589442 4294 589498 4350
rect 589566 4294 589622 4350
rect 589194 4170 589250 4226
rect 589318 4170 589374 4226
rect 589442 4170 589498 4226
rect 589566 4170 589622 4226
rect 589194 4046 589250 4102
rect 589318 4046 589374 4102
rect 589442 4046 589498 4102
rect 589566 4046 589622 4102
rect 589194 3922 589250 3978
rect 589318 3922 589374 3978
rect 589442 3922 589498 3978
rect 589566 3922 589622 3978
rect 589194 -216 589250 -160
rect 589318 -216 589374 -160
rect 589442 -216 589498 -160
rect 589566 -216 589622 -160
rect 589194 -340 589250 -284
rect 589318 -340 589374 -284
rect 589442 -340 589498 -284
rect 589566 -340 589622 -284
rect 589194 -464 589250 -408
rect 589318 -464 589374 -408
rect 589442 -464 589498 -408
rect 589566 -464 589622 -408
rect 589194 -588 589250 -532
rect 589318 -588 589374 -532
rect 589442 -588 589498 -532
rect 589566 -588 589622 -532
rect 592914 598116 592970 598172
rect 593038 598116 593094 598172
rect 593162 598116 593218 598172
rect 593286 598116 593342 598172
rect 592914 597992 592970 598048
rect 593038 597992 593094 598048
rect 593162 597992 593218 598048
rect 593286 597992 593342 598048
rect 592914 597868 592970 597924
rect 593038 597868 593094 597924
rect 593162 597868 593218 597924
rect 593286 597868 593342 597924
rect 592914 597744 592970 597800
rect 593038 597744 593094 597800
rect 593162 597744 593218 597800
rect 593286 597744 593342 597800
rect 597456 598116 597512 598172
rect 597580 598116 597636 598172
rect 597704 598116 597760 598172
rect 597828 598116 597884 598172
rect 597456 597992 597512 598048
rect 597580 597992 597636 598048
rect 597704 597992 597760 598048
rect 597828 597992 597884 598048
rect 597456 597868 597512 597924
rect 597580 597868 597636 597924
rect 597704 597868 597760 597924
rect 597828 597868 597884 597924
rect 597456 597744 597512 597800
rect 597580 597744 597636 597800
rect 597704 597744 597760 597800
rect 597828 597744 597884 597800
rect 592914 586294 592970 586350
rect 593038 586294 593094 586350
rect 593162 586294 593218 586350
rect 593286 586294 593342 586350
rect 592914 586170 592970 586226
rect 593038 586170 593094 586226
rect 593162 586170 593218 586226
rect 593286 586170 593342 586226
rect 592914 586046 592970 586102
rect 593038 586046 593094 586102
rect 593162 586046 593218 586102
rect 593286 586046 593342 586102
rect 592914 585922 592970 585978
rect 593038 585922 593094 585978
rect 593162 585922 593218 585978
rect 593286 585922 593342 585978
rect 592914 568294 592970 568350
rect 593038 568294 593094 568350
rect 593162 568294 593218 568350
rect 593286 568294 593342 568350
rect 592914 568170 592970 568226
rect 593038 568170 593094 568226
rect 593162 568170 593218 568226
rect 593286 568170 593342 568226
rect 592914 568046 592970 568102
rect 593038 568046 593094 568102
rect 593162 568046 593218 568102
rect 593286 568046 593342 568102
rect 592914 567922 592970 567978
rect 593038 567922 593094 567978
rect 593162 567922 593218 567978
rect 593286 567922 593342 567978
rect 592914 550294 592970 550350
rect 593038 550294 593094 550350
rect 593162 550294 593218 550350
rect 593286 550294 593342 550350
rect 592914 550170 592970 550226
rect 593038 550170 593094 550226
rect 593162 550170 593218 550226
rect 593286 550170 593342 550226
rect 592914 550046 592970 550102
rect 593038 550046 593094 550102
rect 593162 550046 593218 550102
rect 593286 550046 593342 550102
rect 592914 549922 592970 549978
rect 593038 549922 593094 549978
rect 593162 549922 593218 549978
rect 593286 549922 593342 549978
rect 592914 532294 592970 532350
rect 593038 532294 593094 532350
rect 593162 532294 593218 532350
rect 593286 532294 593342 532350
rect 592914 532170 592970 532226
rect 593038 532170 593094 532226
rect 593162 532170 593218 532226
rect 593286 532170 593342 532226
rect 592914 532046 592970 532102
rect 593038 532046 593094 532102
rect 593162 532046 593218 532102
rect 593286 532046 593342 532102
rect 592914 531922 592970 531978
rect 593038 531922 593094 531978
rect 593162 531922 593218 531978
rect 593286 531922 593342 531978
rect 592914 514294 592970 514350
rect 593038 514294 593094 514350
rect 593162 514294 593218 514350
rect 593286 514294 593342 514350
rect 592914 514170 592970 514226
rect 593038 514170 593094 514226
rect 593162 514170 593218 514226
rect 593286 514170 593342 514226
rect 592914 514046 592970 514102
rect 593038 514046 593094 514102
rect 593162 514046 593218 514102
rect 593286 514046 593342 514102
rect 592914 513922 592970 513978
rect 593038 513922 593094 513978
rect 593162 513922 593218 513978
rect 593286 513922 593342 513978
rect 592914 496294 592970 496350
rect 593038 496294 593094 496350
rect 593162 496294 593218 496350
rect 593286 496294 593342 496350
rect 592914 496170 592970 496226
rect 593038 496170 593094 496226
rect 593162 496170 593218 496226
rect 593286 496170 593342 496226
rect 592914 496046 592970 496102
rect 593038 496046 593094 496102
rect 593162 496046 593218 496102
rect 593286 496046 593342 496102
rect 592914 495922 592970 495978
rect 593038 495922 593094 495978
rect 593162 495922 593218 495978
rect 593286 495922 593342 495978
rect 592914 478294 592970 478350
rect 593038 478294 593094 478350
rect 593162 478294 593218 478350
rect 593286 478294 593342 478350
rect 592914 478170 592970 478226
rect 593038 478170 593094 478226
rect 593162 478170 593218 478226
rect 593286 478170 593342 478226
rect 592914 478046 592970 478102
rect 593038 478046 593094 478102
rect 593162 478046 593218 478102
rect 593286 478046 593342 478102
rect 592914 477922 592970 477978
rect 593038 477922 593094 477978
rect 593162 477922 593218 477978
rect 593286 477922 593342 477978
rect 592914 460294 592970 460350
rect 593038 460294 593094 460350
rect 593162 460294 593218 460350
rect 593286 460294 593342 460350
rect 592914 460170 592970 460226
rect 593038 460170 593094 460226
rect 593162 460170 593218 460226
rect 593286 460170 593342 460226
rect 592914 460046 592970 460102
rect 593038 460046 593094 460102
rect 593162 460046 593218 460102
rect 593286 460046 593342 460102
rect 592914 459922 592970 459978
rect 593038 459922 593094 459978
rect 593162 459922 593218 459978
rect 593286 459922 593342 459978
rect 592914 442294 592970 442350
rect 593038 442294 593094 442350
rect 593162 442294 593218 442350
rect 593286 442294 593342 442350
rect 592914 442170 592970 442226
rect 593038 442170 593094 442226
rect 593162 442170 593218 442226
rect 593286 442170 593342 442226
rect 592914 442046 592970 442102
rect 593038 442046 593094 442102
rect 593162 442046 593218 442102
rect 593286 442046 593342 442102
rect 592914 441922 592970 441978
rect 593038 441922 593094 441978
rect 593162 441922 593218 441978
rect 593286 441922 593342 441978
rect 592914 424294 592970 424350
rect 593038 424294 593094 424350
rect 593162 424294 593218 424350
rect 593286 424294 593342 424350
rect 592914 424170 592970 424226
rect 593038 424170 593094 424226
rect 593162 424170 593218 424226
rect 593286 424170 593342 424226
rect 592914 424046 592970 424102
rect 593038 424046 593094 424102
rect 593162 424046 593218 424102
rect 593286 424046 593342 424102
rect 592914 423922 592970 423978
rect 593038 423922 593094 423978
rect 593162 423922 593218 423978
rect 593286 423922 593342 423978
rect 592914 406294 592970 406350
rect 593038 406294 593094 406350
rect 593162 406294 593218 406350
rect 593286 406294 593342 406350
rect 592914 406170 592970 406226
rect 593038 406170 593094 406226
rect 593162 406170 593218 406226
rect 593286 406170 593342 406226
rect 592914 406046 592970 406102
rect 593038 406046 593094 406102
rect 593162 406046 593218 406102
rect 593286 406046 593342 406102
rect 592914 405922 592970 405978
rect 593038 405922 593094 405978
rect 593162 405922 593218 405978
rect 593286 405922 593342 405978
rect 592914 388294 592970 388350
rect 593038 388294 593094 388350
rect 593162 388294 593218 388350
rect 593286 388294 593342 388350
rect 592914 388170 592970 388226
rect 593038 388170 593094 388226
rect 593162 388170 593218 388226
rect 593286 388170 593342 388226
rect 592914 388046 592970 388102
rect 593038 388046 593094 388102
rect 593162 388046 593218 388102
rect 593286 388046 593342 388102
rect 592914 387922 592970 387978
rect 593038 387922 593094 387978
rect 593162 387922 593218 387978
rect 593286 387922 593342 387978
rect 592914 370294 592970 370350
rect 593038 370294 593094 370350
rect 593162 370294 593218 370350
rect 593286 370294 593342 370350
rect 592914 370170 592970 370226
rect 593038 370170 593094 370226
rect 593162 370170 593218 370226
rect 593286 370170 593342 370226
rect 592914 370046 592970 370102
rect 593038 370046 593094 370102
rect 593162 370046 593218 370102
rect 593286 370046 593342 370102
rect 592914 369922 592970 369978
rect 593038 369922 593094 369978
rect 593162 369922 593218 369978
rect 593286 369922 593342 369978
rect 592914 352294 592970 352350
rect 593038 352294 593094 352350
rect 593162 352294 593218 352350
rect 593286 352294 593342 352350
rect 592914 352170 592970 352226
rect 593038 352170 593094 352226
rect 593162 352170 593218 352226
rect 593286 352170 593342 352226
rect 592914 352046 592970 352102
rect 593038 352046 593094 352102
rect 593162 352046 593218 352102
rect 593286 352046 593342 352102
rect 592914 351922 592970 351978
rect 593038 351922 593094 351978
rect 593162 351922 593218 351978
rect 593286 351922 593342 351978
rect 592914 334294 592970 334350
rect 593038 334294 593094 334350
rect 593162 334294 593218 334350
rect 593286 334294 593342 334350
rect 592914 334170 592970 334226
rect 593038 334170 593094 334226
rect 593162 334170 593218 334226
rect 593286 334170 593342 334226
rect 592914 334046 592970 334102
rect 593038 334046 593094 334102
rect 593162 334046 593218 334102
rect 593286 334046 593342 334102
rect 592914 333922 592970 333978
rect 593038 333922 593094 333978
rect 593162 333922 593218 333978
rect 593286 333922 593342 333978
rect 592914 316294 592970 316350
rect 593038 316294 593094 316350
rect 593162 316294 593218 316350
rect 593286 316294 593342 316350
rect 592914 316170 592970 316226
rect 593038 316170 593094 316226
rect 593162 316170 593218 316226
rect 593286 316170 593342 316226
rect 592914 316046 592970 316102
rect 593038 316046 593094 316102
rect 593162 316046 593218 316102
rect 593286 316046 593342 316102
rect 592914 315922 592970 315978
rect 593038 315922 593094 315978
rect 593162 315922 593218 315978
rect 593286 315922 593342 315978
rect 592914 298294 592970 298350
rect 593038 298294 593094 298350
rect 593162 298294 593218 298350
rect 593286 298294 593342 298350
rect 592914 298170 592970 298226
rect 593038 298170 593094 298226
rect 593162 298170 593218 298226
rect 593286 298170 593342 298226
rect 592914 298046 592970 298102
rect 593038 298046 593094 298102
rect 593162 298046 593218 298102
rect 593286 298046 593342 298102
rect 592914 297922 592970 297978
rect 593038 297922 593094 297978
rect 593162 297922 593218 297978
rect 593286 297922 593342 297978
rect 592914 280294 592970 280350
rect 593038 280294 593094 280350
rect 593162 280294 593218 280350
rect 593286 280294 593342 280350
rect 592914 280170 592970 280226
rect 593038 280170 593094 280226
rect 593162 280170 593218 280226
rect 593286 280170 593342 280226
rect 592914 280046 592970 280102
rect 593038 280046 593094 280102
rect 593162 280046 593218 280102
rect 593286 280046 593342 280102
rect 592914 279922 592970 279978
rect 593038 279922 593094 279978
rect 593162 279922 593218 279978
rect 593286 279922 593342 279978
rect 592914 262294 592970 262350
rect 593038 262294 593094 262350
rect 593162 262294 593218 262350
rect 593286 262294 593342 262350
rect 592914 262170 592970 262226
rect 593038 262170 593094 262226
rect 593162 262170 593218 262226
rect 593286 262170 593342 262226
rect 592914 262046 592970 262102
rect 593038 262046 593094 262102
rect 593162 262046 593218 262102
rect 593286 262046 593342 262102
rect 592914 261922 592970 261978
rect 593038 261922 593094 261978
rect 593162 261922 593218 261978
rect 593286 261922 593342 261978
rect 592914 244294 592970 244350
rect 593038 244294 593094 244350
rect 593162 244294 593218 244350
rect 593286 244294 593342 244350
rect 592914 244170 592970 244226
rect 593038 244170 593094 244226
rect 593162 244170 593218 244226
rect 593286 244170 593342 244226
rect 592914 244046 592970 244102
rect 593038 244046 593094 244102
rect 593162 244046 593218 244102
rect 593286 244046 593342 244102
rect 592914 243922 592970 243978
rect 593038 243922 593094 243978
rect 593162 243922 593218 243978
rect 593286 243922 593342 243978
rect 592914 226294 592970 226350
rect 593038 226294 593094 226350
rect 593162 226294 593218 226350
rect 593286 226294 593342 226350
rect 592914 226170 592970 226226
rect 593038 226170 593094 226226
rect 593162 226170 593218 226226
rect 593286 226170 593342 226226
rect 592914 226046 592970 226102
rect 593038 226046 593094 226102
rect 593162 226046 593218 226102
rect 593286 226046 593342 226102
rect 592914 225922 592970 225978
rect 593038 225922 593094 225978
rect 593162 225922 593218 225978
rect 593286 225922 593342 225978
rect 592914 208294 592970 208350
rect 593038 208294 593094 208350
rect 593162 208294 593218 208350
rect 593286 208294 593342 208350
rect 592914 208170 592970 208226
rect 593038 208170 593094 208226
rect 593162 208170 593218 208226
rect 593286 208170 593342 208226
rect 592914 208046 592970 208102
rect 593038 208046 593094 208102
rect 593162 208046 593218 208102
rect 593286 208046 593342 208102
rect 592914 207922 592970 207978
rect 593038 207922 593094 207978
rect 593162 207922 593218 207978
rect 593286 207922 593342 207978
rect 592914 190294 592970 190350
rect 593038 190294 593094 190350
rect 593162 190294 593218 190350
rect 593286 190294 593342 190350
rect 592914 190170 592970 190226
rect 593038 190170 593094 190226
rect 593162 190170 593218 190226
rect 593286 190170 593342 190226
rect 592914 190046 592970 190102
rect 593038 190046 593094 190102
rect 593162 190046 593218 190102
rect 593286 190046 593342 190102
rect 592914 189922 592970 189978
rect 593038 189922 593094 189978
rect 593162 189922 593218 189978
rect 593286 189922 593342 189978
rect 592914 172294 592970 172350
rect 593038 172294 593094 172350
rect 593162 172294 593218 172350
rect 593286 172294 593342 172350
rect 592914 172170 592970 172226
rect 593038 172170 593094 172226
rect 593162 172170 593218 172226
rect 593286 172170 593342 172226
rect 592914 172046 592970 172102
rect 593038 172046 593094 172102
rect 593162 172046 593218 172102
rect 593286 172046 593342 172102
rect 592914 171922 592970 171978
rect 593038 171922 593094 171978
rect 593162 171922 593218 171978
rect 593286 171922 593342 171978
rect 592914 154294 592970 154350
rect 593038 154294 593094 154350
rect 593162 154294 593218 154350
rect 593286 154294 593342 154350
rect 592914 154170 592970 154226
rect 593038 154170 593094 154226
rect 593162 154170 593218 154226
rect 593286 154170 593342 154226
rect 592914 154046 592970 154102
rect 593038 154046 593094 154102
rect 593162 154046 593218 154102
rect 593286 154046 593342 154102
rect 592914 153922 592970 153978
rect 593038 153922 593094 153978
rect 593162 153922 593218 153978
rect 593286 153922 593342 153978
rect 592914 136294 592970 136350
rect 593038 136294 593094 136350
rect 593162 136294 593218 136350
rect 593286 136294 593342 136350
rect 592914 136170 592970 136226
rect 593038 136170 593094 136226
rect 593162 136170 593218 136226
rect 593286 136170 593342 136226
rect 592914 136046 592970 136102
rect 593038 136046 593094 136102
rect 593162 136046 593218 136102
rect 593286 136046 593342 136102
rect 592914 135922 592970 135978
rect 593038 135922 593094 135978
rect 593162 135922 593218 135978
rect 593286 135922 593342 135978
rect 592914 118294 592970 118350
rect 593038 118294 593094 118350
rect 593162 118294 593218 118350
rect 593286 118294 593342 118350
rect 592914 118170 592970 118226
rect 593038 118170 593094 118226
rect 593162 118170 593218 118226
rect 593286 118170 593342 118226
rect 592914 118046 592970 118102
rect 593038 118046 593094 118102
rect 593162 118046 593218 118102
rect 593286 118046 593342 118102
rect 592914 117922 592970 117978
rect 593038 117922 593094 117978
rect 593162 117922 593218 117978
rect 593286 117922 593342 117978
rect 592914 100294 592970 100350
rect 593038 100294 593094 100350
rect 593162 100294 593218 100350
rect 593286 100294 593342 100350
rect 592914 100170 592970 100226
rect 593038 100170 593094 100226
rect 593162 100170 593218 100226
rect 593286 100170 593342 100226
rect 592914 100046 592970 100102
rect 593038 100046 593094 100102
rect 593162 100046 593218 100102
rect 593286 100046 593342 100102
rect 592914 99922 592970 99978
rect 593038 99922 593094 99978
rect 593162 99922 593218 99978
rect 593286 99922 593342 99978
rect 592914 82294 592970 82350
rect 593038 82294 593094 82350
rect 593162 82294 593218 82350
rect 593286 82294 593342 82350
rect 592914 82170 592970 82226
rect 593038 82170 593094 82226
rect 593162 82170 593218 82226
rect 593286 82170 593342 82226
rect 592914 82046 592970 82102
rect 593038 82046 593094 82102
rect 593162 82046 593218 82102
rect 593286 82046 593342 82102
rect 592914 81922 592970 81978
rect 593038 81922 593094 81978
rect 593162 81922 593218 81978
rect 593286 81922 593342 81978
rect 592914 64294 592970 64350
rect 593038 64294 593094 64350
rect 593162 64294 593218 64350
rect 593286 64294 593342 64350
rect 592914 64170 592970 64226
rect 593038 64170 593094 64226
rect 593162 64170 593218 64226
rect 593286 64170 593342 64226
rect 592914 64046 592970 64102
rect 593038 64046 593094 64102
rect 593162 64046 593218 64102
rect 593286 64046 593342 64102
rect 592914 63922 592970 63978
rect 593038 63922 593094 63978
rect 593162 63922 593218 63978
rect 593286 63922 593342 63978
rect 592914 46294 592970 46350
rect 593038 46294 593094 46350
rect 593162 46294 593218 46350
rect 593286 46294 593342 46350
rect 592914 46170 592970 46226
rect 593038 46170 593094 46226
rect 593162 46170 593218 46226
rect 593286 46170 593342 46226
rect 592914 46046 592970 46102
rect 593038 46046 593094 46102
rect 593162 46046 593218 46102
rect 593286 46046 593342 46102
rect 592914 45922 592970 45978
rect 593038 45922 593094 45978
rect 593162 45922 593218 45978
rect 593286 45922 593342 45978
rect 592914 28294 592970 28350
rect 593038 28294 593094 28350
rect 593162 28294 593218 28350
rect 593286 28294 593342 28350
rect 592914 28170 592970 28226
rect 593038 28170 593094 28226
rect 593162 28170 593218 28226
rect 593286 28170 593342 28226
rect 592914 28046 592970 28102
rect 593038 28046 593094 28102
rect 593162 28046 593218 28102
rect 593286 28046 593342 28102
rect 592914 27922 592970 27978
rect 593038 27922 593094 27978
rect 593162 27922 593218 27978
rect 593286 27922 593342 27978
rect 592914 10294 592970 10350
rect 593038 10294 593094 10350
rect 593162 10294 593218 10350
rect 593286 10294 593342 10350
rect 592914 10170 592970 10226
rect 593038 10170 593094 10226
rect 593162 10170 593218 10226
rect 593286 10170 593342 10226
rect 592914 10046 592970 10102
rect 593038 10046 593094 10102
rect 593162 10046 593218 10102
rect 593286 10046 593342 10102
rect 592914 9922 592970 9978
rect 593038 9922 593094 9978
rect 593162 9922 593218 9978
rect 593286 9922 593342 9978
rect 596496 597156 596552 597212
rect 596620 597156 596676 597212
rect 596744 597156 596800 597212
rect 596868 597156 596924 597212
rect 596496 597032 596552 597088
rect 596620 597032 596676 597088
rect 596744 597032 596800 597088
rect 596868 597032 596924 597088
rect 596496 596908 596552 596964
rect 596620 596908 596676 596964
rect 596744 596908 596800 596964
rect 596868 596908 596924 596964
rect 596496 596784 596552 596840
rect 596620 596784 596676 596840
rect 596744 596784 596800 596840
rect 596868 596784 596924 596840
rect 596496 580294 596552 580350
rect 596620 580294 596676 580350
rect 596744 580294 596800 580350
rect 596868 580294 596924 580350
rect 596496 580170 596552 580226
rect 596620 580170 596676 580226
rect 596744 580170 596800 580226
rect 596868 580170 596924 580226
rect 596496 580046 596552 580102
rect 596620 580046 596676 580102
rect 596744 580046 596800 580102
rect 596868 580046 596924 580102
rect 596496 579922 596552 579978
rect 596620 579922 596676 579978
rect 596744 579922 596800 579978
rect 596868 579922 596924 579978
rect 596496 562294 596552 562350
rect 596620 562294 596676 562350
rect 596744 562294 596800 562350
rect 596868 562294 596924 562350
rect 596496 562170 596552 562226
rect 596620 562170 596676 562226
rect 596744 562170 596800 562226
rect 596868 562170 596924 562226
rect 596496 562046 596552 562102
rect 596620 562046 596676 562102
rect 596744 562046 596800 562102
rect 596868 562046 596924 562102
rect 596496 561922 596552 561978
rect 596620 561922 596676 561978
rect 596744 561922 596800 561978
rect 596868 561922 596924 561978
rect 596496 544294 596552 544350
rect 596620 544294 596676 544350
rect 596744 544294 596800 544350
rect 596868 544294 596924 544350
rect 596496 544170 596552 544226
rect 596620 544170 596676 544226
rect 596744 544170 596800 544226
rect 596868 544170 596924 544226
rect 596496 544046 596552 544102
rect 596620 544046 596676 544102
rect 596744 544046 596800 544102
rect 596868 544046 596924 544102
rect 596496 543922 596552 543978
rect 596620 543922 596676 543978
rect 596744 543922 596800 543978
rect 596868 543922 596924 543978
rect 596496 526294 596552 526350
rect 596620 526294 596676 526350
rect 596744 526294 596800 526350
rect 596868 526294 596924 526350
rect 596496 526170 596552 526226
rect 596620 526170 596676 526226
rect 596744 526170 596800 526226
rect 596868 526170 596924 526226
rect 596496 526046 596552 526102
rect 596620 526046 596676 526102
rect 596744 526046 596800 526102
rect 596868 526046 596924 526102
rect 596496 525922 596552 525978
rect 596620 525922 596676 525978
rect 596744 525922 596800 525978
rect 596868 525922 596924 525978
rect 596496 508294 596552 508350
rect 596620 508294 596676 508350
rect 596744 508294 596800 508350
rect 596868 508294 596924 508350
rect 596496 508170 596552 508226
rect 596620 508170 596676 508226
rect 596744 508170 596800 508226
rect 596868 508170 596924 508226
rect 596496 508046 596552 508102
rect 596620 508046 596676 508102
rect 596744 508046 596800 508102
rect 596868 508046 596924 508102
rect 596496 507922 596552 507978
rect 596620 507922 596676 507978
rect 596744 507922 596800 507978
rect 596868 507922 596924 507978
rect 596496 490294 596552 490350
rect 596620 490294 596676 490350
rect 596744 490294 596800 490350
rect 596868 490294 596924 490350
rect 596496 490170 596552 490226
rect 596620 490170 596676 490226
rect 596744 490170 596800 490226
rect 596868 490170 596924 490226
rect 596496 490046 596552 490102
rect 596620 490046 596676 490102
rect 596744 490046 596800 490102
rect 596868 490046 596924 490102
rect 596496 489922 596552 489978
rect 596620 489922 596676 489978
rect 596744 489922 596800 489978
rect 596868 489922 596924 489978
rect 596496 472294 596552 472350
rect 596620 472294 596676 472350
rect 596744 472294 596800 472350
rect 596868 472294 596924 472350
rect 596496 472170 596552 472226
rect 596620 472170 596676 472226
rect 596744 472170 596800 472226
rect 596868 472170 596924 472226
rect 596496 472046 596552 472102
rect 596620 472046 596676 472102
rect 596744 472046 596800 472102
rect 596868 472046 596924 472102
rect 596496 471922 596552 471978
rect 596620 471922 596676 471978
rect 596744 471922 596800 471978
rect 596868 471922 596924 471978
rect 596496 454294 596552 454350
rect 596620 454294 596676 454350
rect 596744 454294 596800 454350
rect 596868 454294 596924 454350
rect 596496 454170 596552 454226
rect 596620 454170 596676 454226
rect 596744 454170 596800 454226
rect 596868 454170 596924 454226
rect 596496 454046 596552 454102
rect 596620 454046 596676 454102
rect 596744 454046 596800 454102
rect 596868 454046 596924 454102
rect 596496 453922 596552 453978
rect 596620 453922 596676 453978
rect 596744 453922 596800 453978
rect 596868 453922 596924 453978
rect 596496 436294 596552 436350
rect 596620 436294 596676 436350
rect 596744 436294 596800 436350
rect 596868 436294 596924 436350
rect 596496 436170 596552 436226
rect 596620 436170 596676 436226
rect 596744 436170 596800 436226
rect 596868 436170 596924 436226
rect 596496 436046 596552 436102
rect 596620 436046 596676 436102
rect 596744 436046 596800 436102
rect 596868 436046 596924 436102
rect 596496 435922 596552 435978
rect 596620 435922 596676 435978
rect 596744 435922 596800 435978
rect 596868 435922 596924 435978
rect 596496 418294 596552 418350
rect 596620 418294 596676 418350
rect 596744 418294 596800 418350
rect 596868 418294 596924 418350
rect 596496 418170 596552 418226
rect 596620 418170 596676 418226
rect 596744 418170 596800 418226
rect 596868 418170 596924 418226
rect 596496 418046 596552 418102
rect 596620 418046 596676 418102
rect 596744 418046 596800 418102
rect 596868 418046 596924 418102
rect 596496 417922 596552 417978
rect 596620 417922 596676 417978
rect 596744 417922 596800 417978
rect 596868 417922 596924 417978
rect 596496 400294 596552 400350
rect 596620 400294 596676 400350
rect 596744 400294 596800 400350
rect 596868 400294 596924 400350
rect 596496 400170 596552 400226
rect 596620 400170 596676 400226
rect 596744 400170 596800 400226
rect 596868 400170 596924 400226
rect 596496 400046 596552 400102
rect 596620 400046 596676 400102
rect 596744 400046 596800 400102
rect 596868 400046 596924 400102
rect 596496 399922 596552 399978
rect 596620 399922 596676 399978
rect 596744 399922 596800 399978
rect 596868 399922 596924 399978
rect 596496 382294 596552 382350
rect 596620 382294 596676 382350
rect 596744 382294 596800 382350
rect 596868 382294 596924 382350
rect 596496 382170 596552 382226
rect 596620 382170 596676 382226
rect 596744 382170 596800 382226
rect 596868 382170 596924 382226
rect 596496 382046 596552 382102
rect 596620 382046 596676 382102
rect 596744 382046 596800 382102
rect 596868 382046 596924 382102
rect 596496 381922 596552 381978
rect 596620 381922 596676 381978
rect 596744 381922 596800 381978
rect 596868 381922 596924 381978
rect 596496 364294 596552 364350
rect 596620 364294 596676 364350
rect 596744 364294 596800 364350
rect 596868 364294 596924 364350
rect 596496 364170 596552 364226
rect 596620 364170 596676 364226
rect 596744 364170 596800 364226
rect 596868 364170 596924 364226
rect 596496 364046 596552 364102
rect 596620 364046 596676 364102
rect 596744 364046 596800 364102
rect 596868 364046 596924 364102
rect 596496 363922 596552 363978
rect 596620 363922 596676 363978
rect 596744 363922 596800 363978
rect 596868 363922 596924 363978
rect 596496 346294 596552 346350
rect 596620 346294 596676 346350
rect 596744 346294 596800 346350
rect 596868 346294 596924 346350
rect 596496 346170 596552 346226
rect 596620 346170 596676 346226
rect 596744 346170 596800 346226
rect 596868 346170 596924 346226
rect 596496 346046 596552 346102
rect 596620 346046 596676 346102
rect 596744 346046 596800 346102
rect 596868 346046 596924 346102
rect 596496 345922 596552 345978
rect 596620 345922 596676 345978
rect 596744 345922 596800 345978
rect 596868 345922 596924 345978
rect 596496 328294 596552 328350
rect 596620 328294 596676 328350
rect 596744 328294 596800 328350
rect 596868 328294 596924 328350
rect 596496 328170 596552 328226
rect 596620 328170 596676 328226
rect 596744 328170 596800 328226
rect 596868 328170 596924 328226
rect 596496 328046 596552 328102
rect 596620 328046 596676 328102
rect 596744 328046 596800 328102
rect 596868 328046 596924 328102
rect 596496 327922 596552 327978
rect 596620 327922 596676 327978
rect 596744 327922 596800 327978
rect 596868 327922 596924 327978
rect 596496 310294 596552 310350
rect 596620 310294 596676 310350
rect 596744 310294 596800 310350
rect 596868 310294 596924 310350
rect 596496 310170 596552 310226
rect 596620 310170 596676 310226
rect 596744 310170 596800 310226
rect 596868 310170 596924 310226
rect 596496 310046 596552 310102
rect 596620 310046 596676 310102
rect 596744 310046 596800 310102
rect 596868 310046 596924 310102
rect 596496 309922 596552 309978
rect 596620 309922 596676 309978
rect 596744 309922 596800 309978
rect 596868 309922 596924 309978
rect 596496 292294 596552 292350
rect 596620 292294 596676 292350
rect 596744 292294 596800 292350
rect 596868 292294 596924 292350
rect 596496 292170 596552 292226
rect 596620 292170 596676 292226
rect 596744 292170 596800 292226
rect 596868 292170 596924 292226
rect 596496 292046 596552 292102
rect 596620 292046 596676 292102
rect 596744 292046 596800 292102
rect 596868 292046 596924 292102
rect 596496 291922 596552 291978
rect 596620 291922 596676 291978
rect 596744 291922 596800 291978
rect 596868 291922 596924 291978
rect 596496 274294 596552 274350
rect 596620 274294 596676 274350
rect 596744 274294 596800 274350
rect 596868 274294 596924 274350
rect 596496 274170 596552 274226
rect 596620 274170 596676 274226
rect 596744 274170 596800 274226
rect 596868 274170 596924 274226
rect 596496 274046 596552 274102
rect 596620 274046 596676 274102
rect 596744 274046 596800 274102
rect 596868 274046 596924 274102
rect 596496 273922 596552 273978
rect 596620 273922 596676 273978
rect 596744 273922 596800 273978
rect 596868 273922 596924 273978
rect 596496 256294 596552 256350
rect 596620 256294 596676 256350
rect 596744 256294 596800 256350
rect 596868 256294 596924 256350
rect 596496 256170 596552 256226
rect 596620 256170 596676 256226
rect 596744 256170 596800 256226
rect 596868 256170 596924 256226
rect 596496 256046 596552 256102
rect 596620 256046 596676 256102
rect 596744 256046 596800 256102
rect 596868 256046 596924 256102
rect 596496 255922 596552 255978
rect 596620 255922 596676 255978
rect 596744 255922 596800 255978
rect 596868 255922 596924 255978
rect 596496 238294 596552 238350
rect 596620 238294 596676 238350
rect 596744 238294 596800 238350
rect 596868 238294 596924 238350
rect 596496 238170 596552 238226
rect 596620 238170 596676 238226
rect 596744 238170 596800 238226
rect 596868 238170 596924 238226
rect 596496 238046 596552 238102
rect 596620 238046 596676 238102
rect 596744 238046 596800 238102
rect 596868 238046 596924 238102
rect 596496 237922 596552 237978
rect 596620 237922 596676 237978
rect 596744 237922 596800 237978
rect 596868 237922 596924 237978
rect 596496 220294 596552 220350
rect 596620 220294 596676 220350
rect 596744 220294 596800 220350
rect 596868 220294 596924 220350
rect 596496 220170 596552 220226
rect 596620 220170 596676 220226
rect 596744 220170 596800 220226
rect 596868 220170 596924 220226
rect 596496 220046 596552 220102
rect 596620 220046 596676 220102
rect 596744 220046 596800 220102
rect 596868 220046 596924 220102
rect 596496 219922 596552 219978
rect 596620 219922 596676 219978
rect 596744 219922 596800 219978
rect 596868 219922 596924 219978
rect 596496 202294 596552 202350
rect 596620 202294 596676 202350
rect 596744 202294 596800 202350
rect 596868 202294 596924 202350
rect 596496 202170 596552 202226
rect 596620 202170 596676 202226
rect 596744 202170 596800 202226
rect 596868 202170 596924 202226
rect 596496 202046 596552 202102
rect 596620 202046 596676 202102
rect 596744 202046 596800 202102
rect 596868 202046 596924 202102
rect 596496 201922 596552 201978
rect 596620 201922 596676 201978
rect 596744 201922 596800 201978
rect 596868 201922 596924 201978
rect 596496 184294 596552 184350
rect 596620 184294 596676 184350
rect 596744 184294 596800 184350
rect 596868 184294 596924 184350
rect 596496 184170 596552 184226
rect 596620 184170 596676 184226
rect 596744 184170 596800 184226
rect 596868 184170 596924 184226
rect 596496 184046 596552 184102
rect 596620 184046 596676 184102
rect 596744 184046 596800 184102
rect 596868 184046 596924 184102
rect 596496 183922 596552 183978
rect 596620 183922 596676 183978
rect 596744 183922 596800 183978
rect 596868 183922 596924 183978
rect 596496 166294 596552 166350
rect 596620 166294 596676 166350
rect 596744 166294 596800 166350
rect 596868 166294 596924 166350
rect 596496 166170 596552 166226
rect 596620 166170 596676 166226
rect 596744 166170 596800 166226
rect 596868 166170 596924 166226
rect 596496 166046 596552 166102
rect 596620 166046 596676 166102
rect 596744 166046 596800 166102
rect 596868 166046 596924 166102
rect 596496 165922 596552 165978
rect 596620 165922 596676 165978
rect 596744 165922 596800 165978
rect 596868 165922 596924 165978
rect 596496 148294 596552 148350
rect 596620 148294 596676 148350
rect 596744 148294 596800 148350
rect 596868 148294 596924 148350
rect 596496 148170 596552 148226
rect 596620 148170 596676 148226
rect 596744 148170 596800 148226
rect 596868 148170 596924 148226
rect 596496 148046 596552 148102
rect 596620 148046 596676 148102
rect 596744 148046 596800 148102
rect 596868 148046 596924 148102
rect 596496 147922 596552 147978
rect 596620 147922 596676 147978
rect 596744 147922 596800 147978
rect 596868 147922 596924 147978
rect 596496 130294 596552 130350
rect 596620 130294 596676 130350
rect 596744 130294 596800 130350
rect 596868 130294 596924 130350
rect 596496 130170 596552 130226
rect 596620 130170 596676 130226
rect 596744 130170 596800 130226
rect 596868 130170 596924 130226
rect 596496 130046 596552 130102
rect 596620 130046 596676 130102
rect 596744 130046 596800 130102
rect 596868 130046 596924 130102
rect 596496 129922 596552 129978
rect 596620 129922 596676 129978
rect 596744 129922 596800 129978
rect 596868 129922 596924 129978
rect 596496 112294 596552 112350
rect 596620 112294 596676 112350
rect 596744 112294 596800 112350
rect 596868 112294 596924 112350
rect 596496 112170 596552 112226
rect 596620 112170 596676 112226
rect 596744 112170 596800 112226
rect 596868 112170 596924 112226
rect 596496 112046 596552 112102
rect 596620 112046 596676 112102
rect 596744 112046 596800 112102
rect 596868 112046 596924 112102
rect 596496 111922 596552 111978
rect 596620 111922 596676 111978
rect 596744 111922 596800 111978
rect 596868 111922 596924 111978
rect 596496 94294 596552 94350
rect 596620 94294 596676 94350
rect 596744 94294 596800 94350
rect 596868 94294 596924 94350
rect 596496 94170 596552 94226
rect 596620 94170 596676 94226
rect 596744 94170 596800 94226
rect 596868 94170 596924 94226
rect 596496 94046 596552 94102
rect 596620 94046 596676 94102
rect 596744 94046 596800 94102
rect 596868 94046 596924 94102
rect 596496 93922 596552 93978
rect 596620 93922 596676 93978
rect 596744 93922 596800 93978
rect 596868 93922 596924 93978
rect 596496 76294 596552 76350
rect 596620 76294 596676 76350
rect 596744 76294 596800 76350
rect 596868 76294 596924 76350
rect 596496 76170 596552 76226
rect 596620 76170 596676 76226
rect 596744 76170 596800 76226
rect 596868 76170 596924 76226
rect 596496 76046 596552 76102
rect 596620 76046 596676 76102
rect 596744 76046 596800 76102
rect 596868 76046 596924 76102
rect 596496 75922 596552 75978
rect 596620 75922 596676 75978
rect 596744 75922 596800 75978
rect 596868 75922 596924 75978
rect 596496 58294 596552 58350
rect 596620 58294 596676 58350
rect 596744 58294 596800 58350
rect 596868 58294 596924 58350
rect 596496 58170 596552 58226
rect 596620 58170 596676 58226
rect 596744 58170 596800 58226
rect 596868 58170 596924 58226
rect 596496 58046 596552 58102
rect 596620 58046 596676 58102
rect 596744 58046 596800 58102
rect 596868 58046 596924 58102
rect 596496 57922 596552 57978
rect 596620 57922 596676 57978
rect 596744 57922 596800 57978
rect 596868 57922 596924 57978
rect 596496 40294 596552 40350
rect 596620 40294 596676 40350
rect 596744 40294 596800 40350
rect 596868 40294 596924 40350
rect 596496 40170 596552 40226
rect 596620 40170 596676 40226
rect 596744 40170 596800 40226
rect 596868 40170 596924 40226
rect 596496 40046 596552 40102
rect 596620 40046 596676 40102
rect 596744 40046 596800 40102
rect 596868 40046 596924 40102
rect 596496 39922 596552 39978
rect 596620 39922 596676 39978
rect 596744 39922 596800 39978
rect 596868 39922 596924 39978
rect 596496 22294 596552 22350
rect 596620 22294 596676 22350
rect 596744 22294 596800 22350
rect 596868 22294 596924 22350
rect 596496 22170 596552 22226
rect 596620 22170 596676 22226
rect 596744 22170 596800 22226
rect 596868 22170 596924 22226
rect 596496 22046 596552 22102
rect 596620 22046 596676 22102
rect 596744 22046 596800 22102
rect 596868 22046 596924 22102
rect 596496 21922 596552 21978
rect 596620 21922 596676 21978
rect 596744 21922 596800 21978
rect 596868 21922 596924 21978
rect 596496 4294 596552 4350
rect 596620 4294 596676 4350
rect 596744 4294 596800 4350
rect 596868 4294 596924 4350
rect 596496 4170 596552 4226
rect 596620 4170 596676 4226
rect 596744 4170 596800 4226
rect 596868 4170 596924 4226
rect 596496 4046 596552 4102
rect 596620 4046 596676 4102
rect 596744 4046 596800 4102
rect 596868 4046 596924 4102
rect 596496 3922 596552 3978
rect 596620 3922 596676 3978
rect 596744 3922 596800 3978
rect 596868 3922 596924 3978
rect 596496 -216 596552 -160
rect 596620 -216 596676 -160
rect 596744 -216 596800 -160
rect 596868 -216 596924 -160
rect 596496 -340 596552 -284
rect 596620 -340 596676 -284
rect 596744 -340 596800 -284
rect 596868 -340 596924 -284
rect 596496 -464 596552 -408
rect 596620 -464 596676 -408
rect 596744 -464 596800 -408
rect 596868 -464 596924 -408
rect 596496 -588 596552 -532
rect 596620 -588 596676 -532
rect 596744 -588 596800 -532
rect 596868 -588 596924 -532
rect 597456 586294 597512 586350
rect 597580 586294 597636 586350
rect 597704 586294 597760 586350
rect 597828 586294 597884 586350
rect 597456 586170 597512 586226
rect 597580 586170 597636 586226
rect 597704 586170 597760 586226
rect 597828 586170 597884 586226
rect 597456 586046 597512 586102
rect 597580 586046 597636 586102
rect 597704 586046 597760 586102
rect 597828 586046 597884 586102
rect 597456 585922 597512 585978
rect 597580 585922 597636 585978
rect 597704 585922 597760 585978
rect 597828 585922 597884 585978
rect 597456 568294 597512 568350
rect 597580 568294 597636 568350
rect 597704 568294 597760 568350
rect 597828 568294 597884 568350
rect 597456 568170 597512 568226
rect 597580 568170 597636 568226
rect 597704 568170 597760 568226
rect 597828 568170 597884 568226
rect 597456 568046 597512 568102
rect 597580 568046 597636 568102
rect 597704 568046 597760 568102
rect 597828 568046 597884 568102
rect 597456 567922 597512 567978
rect 597580 567922 597636 567978
rect 597704 567922 597760 567978
rect 597828 567922 597884 567978
rect 597456 550294 597512 550350
rect 597580 550294 597636 550350
rect 597704 550294 597760 550350
rect 597828 550294 597884 550350
rect 597456 550170 597512 550226
rect 597580 550170 597636 550226
rect 597704 550170 597760 550226
rect 597828 550170 597884 550226
rect 597456 550046 597512 550102
rect 597580 550046 597636 550102
rect 597704 550046 597760 550102
rect 597828 550046 597884 550102
rect 597456 549922 597512 549978
rect 597580 549922 597636 549978
rect 597704 549922 597760 549978
rect 597828 549922 597884 549978
rect 597456 532294 597512 532350
rect 597580 532294 597636 532350
rect 597704 532294 597760 532350
rect 597828 532294 597884 532350
rect 597456 532170 597512 532226
rect 597580 532170 597636 532226
rect 597704 532170 597760 532226
rect 597828 532170 597884 532226
rect 597456 532046 597512 532102
rect 597580 532046 597636 532102
rect 597704 532046 597760 532102
rect 597828 532046 597884 532102
rect 597456 531922 597512 531978
rect 597580 531922 597636 531978
rect 597704 531922 597760 531978
rect 597828 531922 597884 531978
rect 597456 514294 597512 514350
rect 597580 514294 597636 514350
rect 597704 514294 597760 514350
rect 597828 514294 597884 514350
rect 597456 514170 597512 514226
rect 597580 514170 597636 514226
rect 597704 514170 597760 514226
rect 597828 514170 597884 514226
rect 597456 514046 597512 514102
rect 597580 514046 597636 514102
rect 597704 514046 597760 514102
rect 597828 514046 597884 514102
rect 597456 513922 597512 513978
rect 597580 513922 597636 513978
rect 597704 513922 597760 513978
rect 597828 513922 597884 513978
rect 597456 496294 597512 496350
rect 597580 496294 597636 496350
rect 597704 496294 597760 496350
rect 597828 496294 597884 496350
rect 597456 496170 597512 496226
rect 597580 496170 597636 496226
rect 597704 496170 597760 496226
rect 597828 496170 597884 496226
rect 597456 496046 597512 496102
rect 597580 496046 597636 496102
rect 597704 496046 597760 496102
rect 597828 496046 597884 496102
rect 597456 495922 597512 495978
rect 597580 495922 597636 495978
rect 597704 495922 597760 495978
rect 597828 495922 597884 495978
rect 597456 478294 597512 478350
rect 597580 478294 597636 478350
rect 597704 478294 597760 478350
rect 597828 478294 597884 478350
rect 597456 478170 597512 478226
rect 597580 478170 597636 478226
rect 597704 478170 597760 478226
rect 597828 478170 597884 478226
rect 597456 478046 597512 478102
rect 597580 478046 597636 478102
rect 597704 478046 597760 478102
rect 597828 478046 597884 478102
rect 597456 477922 597512 477978
rect 597580 477922 597636 477978
rect 597704 477922 597760 477978
rect 597828 477922 597884 477978
rect 597456 460294 597512 460350
rect 597580 460294 597636 460350
rect 597704 460294 597760 460350
rect 597828 460294 597884 460350
rect 597456 460170 597512 460226
rect 597580 460170 597636 460226
rect 597704 460170 597760 460226
rect 597828 460170 597884 460226
rect 597456 460046 597512 460102
rect 597580 460046 597636 460102
rect 597704 460046 597760 460102
rect 597828 460046 597884 460102
rect 597456 459922 597512 459978
rect 597580 459922 597636 459978
rect 597704 459922 597760 459978
rect 597828 459922 597884 459978
rect 597456 442294 597512 442350
rect 597580 442294 597636 442350
rect 597704 442294 597760 442350
rect 597828 442294 597884 442350
rect 597456 442170 597512 442226
rect 597580 442170 597636 442226
rect 597704 442170 597760 442226
rect 597828 442170 597884 442226
rect 597456 442046 597512 442102
rect 597580 442046 597636 442102
rect 597704 442046 597760 442102
rect 597828 442046 597884 442102
rect 597456 441922 597512 441978
rect 597580 441922 597636 441978
rect 597704 441922 597760 441978
rect 597828 441922 597884 441978
rect 597456 424294 597512 424350
rect 597580 424294 597636 424350
rect 597704 424294 597760 424350
rect 597828 424294 597884 424350
rect 597456 424170 597512 424226
rect 597580 424170 597636 424226
rect 597704 424170 597760 424226
rect 597828 424170 597884 424226
rect 597456 424046 597512 424102
rect 597580 424046 597636 424102
rect 597704 424046 597760 424102
rect 597828 424046 597884 424102
rect 597456 423922 597512 423978
rect 597580 423922 597636 423978
rect 597704 423922 597760 423978
rect 597828 423922 597884 423978
rect 597456 406294 597512 406350
rect 597580 406294 597636 406350
rect 597704 406294 597760 406350
rect 597828 406294 597884 406350
rect 597456 406170 597512 406226
rect 597580 406170 597636 406226
rect 597704 406170 597760 406226
rect 597828 406170 597884 406226
rect 597456 406046 597512 406102
rect 597580 406046 597636 406102
rect 597704 406046 597760 406102
rect 597828 406046 597884 406102
rect 597456 405922 597512 405978
rect 597580 405922 597636 405978
rect 597704 405922 597760 405978
rect 597828 405922 597884 405978
rect 597456 388294 597512 388350
rect 597580 388294 597636 388350
rect 597704 388294 597760 388350
rect 597828 388294 597884 388350
rect 597456 388170 597512 388226
rect 597580 388170 597636 388226
rect 597704 388170 597760 388226
rect 597828 388170 597884 388226
rect 597456 388046 597512 388102
rect 597580 388046 597636 388102
rect 597704 388046 597760 388102
rect 597828 388046 597884 388102
rect 597456 387922 597512 387978
rect 597580 387922 597636 387978
rect 597704 387922 597760 387978
rect 597828 387922 597884 387978
rect 597456 370294 597512 370350
rect 597580 370294 597636 370350
rect 597704 370294 597760 370350
rect 597828 370294 597884 370350
rect 597456 370170 597512 370226
rect 597580 370170 597636 370226
rect 597704 370170 597760 370226
rect 597828 370170 597884 370226
rect 597456 370046 597512 370102
rect 597580 370046 597636 370102
rect 597704 370046 597760 370102
rect 597828 370046 597884 370102
rect 597456 369922 597512 369978
rect 597580 369922 597636 369978
rect 597704 369922 597760 369978
rect 597828 369922 597884 369978
rect 597456 352294 597512 352350
rect 597580 352294 597636 352350
rect 597704 352294 597760 352350
rect 597828 352294 597884 352350
rect 597456 352170 597512 352226
rect 597580 352170 597636 352226
rect 597704 352170 597760 352226
rect 597828 352170 597884 352226
rect 597456 352046 597512 352102
rect 597580 352046 597636 352102
rect 597704 352046 597760 352102
rect 597828 352046 597884 352102
rect 597456 351922 597512 351978
rect 597580 351922 597636 351978
rect 597704 351922 597760 351978
rect 597828 351922 597884 351978
rect 597456 334294 597512 334350
rect 597580 334294 597636 334350
rect 597704 334294 597760 334350
rect 597828 334294 597884 334350
rect 597456 334170 597512 334226
rect 597580 334170 597636 334226
rect 597704 334170 597760 334226
rect 597828 334170 597884 334226
rect 597456 334046 597512 334102
rect 597580 334046 597636 334102
rect 597704 334046 597760 334102
rect 597828 334046 597884 334102
rect 597456 333922 597512 333978
rect 597580 333922 597636 333978
rect 597704 333922 597760 333978
rect 597828 333922 597884 333978
rect 597456 316294 597512 316350
rect 597580 316294 597636 316350
rect 597704 316294 597760 316350
rect 597828 316294 597884 316350
rect 597456 316170 597512 316226
rect 597580 316170 597636 316226
rect 597704 316170 597760 316226
rect 597828 316170 597884 316226
rect 597456 316046 597512 316102
rect 597580 316046 597636 316102
rect 597704 316046 597760 316102
rect 597828 316046 597884 316102
rect 597456 315922 597512 315978
rect 597580 315922 597636 315978
rect 597704 315922 597760 315978
rect 597828 315922 597884 315978
rect 597456 298294 597512 298350
rect 597580 298294 597636 298350
rect 597704 298294 597760 298350
rect 597828 298294 597884 298350
rect 597456 298170 597512 298226
rect 597580 298170 597636 298226
rect 597704 298170 597760 298226
rect 597828 298170 597884 298226
rect 597456 298046 597512 298102
rect 597580 298046 597636 298102
rect 597704 298046 597760 298102
rect 597828 298046 597884 298102
rect 597456 297922 597512 297978
rect 597580 297922 597636 297978
rect 597704 297922 597760 297978
rect 597828 297922 597884 297978
rect 597456 280294 597512 280350
rect 597580 280294 597636 280350
rect 597704 280294 597760 280350
rect 597828 280294 597884 280350
rect 597456 280170 597512 280226
rect 597580 280170 597636 280226
rect 597704 280170 597760 280226
rect 597828 280170 597884 280226
rect 597456 280046 597512 280102
rect 597580 280046 597636 280102
rect 597704 280046 597760 280102
rect 597828 280046 597884 280102
rect 597456 279922 597512 279978
rect 597580 279922 597636 279978
rect 597704 279922 597760 279978
rect 597828 279922 597884 279978
rect 597456 262294 597512 262350
rect 597580 262294 597636 262350
rect 597704 262294 597760 262350
rect 597828 262294 597884 262350
rect 597456 262170 597512 262226
rect 597580 262170 597636 262226
rect 597704 262170 597760 262226
rect 597828 262170 597884 262226
rect 597456 262046 597512 262102
rect 597580 262046 597636 262102
rect 597704 262046 597760 262102
rect 597828 262046 597884 262102
rect 597456 261922 597512 261978
rect 597580 261922 597636 261978
rect 597704 261922 597760 261978
rect 597828 261922 597884 261978
rect 597456 244294 597512 244350
rect 597580 244294 597636 244350
rect 597704 244294 597760 244350
rect 597828 244294 597884 244350
rect 597456 244170 597512 244226
rect 597580 244170 597636 244226
rect 597704 244170 597760 244226
rect 597828 244170 597884 244226
rect 597456 244046 597512 244102
rect 597580 244046 597636 244102
rect 597704 244046 597760 244102
rect 597828 244046 597884 244102
rect 597456 243922 597512 243978
rect 597580 243922 597636 243978
rect 597704 243922 597760 243978
rect 597828 243922 597884 243978
rect 597456 226294 597512 226350
rect 597580 226294 597636 226350
rect 597704 226294 597760 226350
rect 597828 226294 597884 226350
rect 597456 226170 597512 226226
rect 597580 226170 597636 226226
rect 597704 226170 597760 226226
rect 597828 226170 597884 226226
rect 597456 226046 597512 226102
rect 597580 226046 597636 226102
rect 597704 226046 597760 226102
rect 597828 226046 597884 226102
rect 597456 225922 597512 225978
rect 597580 225922 597636 225978
rect 597704 225922 597760 225978
rect 597828 225922 597884 225978
rect 597456 208294 597512 208350
rect 597580 208294 597636 208350
rect 597704 208294 597760 208350
rect 597828 208294 597884 208350
rect 597456 208170 597512 208226
rect 597580 208170 597636 208226
rect 597704 208170 597760 208226
rect 597828 208170 597884 208226
rect 597456 208046 597512 208102
rect 597580 208046 597636 208102
rect 597704 208046 597760 208102
rect 597828 208046 597884 208102
rect 597456 207922 597512 207978
rect 597580 207922 597636 207978
rect 597704 207922 597760 207978
rect 597828 207922 597884 207978
rect 597456 190294 597512 190350
rect 597580 190294 597636 190350
rect 597704 190294 597760 190350
rect 597828 190294 597884 190350
rect 597456 190170 597512 190226
rect 597580 190170 597636 190226
rect 597704 190170 597760 190226
rect 597828 190170 597884 190226
rect 597456 190046 597512 190102
rect 597580 190046 597636 190102
rect 597704 190046 597760 190102
rect 597828 190046 597884 190102
rect 597456 189922 597512 189978
rect 597580 189922 597636 189978
rect 597704 189922 597760 189978
rect 597828 189922 597884 189978
rect 597456 172294 597512 172350
rect 597580 172294 597636 172350
rect 597704 172294 597760 172350
rect 597828 172294 597884 172350
rect 597456 172170 597512 172226
rect 597580 172170 597636 172226
rect 597704 172170 597760 172226
rect 597828 172170 597884 172226
rect 597456 172046 597512 172102
rect 597580 172046 597636 172102
rect 597704 172046 597760 172102
rect 597828 172046 597884 172102
rect 597456 171922 597512 171978
rect 597580 171922 597636 171978
rect 597704 171922 597760 171978
rect 597828 171922 597884 171978
rect 597456 154294 597512 154350
rect 597580 154294 597636 154350
rect 597704 154294 597760 154350
rect 597828 154294 597884 154350
rect 597456 154170 597512 154226
rect 597580 154170 597636 154226
rect 597704 154170 597760 154226
rect 597828 154170 597884 154226
rect 597456 154046 597512 154102
rect 597580 154046 597636 154102
rect 597704 154046 597760 154102
rect 597828 154046 597884 154102
rect 597456 153922 597512 153978
rect 597580 153922 597636 153978
rect 597704 153922 597760 153978
rect 597828 153922 597884 153978
rect 597456 136294 597512 136350
rect 597580 136294 597636 136350
rect 597704 136294 597760 136350
rect 597828 136294 597884 136350
rect 597456 136170 597512 136226
rect 597580 136170 597636 136226
rect 597704 136170 597760 136226
rect 597828 136170 597884 136226
rect 597456 136046 597512 136102
rect 597580 136046 597636 136102
rect 597704 136046 597760 136102
rect 597828 136046 597884 136102
rect 597456 135922 597512 135978
rect 597580 135922 597636 135978
rect 597704 135922 597760 135978
rect 597828 135922 597884 135978
rect 597456 118294 597512 118350
rect 597580 118294 597636 118350
rect 597704 118294 597760 118350
rect 597828 118294 597884 118350
rect 597456 118170 597512 118226
rect 597580 118170 597636 118226
rect 597704 118170 597760 118226
rect 597828 118170 597884 118226
rect 597456 118046 597512 118102
rect 597580 118046 597636 118102
rect 597704 118046 597760 118102
rect 597828 118046 597884 118102
rect 597456 117922 597512 117978
rect 597580 117922 597636 117978
rect 597704 117922 597760 117978
rect 597828 117922 597884 117978
rect 597456 100294 597512 100350
rect 597580 100294 597636 100350
rect 597704 100294 597760 100350
rect 597828 100294 597884 100350
rect 597456 100170 597512 100226
rect 597580 100170 597636 100226
rect 597704 100170 597760 100226
rect 597828 100170 597884 100226
rect 597456 100046 597512 100102
rect 597580 100046 597636 100102
rect 597704 100046 597760 100102
rect 597828 100046 597884 100102
rect 597456 99922 597512 99978
rect 597580 99922 597636 99978
rect 597704 99922 597760 99978
rect 597828 99922 597884 99978
rect 597456 82294 597512 82350
rect 597580 82294 597636 82350
rect 597704 82294 597760 82350
rect 597828 82294 597884 82350
rect 597456 82170 597512 82226
rect 597580 82170 597636 82226
rect 597704 82170 597760 82226
rect 597828 82170 597884 82226
rect 597456 82046 597512 82102
rect 597580 82046 597636 82102
rect 597704 82046 597760 82102
rect 597828 82046 597884 82102
rect 597456 81922 597512 81978
rect 597580 81922 597636 81978
rect 597704 81922 597760 81978
rect 597828 81922 597884 81978
rect 597456 64294 597512 64350
rect 597580 64294 597636 64350
rect 597704 64294 597760 64350
rect 597828 64294 597884 64350
rect 597456 64170 597512 64226
rect 597580 64170 597636 64226
rect 597704 64170 597760 64226
rect 597828 64170 597884 64226
rect 597456 64046 597512 64102
rect 597580 64046 597636 64102
rect 597704 64046 597760 64102
rect 597828 64046 597884 64102
rect 597456 63922 597512 63978
rect 597580 63922 597636 63978
rect 597704 63922 597760 63978
rect 597828 63922 597884 63978
rect 597456 46294 597512 46350
rect 597580 46294 597636 46350
rect 597704 46294 597760 46350
rect 597828 46294 597884 46350
rect 597456 46170 597512 46226
rect 597580 46170 597636 46226
rect 597704 46170 597760 46226
rect 597828 46170 597884 46226
rect 597456 46046 597512 46102
rect 597580 46046 597636 46102
rect 597704 46046 597760 46102
rect 597828 46046 597884 46102
rect 597456 45922 597512 45978
rect 597580 45922 597636 45978
rect 597704 45922 597760 45978
rect 597828 45922 597884 45978
rect 597456 28294 597512 28350
rect 597580 28294 597636 28350
rect 597704 28294 597760 28350
rect 597828 28294 597884 28350
rect 597456 28170 597512 28226
rect 597580 28170 597636 28226
rect 597704 28170 597760 28226
rect 597828 28170 597884 28226
rect 597456 28046 597512 28102
rect 597580 28046 597636 28102
rect 597704 28046 597760 28102
rect 597828 28046 597884 28102
rect 597456 27922 597512 27978
rect 597580 27922 597636 27978
rect 597704 27922 597760 27978
rect 597828 27922 597884 27978
rect 597456 10294 597512 10350
rect 597580 10294 597636 10350
rect 597704 10294 597760 10350
rect 597828 10294 597884 10350
rect 597456 10170 597512 10226
rect 597580 10170 597636 10226
rect 597704 10170 597760 10226
rect 597828 10170 597884 10226
rect 597456 10046 597512 10102
rect 597580 10046 597636 10102
rect 597704 10046 597760 10102
rect 597828 10046 597884 10102
rect 597456 9922 597512 9978
rect 597580 9922 597636 9978
rect 597704 9922 597760 9978
rect 597828 9922 597884 9978
rect 592914 -1176 592970 -1120
rect 593038 -1176 593094 -1120
rect 593162 -1176 593218 -1120
rect 593286 -1176 593342 -1120
rect 592914 -1300 592970 -1244
rect 593038 -1300 593094 -1244
rect 593162 -1300 593218 -1244
rect 593286 -1300 593342 -1244
rect 592914 -1424 592970 -1368
rect 593038 -1424 593094 -1368
rect 593162 -1424 593218 -1368
rect 593286 -1424 593342 -1368
rect 592914 -1548 592970 -1492
rect 593038 -1548 593094 -1492
rect 593162 -1548 593218 -1492
rect 593286 -1548 593342 -1492
rect 597456 -1176 597512 -1120
rect 597580 -1176 597636 -1120
rect 597704 -1176 597760 -1120
rect 597828 -1176 597884 -1120
rect 597456 -1300 597512 -1244
rect 597580 -1300 597636 -1244
rect 597704 -1300 597760 -1244
rect 597828 -1300 597884 -1244
rect 597456 -1424 597512 -1368
rect 597580 -1424 597636 -1368
rect 597704 -1424 597760 -1368
rect 597828 -1424 597884 -1368
rect 597456 -1548 597512 -1492
rect 597580 -1548 597636 -1492
rect 597704 -1548 597760 -1492
rect 597828 -1548 597884 -1492
<< metal5 >>
rect -1916 598172 597980 598268
rect -1916 598116 -1820 598172
rect -1764 598116 -1696 598172
rect -1640 598116 -1572 598172
rect -1516 598116 -1448 598172
rect -1392 598116 9234 598172
rect 9290 598116 9358 598172
rect 9414 598116 9482 598172
rect 9538 598116 9606 598172
rect 9662 598116 39954 598172
rect 40010 598116 40078 598172
rect 40134 598116 40202 598172
rect 40258 598116 40326 598172
rect 40382 598116 70674 598172
rect 70730 598116 70798 598172
rect 70854 598116 70922 598172
rect 70978 598116 71046 598172
rect 71102 598116 101394 598172
rect 101450 598116 101518 598172
rect 101574 598116 101642 598172
rect 101698 598116 101766 598172
rect 101822 598116 132114 598172
rect 132170 598116 132238 598172
rect 132294 598116 132362 598172
rect 132418 598116 132486 598172
rect 132542 598116 162834 598172
rect 162890 598116 162958 598172
rect 163014 598116 163082 598172
rect 163138 598116 163206 598172
rect 163262 598116 193554 598172
rect 193610 598116 193678 598172
rect 193734 598116 193802 598172
rect 193858 598116 193926 598172
rect 193982 598116 224274 598172
rect 224330 598116 224398 598172
rect 224454 598116 224522 598172
rect 224578 598116 224646 598172
rect 224702 598116 254994 598172
rect 255050 598116 255118 598172
rect 255174 598116 255242 598172
rect 255298 598116 255366 598172
rect 255422 598116 285714 598172
rect 285770 598116 285838 598172
rect 285894 598116 285962 598172
rect 286018 598116 286086 598172
rect 286142 598116 316434 598172
rect 316490 598116 316558 598172
rect 316614 598116 316682 598172
rect 316738 598116 316806 598172
rect 316862 598116 347154 598172
rect 347210 598116 347278 598172
rect 347334 598116 347402 598172
rect 347458 598116 347526 598172
rect 347582 598116 377874 598172
rect 377930 598116 377998 598172
rect 378054 598116 378122 598172
rect 378178 598116 378246 598172
rect 378302 598116 408594 598172
rect 408650 598116 408718 598172
rect 408774 598116 408842 598172
rect 408898 598116 408966 598172
rect 409022 598116 439314 598172
rect 439370 598116 439438 598172
rect 439494 598116 439562 598172
rect 439618 598116 439686 598172
rect 439742 598116 470034 598172
rect 470090 598116 470158 598172
rect 470214 598116 470282 598172
rect 470338 598116 470406 598172
rect 470462 598116 500754 598172
rect 500810 598116 500878 598172
rect 500934 598116 501002 598172
rect 501058 598116 501126 598172
rect 501182 598116 531474 598172
rect 531530 598116 531598 598172
rect 531654 598116 531722 598172
rect 531778 598116 531846 598172
rect 531902 598116 562194 598172
rect 562250 598116 562318 598172
rect 562374 598116 562442 598172
rect 562498 598116 562566 598172
rect 562622 598116 592914 598172
rect 592970 598116 593038 598172
rect 593094 598116 593162 598172
rect 593218 598116 593286 598172
rect 593342 598116 597456 598172
rect 597512 598116 597580 598172
rect 597636 598116 597704 598172
rect 597760 598116 597828 598172
rect 597884 598116 597980 598172
rect -1916 598048 597980 598116
rect -1916 597992 -1820 598048
rect -1764 597992 -1696 598048
rect -1640 597992 -1572 598048
rect -1516 597992 -1448 598048
rect -1392 597992 9234 598048
rect 9290 597992 9358 598048
rect 9414 597992 9482 598048
rect 9538 597992 9606 598048
rect 9662 597992 39954 598048
rect 40010 597992 40078 598048
rect 40134 597992 40202 598048
rect 40258 597992 40326 598048
rect 40382 597992 70674 598048
rect 70730 597992 70798 598048
rect 70854 597992 70922 598048
rect 70978 597992 71046 598048
rect 71102 597992 101394 598048
rect 101450 597992 101518 598048
rect 101574 597992 101642 598048
rect 101698 597992 101766 598048
rect 101822 597992 132114 598048
rect 132170 597992 132238 598048
rect 132294 597992 132362 598048
rect 132418 597992 132486 598048
rect 132542 597992 162834 598048
rect 162890 597992 162958 598048
rect 163014 597992 163082 598048
rect 163138 597992 163206 598048
rect 163262 597992 193554 598048
rect 193610 597992 193678 598048
rect 193734 597992 193802 598048
rect 193858 597992 193926 598048
rect 193982 597992 224274 598048
rect 224330 597992 224398 598048
rect 224454 597992 224522 598048
rect 224578 597992 224646 598048
rect 224702 597992 254994 598048
rect 255050 597992 255118 598048
rect 255174 597992 255242 598048
rect 255298 597992 255366 598048
rect 255422 597992 285714 598048
rect 285770 597992 285838 598048
rect 285894 597992 285962 598048
rect 286018 597992 286086 598048
rect 286142 597992 316434 598048
rect 316490 597992 316558 598048
rect 316614 597992 316682 598048
rect 316738 597992 316806 598048
rect 316862 597992 347154 598048
rect 347210 597992 347278 598048
rect 347334 597992 347402 598048
rect 347458 597992 347526 598048
rect 347582 597992 377874 598048
rect 377930 597992 377998 598048
rect 378054 597992 378122 598048
rect 378178 597992 378246 598048
rect 378302 597992 408594 598048
rect 408650 597992 408718 598048
rect 408774 597992 408842 598048
rect 408898 597992 408966 598048
rect 409022 597992 439314 598048
rect 439370 597992 439438 598048
rect 439494 597992 439562 598048
rect 439618 597992 439686 598048
rect 439742 597992 470034 598048
rect 470090 597992 470158 598048
rect 470214 597992 470282 598048
rect 470338 597992 470406 598048
rect 470462 597992 500754 598048
rect 500810 597992 500878 598048
rect 500934 597992 501002 598048
rect 501058 597992 501126 598048
rect 501182 597992 531474 598048
rect 531530 597992 531598 598048
rect 531654 597992 531722 598048
rect 531778 597992 531846 598048
rect 531902 597992 562194 598048
rect 562250 597992 562318 598048
rect 562374 597992 562442 598048
rect 562498 597992 562566 598048
rect 562622 597992 592914 598048
rect 592970 597992 593038 598048
rect 593094 597992 593162 598048
rect 593218 597992 593286 598048
rect 593342 597992 597456 598048
rect 597512 597992 597580 598048
rect 597636 597992 597704 598048
rect 597760 597992 597828 598048
rect 597884 597992 597980 598048
rect -1916 597924 597980 597992
rect -1916 597868 -1820 597924
rect -1764 597868 -1696 597924
rect -1640 597868 -1572 597924
rect -1516 597868 -1448 597924
rect -1392 597868 9234 597924
rect 9290 597868 9358 597924
rect 9414 597868 9482 597924
rect 9538 597868 9606 597924
rect 9662 597868 39954 597924
rect 40010 597868 40078 597924
rect 40134 597868 40202 597924
rect 40258 597868 40326 597924
rect 40382 597868 70674 597924
rect 70730 597868 70798 597924
rect 70854 597868 70922 597924
rect 70978 597868 71046 597924
rect 71102 597868 101394 597924
rect 101450 597868 101518 597924
rect 101574 597868 101642 597924
rect 101698 597868 101766 597924
rect 101822 597868 132114 597924
rect 132170 597868 132238 597924
rect 132294 597868 132362 597924
rect 132418 597868 132486 597924
rect 132542 597868 162834 597924
rect 162890 597868 162958 597924
rect 163014 597868 163082 597924
rect 163138 597868 163206 597924
rect 163262 597868 193554 597924
rect 193610 597868 193678 597924
rect 193734 597868 193802 597924
rect 193858 597868 193926 597924
rect 193982 597868 224274 597924
rect 224330 597868 224398 597924
rect 224454 597868 224522 597924
rect 224578 597868 224646 597924
rect 224702 597868 254994 597924
rect 255050 597868 255118 597924
rect 255174 597868 255242 597924
rect 255298 597868 255366 597924
rect 255422 597868 285714 597924
rect 285770 597868 285838 597924
rect 285894 597868 285962 597924
rect 286018 597868 286086 597924
rect 286142 597868 316434 597924
rect 316490 597868 316558 597924
rect 316614 597868 316682 597924
rect 316738 597868 316806 597924
rect 316862 597868 347154 597924
rect 347210 597868 347278 597924
rect 347334 597868 347402 597924
rect 347458 597868 347526 597924
rect 347582 597868 377874 597924
rect 377930 597868 377998 597924
rect 378054 597868 378122 597924
rect 378178 597868 378246 597924
rect 378302 597868 408594 597924
rect 408650 597868 408718 597924
rect 408774 597868 408842 597924
rect 408898 597868 408966 597924
rect 409022 597868 439314 597924
rect 439370 597868 439438 597924
rect 439494 597868 439562 597924
rect 439618 597868 439686 597924
rect 439742 597868 470034 597924
rect 470090 597868 470158 597924
rect 470214 597868 470282 597924
rect 470338 597868 470406 597924
rect 470462 597868 500754 597924
rect 500810 597868 500878 597924
rect 500934 597868 501002 597924
rect 501058 597868 501126 597924
rect 501182 597868 531474 597924
rect 531530 597868 531598 597924
rect 531654 597868 531722 597924
rect 531778 597868 531846 597924
rect 531902 597868 562194 597924
rect 562250 597868 562318 597924
rect 562374 597868 562442 597924
rect 562498 597868 562566 597924
rect 562622 597868 592914 597924
rect 592970 597868 593038 597924
rect 593094 597868 593162 597924
rect 593218 597868 593286 597924
rect 593342 597868 597456 597924
rect 597512 597868 597580 597924
rect 597636 597868 597704 597924
rect 597760 597868 597828 597924
rect 597884 597868 597980 597924
rect -1916 597800 597980 597868
rect -1916 597744 -1820 597800
rect -1764 597744 -1696 597800
rect -1640 597744 -1572 597800
rect -1516 597744 -1448 597800
rect -1392 597744 9234 597800
rect 9290 597744 9358 597800
rect 9414 597744 9482 597800
rect 9538 597744 9606 597800
rect 9662 597744 39954 597800
rect 40010 597744 40078 597800
rect 40134 597744 40202 597800
rect 40258 597744 40326 597800
rect 40382 597744 70674 597800
rect 70730 597744 70798 597800
rect 70854 597744 70922 597800
rect 70978 597744 71046 597800
rect 71102 597744 101394 597800
rect 101450 597744 101518 597800
rect 101574 597744 101642 597800
rect 101698 597744 101766 597800
rect 101822 597744 132114 597800
rect 132170 597744 132238 597800
rect 132294 597744 132362 597800
rect 132418 597744 132486 597800
rect 132542 597744 162834 597800
rect 162890 597744 162958 597800
rect 163014 597744 163082 597800
rect 163138 597744 163206 597800
rect 163262 597744 193554 597800
rect 193610 597744 193678 597800
rect 193734 597744 193802 597800
rect 193858 597744 193926 597800
rect 193982 597744 224274 597800
rect 224330 597744 224398 597800
rect 224454 597744 224522 597800
rect 224578 597744 224646 597800
rect 224702 597744 254994 597800
rect 255050 597744 255118 597800
rect 255174 597744 255242 597800
rect 255298 597744 255366 597800
rect 255422 597744 285714 597800
rect 285770 597744 285838 597800
rect 285894 597744 285962 597800
rect 286018 597744 286086 597800
rect 286142 597744 316434 597800
rect 316490 597744 316558 597800
rect 316614 597744 316682 597800
rect 316738 597744 316806 597800
rect 316862 597744 347154 597800
rect 347210 597744 347278 597800
rect 347334 597744 347402 597800
rect 347458 597744 347526 597800
rect 347582 597744 377874 597800
rect 377930 597744 377998 597800
rect 378054 597744 378122 597800
rect 378178 597744 378246 597800
rect 378302 597744 408594 597800
rect 408650 597744 408718 597800
rect 408774 597744 408842 597800
rect 408898 597744 408966 597800
rect 409022 597744 439314 597800
rect 439370 597744 439438 597800
rect 439494 597744 439562 597800
rect 439618 597744 439686 597800
rect 439742 597744 470034 597800
rect 470090 597744 470158 597800
rect 470214 597744 470282 597800
rect 470338 597744 470406 597800
rect 470462 597744 500754 597800
rect 500810 597744 500878 597800
rect 500934 597744 501002 597800
rect 501058 597744 501126 597800
rect 501182 597744 531474 597800
rect 531530 597744 531598 597800
rect 531654 597744 531722 597800
rect 531778 597744 531846 597800
rect 531902 597744 562194 597800
rect 562250 597744 562318 597800
rect 562374 597744 562442 597800
rect 562498 597744 562566 597800
rect 562622 597744 592914 597800
rect 592970 597744 593038 597800
rect 593094 597744 593162 597800
rect 593218 597744 593286 597800
rect 593342 597744 597456 597800
rect 597512 597744 597580 597800
rect 597636 597744 597704 597800
rect 597760 597744 597828 597800
rect 597884 597744 597980 597800
rect -1916 597648 597980 597744
rect -956 597212 597020 597308
rect -956 597156 -860 597212
rect -804 597156 -736 597212
rect -680 597156 -612 597212
rect -556 597156 -488 597212
rect -432 597156 5514 597212
rect 5570 597156 5638 597212
rect 5694 597156 5762 597212
rect 5818 597156 5886 597212
rect 5942 597156 36234 597212
rect 36290 597156 36358 597212
rect 36414 597156 36482 597212
rect 36538 597156 36606 597212
rect 36662 597156 66954 597212
rect 67010 597156 67078 597212
rect 67134 597156 67202 597212
rect 67258 597156 67326 597212
rect 67382 597156 97674 597212
rect 97730 597156 97798 597212
rect 97854 597156 97922 597212
rect 97978 597156 98046 597212
rect 98102 597156 128394 597212
rect 128450 597156 128518 597212
rect 128574 597156 128642 597212
rect 128698 597156 128766 597212
rect 128822 597156 159114 597212
rect 159170 597156 159238 597212
rect 159294 597156 159362 597212
rect 159418 597156 159486 597212
rect 159542 597156 189834 597212
rect 189890 597156 189958 597212
rect 190014 597156 190082 597212
rect 190138 597156 190206 597212
rect 190262 597156 220554 597212
rect 220610 597156 220678 597212
rect 220734 597156 220802 597212
rect 220858 597156 220926 597212
rect 220982 597156 251274 597212
rect 251330 597156 251398 597212
rect 251454 597156 251522 597212
rect 251578 597156 251646 597212
rect 251702 597156 281994 597212
rect 282050 597156 282118 597212
rect 282174 597156 282242 597212
rect 282298 597156 282366 597212
rect 282422 597156 312714 597212
rect 312770 597156 312838 597212
rect 312894 597156 312962 597212
rect 313018 597156 313086 597212
rect 313142 597156 343434 597212
rect 343490 597156 343558 597212
rect 343614 597156 343682 597212
rect 343738 597156 343806 597212
rect 343862 597156 374154 597212
rect 374210 597156 374278 597212
rect 374334 597156 374402 597212
rect 374458 597156 374526 597212
rect 374582 597156 404874 597212
rect 404930 597156 404998 597212
rect 405054 597156 405122 597212
rect 405178 597156 405246 597212
rect 405302 597156 435594 597212
rect 435650 597156 435718 597212
rect 435774 597156 435842 597212
rect 435898 597156 435966 597212
rect 436022 597156 466314 597212
rect 466370 597156 466438 597212
rect 466494 597156 466562 597212
rect 466618 597156 466686 597212
rect 466742 597156 497034 597212
rect 497090 597156 497158 597212
rect 497214 597156 497282 597212
rect 497338 597156 497406 597212
rect 497462 597156 527754 597212
rect 527810 597156 527878 597212
rect 527934 597156 528002 597212
rect 528058 597156 528126 597212
rect 528182 597156 558474 597212
rect 558530 597156 558598 597212
rect 558654 597156 558722 597212
rect 558778 597156 558846 597212
rect 558902 597156 589194 597212
rect 589250 597156 589318 597212
rect 589374 597156 589442 597212
rect 589498 597156 589566 597212
rect 589622 597156 596496 597212
rect 596552 597156 596620 597212
rect 596676 597156 596744 597212
rect 596800 597156 596868 597212
rect 596924 597156 597020 597212
rect -956 597088 597020 597156
rect -956 597032 -860 597088
rect -804 597032 -736 597088
rect -680 597032 -612 597088
rect -556 597032 -488 597088
rect -432 597032 5514 597088
rect 5570 597032 5638 597088
rect 5694 597032 5762 597088
rect 5818 597032 5886 597088
rect 5942 597032 36234 597088
rect 36290 597032 36358 597088
rect 36414 597032 36482 597088
rect 36538 597032 36606 597088
rect 36662 597032 66954 597088
rect 67010 597032 67078 597088
rect 67134 597032 67202 597088
rect 67258 597032 67326 597088
rect 67382 597032 97674 597088
rect 97730 597032 97798 597088
rect 97854 597032 97922 597088
rect 97978 597032 98046 597088
rect 98102 597032 128394 597088
rect 128450 597032 128518 597088
rect 128574 597032 128642 597088
rect 128698 597032 128766 597088
rect 128822 597032 159114 597088
rect 159170 597032 159238 597088
rect 159294 597032 159362 597088
rect 159418 597032 159486 597088
rect 159542 597032 189834 597088
rect 189890 597032 189958 597088
rect 190014 597032 190082 597088
rect 190138 597032 190206 597088
rect 190262 597032 220554 597088
rect 220610 597032 220678 597088
rect 220734 597032 220802 597088
rect 220858 597032 220926 597088
rect 220982 597032 251274 597088
rect 251330 597032 251398 597088
rect 251454 597032 251522 597088
rect 251578 597032 251646 597088
rect 251702 597032 281994 597088
rect 282050 597032 282118 597088
rect 282174 597032 282242 597088
rect 282298 597032 282366 597088
rect 282422 597032 312714 597088
rect 312770 597032 312838 597088
rect 312894 597032 312962 597088
rect 313018 597032 313086 597088
rect 313142 597032 343434 597088
rect 343490 597032 343558 597088
rect 343614 597032 343682 597088
rect 343738 597032 343806 597088
rect 343862 597032 374154 597088
rect 374210 597032 374278 597088
rect 374334 597032 374402 597088
rect 374458 597032 374526 597088
rect 374582 597032 404874 597088
rect 404930 597032 404998 597088
rect 405054 597032 405122 597088
rect 405178 597032 405246 597088
rect 405302 597032 435594 597088
rect 435650 597032 435718 597088
rect 435774 597032 435842 597088
rect 435898 597032 435966 597088
rect 436022 597032 466314 597088
rect 466370 597032 466438 597088
rect 466494 597032 466562 597088
rect 466618 597032 466686 597088
rect 466742 597032 497034 597088
rect 497090 597032 497158 597088
rect 497214 597032 497282 597088
rect 497338 597032 497406 597088
rect 497462 597032 527754 597088
rect 527810 597032 527878 597088
rect 527934 597032 528002 597088
rect 528058 597032 528126 597088
rect 528182 597032 558474 597088
rect 558530 597032 558598 597088
rect 558654 597032 558722 597088
rect 558778 597032 558846 597088
rect 558902 597032 589194 597088
rect 589250 597032 589318 597088
rect 589374 597032 589442 597088
rect 589498 597032 589566 597088
rect 589622 597032 596496 597088
rect 596552 597032 596620 597088
rect 596676 597032 596744 597088
rect 596800 597032 596868 597088
rect 596924 597032 597020 597088
rect -956 596964 597020 597032
rect -956 596908 -860 596964
rect -804 596908 -736 596964
rect -680 596908 -612 596964
rect -556 596908 -488 596964
rect -432 596908 5514 596964
rect 5570 596908 5638 596964
rect 5694 596908 5762 596964
rect 5818 596908 5886 596964
rect 5942 596908 36234 596964
rect 36290 596908 36358 596964
rect 36414 596908 36482 596964
rect 36538 596908 36606 596964
rect 36662 596908 66954 596964
rect 67010 596908 67078 596964
rect 67134 596908 67202 596964
rect 67258 596908 67326 596964
rect 67382 596908 97674 596964
rect 97730 596908 97798 596964
rect 97854 596908 97922 596964
rect 97978 596908 98046 596964
rect 98102 596908 128394 596964
rect 128450 596908 128518 596964
rect 128574 596908 128642 596964
rect 128698 596908 128766 596964
rect 128822 596908 159114 596964
rect 159170 596908 159238 596964
rect 159294 596908 159362 596964
rect 159418 596908 159486 596964
rect 159542 596908 189834 596964
rect 189890 596908 189958 596964
rect 190014 596908 190082 596964
rect 190138 596908 190206 596964
rect 190262 596908 220554 596964
rect 220610 596908 220678 596964
rect 220734 596908 220802 596964
rect 220858 596908 220926 596964
rect 220982 596908 251274 596964
rect 251330 596908 251398 596964
rect 251454 596908 251522 596964
rect 251578 596908 251646 596964
rect 251702 596908 281994 596964
rect 282050 596908 282118 596964
rect 282174 596908 282242 596964
rect 282298 596908 282366 596964
rect 282422 596908 312714 596964
rect 312770 596908 312838 596964
rect 312894 596908 312962 596964
rect 313018 596908 313086 596964
rect 313142 596908 343434 596964
rect 343490 596908 343558 596964
rect 343614 596908 343682 596964
rect 343738 596908 343806 596964
rect 343862 596908 374154 596964
rect 374210 596908 374278 596964
rect 374334 596908 374402 596964
rect 374458 596908 374526 596964
rect 374582 596908 404874 596964
rect 404930 596908 404998 596964
rect 405054 596908 405122 596964
rect 405178 596908 405246 596964
rect 405302 596908 435594 596964
rect 435650 596908 435718 596964
rect 435774 596908 435842 596964
rect 435898 596908 435966 596964
rect 436022 596908 466314 596964
rect 466370 596908 466438 596964
rect 466494 596908 466562 596964
rect 466618 596908 466686 596964
rect 466742 596908 497034 596964
rect 497090 596908 497158 596964
rect 497214 596908 497282 596964
rect 497338 596908 497406 596964
rect 497462 596908 527754 596964
rect 527810 596908 527878 596964
rect 527934 596908 528002 596964
rect 528058 596908 528126 596964
rect 528182 596908 558474 596964
rect 558530 596908 558598 596964
rect 558654 596908 558722 596964
rect 558778 596908 558846 596964
rect 558902 596908 589194 596964
rect 589250 596908 589318 596964
rect 589374 596908 589442 596964
rect 589498 596908 589566 596964
rect 589622 596908 596496 596964
rect 596552 596908 596620 596964
rect 596676 596908 596744 596964
rect 596800 596908 596868 596964
rect 596924 596908 597020 596964
rect -956 596840 597020 596908
rect -956 596784 -860 596840
rect -804 596784 -736 596840
rect -680 596784 -612 596840
rect -556 596784 -488 596840
rect -432 596784 5514 596840
rect 5570 596784 5638 596840
rect 5694 596784 5762 596840
rect 5818 596784 5886 596840
rect 5942 596784 36234 596840
rect 36290 596784 36358 596840
rect 36414 596784 36482 596840
rect 36538 596784 36606 596840
rect 36662 596784 66954 596840
rect 67010 596784 67078 596840
rect 67134 596784 67202 596840
rect 67258 596784 67326 596840
rect 67382 596784 97674 596840
rect 97730 596784 97798 596840
rect 97854 596784 97922 596840
rect 97978 596784 98046 596840
rect 98102 596784 128394 596840
rect 128450 596784 128518 596840
rect 128574 596784 128642 596840
rect 128698 596784 128766 596840
rect 128822 596784 159114 596840
rect 159170 596784 159238 596840
rect 159294 596784 159362 596840
rect 159418 596784 159486 596840
rect 159542 596784 189834 596840
rect 189890 596784 189958 596840
rect 190014 596784 190082 596840
rect 190138 596784 190206 596840
rect 190262 596784 220554 596840
rect 220610 596784 220678 596840
rect 220734 596784 220802 596840
rect 220858 596784 220926 596840
rect 220982 596784 251274 596840
rect 251330 596784 251398 596840
rect 251454 596784 251522 596840
rect 251578 596784 251646 596840
rect 251702 596784 281994 596840
rect 282050 596784 282118 596840
rect 282174 596784 282242 596840
rect 282298 596784 282366 596840
rect 282422 596784 312714 596840
rect 312770 596784 312838 596840
rect 312894 596784 312962 596840
rect 313018 596784 313086 596840
rect 313142 596784 343434 596840
rect 343490 596784 343558 596840
rect 343614 596784 343682 596840
rect 343738 596784 343806 596840
rect 343862 596784 374154 596840
rect 374210 596784 374278 596840
rect 374334 596784 374402 596840
rect 374458 596784 374526 596840
rect 374582 596784 404874 596840
rect 404930 596784 404998 596840
rect 405054 596784 405122 596840
rect 405178 596784 405246 596840
rect 405302 596784 435594 596840
rect 435650 596784 435718 596840
rect 435774 596784 435842 596840
rect 435898 596784 435966 596840
rect 436022 596784 466314 596840
rect 466370 596784 466438 596840
rect 466494 596784 466562 596840
rect 466618 596784 466686 596840
rect 466742 596784 497034 596840
rect 497090 596784 497158 596840
rect 497214 596784 497282 596840
rect 497338 596784 497406 596840
rect 497462 596784 527754 596840
rect 527810 596784 527878 596840
rect 527934 596784 528002 596840
rect 528058 596784 528126 596840
rect 528182 596784 558474 596840
rect 558530 596784 558598 596840
rect 558654 596784 558722 596840
rect 558778 596784 558846 596840
rect 558902 596784 589194 596840
rect 589250 596784 589318 596840
rect 589374 596784 589442 596840
rect 589498 596784 589566 596840
rect 589622 596784 596496 596840
rect 596552 596784 596620 596840
rect 596676 596784 596744 596840
rect 596800 596784 596868 596840
rect 596924 596784 597020 596840
rect -956 596688 597020 596784
rect -1916 586350 597980 586446
rect -1916 586294 -1820 586350
rect -1764 586294 -1696 586350
rect -1640 586294 -1572 586350
rect -1516 586294 -1448 586350
rect -1392 586294 9234 586350
rect 9290 586294 9358 586350
rect 9414 586294 9482 586350
rect 9538 586294 9606 586350
rect 9662 586294 39954 586350
rect 40010 586294 40078 586350
rect 40134 586294 40202 586350
rect 40258 586294 40326 586350
rect 40382 586294 70674 586350
rect 70730 586294 70798 586350
rect 70854 586294 70922 586350
rect 70978 586294 71046 586350
rect 71102 586294 101394 586350
rect 101450 586294 101518 586350
rect 101574 586294 101642 586350
rect 101698 586294 101766 586350
rect 101822 586294 132114 586350
rect 132170 586294 132238 586350
rect 132294 586294 132362 586350
rect 132418 586294 132486 586350
rect 132542 586294 162834 586350
rect 162890 586294 162958 586350
rect 163014 586294 163082 586350
rect 163138 586294 163206 586350
rect 163262 586294 193554 586350
rect 193610 586294 193678 586350
rect 193734 586294 193802 586350
rect 193858 586294 193926 586350
rect 193982 586294 224274 586350
rect 224330 586294 224398 586350
rect 224454 586294 224522 586350
rect 224578 586294 224646 586350
rect 224702 586294 254994 586350
rect 255050 586294 255118 586350
rect 255174 586294 255242 586350
rect 255298 586294 255366 586350
rect 255422 586294 285714 586350
rect 285770 586294 285838 586350
rect 285894 586294 285962 586350
rect 286018 586294 286086 586350
rect 286142 586294 316434 586350
rect 316490 586294 316558 586350
rect 316614 586294 316682 586350
rect 316738 586294 316806 586350
rect 316862 586294 347154 586350
rect 347210 586294 347278 586350
rect 347334 586294 347402 586350
rect 347458 586294 347526 586350
rect 347582 586294 377874 586350
rect 377930 586294 377998 586350
rect 378054 586294 378122 586350
rect 378178 586294 378246 586350
rect 378302 586294 408594 586350
rect 408650 586294 408718 586350
rect 408774 586294 408842 586350
rect 408898 586294 408966 586350
rect 409022 586294 439314 586350
rect 439370 586294 439438 586350
rect 439494 586294 439562 586350
rect 439618 586294 439686 586350
rect 439742 586294 470034 586350
rect 470090 586294 470158 586350
rect 470214 586294 470282 586350
rect 470338 586294 470406 586350
rect 470462 586294 500754 586350
rect 500810 586294 500878 586350
rect 500934 586294 501002 586350
rect 501058 586294 501126 586350
rect 501182 586294 531474 586350
rect 531530 586294 531598 586350
rect 531654 586294 531722 586350
rect 531778 586294 531846 586350
rect 531902 586294 562194 586350
rect 562250 586294 562318 586350
rect 562374 586294 562442 586350
rect 562498 586294 562566 586350
rect 562622 586294 592914 586350
rect 592970 586294 593038 586350
rect 593094 586294 593162 586350
rect 593218 586294 593286 586350
rect 593342 586294 597456 586350
rect 597512 586294 597580 586350
rect 597636 586294 597704 586350
rect 597760 586294 597828 586350
rect 597884 586294 597980 586350
rect -1916 586226 597980 586294
rect -1916 586170 -1820 586226
rect -1764 586170 -1696 586226
rect -1640 586170 -1572 586226
rect -1516 586170 -1448 586226
rect -1392 586170 9234 586226
rect 9290 586170 9358 586226
rect 9414 586170 9482 586226
rect 9538 586170 9606 586226
rect 9662 586170 39954 586226
rect 40010 586170 40078 586226
rect 40134 586170 40202 586226
rect 40258 586170 40326 586226
rect 40382 586170 70674 586226
rect 70730 586170 70798 586226
rect 70854 586170 70922 586226
rect 70978 586170 71046 586226
rect 71102 586170 101394 586226
rect 101450 586170 101518 586226
rect 101574 586170 101642 586226
rect 101698 586170 101766 586226
rect 101822 586170 132114 586226
rect 132170 586170 132238 586226
rect 132294 586170 132362 586226
rect 132418 586170 132486 586226
rect 132542 586170 162834 586226
rect 162890 586170 162958 586226
rect 163014 586170 163082 586226
rect 163138 586170 163206 586226
rect 163262 586170 193554 586226
rect 193610 586170 193678 586226
rect 193734 586170 193802 586226
rect 193858 586170 193926 586226
rect 193982 586170 224274 586226
rect 224330 586170 224398 586226
rect 224454 586170 224522 586226
rect 224578 586170 224646 586226
rect 224702 586170 254994 586226
rect 255050 586170 255118 586226
rect 255174 586170 255242 586226
rect 255298 586170 255366 586226
rect 255422 586170 285714 586226
rect 285770 586170 285838 586226
rect 285894 586170 285962 586226
rect 286018 586170 286086 586226
rect 286142 586170 316434 586226
rect 316490 586170 316558 586226
rect 316614 586170 316682 586226
rect 316738 586170 316806 586226
rect 316862 586170 347154 586226
rect 347210 586170 347278 586226
rect 347334 586170 347402 586226
rect 347458 586170 347526 586226
rect 347582 586170 377874 586226
rect 377930 586170 377998 586226
rect 378054 586170 378122 586226
rect 378178 586170 378246 586226
rect 378302 586170 408594 586226
rect 408650 586170 408718 586226
rect 408774 586170 408842 586226
rect 408898 586170 408966 586226
rect 409022 586170 439314 586226
rect 439370 586170 439438 586226
rect 439494 586170 439562 586226
rect 439618 586170 439686 586226
rect 439742 586170 470034 586226
rect 470090 586170 470158 586226
rect 470214 586170 470282 586226
rect 470338 586170 470406 586226
rect 470462 586170 500754 586226
rect 500810 586170 500878 586226
rect 500934 586170 501002 586226
rect 501058 586170 501126 586226
rect 501182 586170 531474 586226
rect 531530 586170 531598 586226
rect 531654 586170 531722 586226
rect 531778 586170 531846 586226
rect 531902 586170 562194 586226
rect 562250 586170 562318 586226
rect 562374 586170 562442 586226
rect 562498 586170 562566 586226
rect 562622 586170 592914 586226
rect 592970 586170 593038 586226
rect 593094 586170 593162 586226
rect 593218 586170 593286 586226
rect 593342 586170 597456 586226
rect 597512 586170 597580 586226
rect 597636 586170 597704 586226
rect 597760 586170 597828 586226
rect 597884 586170 597980 586226
rect -1916 586102 597980 586170
rect -1916 586046 -1820 586102
rect -1764 586046 -1696 586102
rect -1640 586046 -1572 586102
rect -1516 586046 -1448 586102
rect -1392 586046 9234 586102
rect 9290 586046 9358 586102
rect 9414 586046 9482 586102
rect 9538 586046 9606 586102
rect 9662 586046 39954 586102
rect 40010 586046 40078 586102
rect 40134 586046 40202 586102
rect 40258 586046 40326 586102
rect 40382 586046 70674 586102
rect 70730 586046 70798 586102
rect 70854 586046 70922 586102
rect 70978 586046 71046 586102
rect 71102 586046 101394 586102
rect 101450 586046 101518 586102
rect 101574 586046 101642 586102
rect 101698 586046 101766 586102
rect 101822 586046 132114 586102
rect 132170 586046 132238 586102
rect 132294 586046 132362 586102
rect 132418 586046 132486 586102
rect 132542 586046 162834 586102
rect 162890 586046 162958 586102
rect 163014 586046 163082 586102
rect 163138 586046 163206 586102
rect 163262 586046 193554 586102
rect 193610 586046 193678 586102
rect 193734 586046 193802 586102
rect 193858 586046 193926 586102
rect 193982 586046 224274 586102
rect 224330 586046 224398 586102
rect 224454 586046 224522 586102
rect 224578 586046 224646 586102
rect 224702 586046 254994 586102
rect 255050 586046 255118 586102
rect 255174 586046 255242 586102
rect 255298 586046 255366 586102
rect 255422 586046 285714 586102
rect 285770 586046 285838 586102
rect 285894 586046 285962 586102
rect 286018 586046 286086 586102
rect 286142 586046 316434 586102
rect 316490 586046 316558 586102
rect 316614 586046 316682 586102
rect 316738 586046 316806 586102
rect 316862 586046 347154 586102
rect 347210 586046 347278 586102
rect 347334 586046 347402 586102
rect 347458 586046 347526 586102
rect 347582 586046 377874 586102
rect 377930 586046 377998 586102
rect 378054 586046 378122 586102
rect 378178 586046 378246 586102
rect 378302 586046 408594 586102
rect 408650 586046 408718 586102
rect 408774 586046 408842 586102
rect 408898 586046 408966 586102
rect 409022 586046 439314 586102
rect 439370 586046 439438 586102
rect 439494 586046 439562 586102
rect 439618 586046 439686 586102
rect 439742 586046 470034 586102
rect 470090 586046 470158 586102
rect 470214 586046 470282 586102
rect 470338 586046 470406 586102
rect 470462 586046 500754 586102
rect 500810 586046 500878 586102
rect 500934 586046 501002 586102
rect 501058 586046 501126 586102
rect 501182 586046 531474 586102
rect 531530 586046 531598 586102
rect 531654 586046 531722 586102
rect 531778 586046 531846 586102
rect 531902 586046 562194 586102
rect 562250 586046 562318 586102
rect 562374 586046 562442 586102
rect 562498 586046 562566 586102
rect 562622 586046 592914 586102
rect 592970 586046 593038 586102
rect 593094 586046 593162 586102
rect 593218 586046 593286 586102
rect 593342 586046 597456 586102
rect 597512 586046 597580 586102
rect 597636 586046 597704 586102
rect 597760 586046 597828 586102
rect 597884 586046 597980 586102
rect -1916 585978 597980 586046
rect -1916 585922 -1820 585978
rect -1764 585922 -1696 585978
rect -1640 585922 -1572 585978
rect -1516 585922 -1448 585978
rect -1392 585922 9234 585978
rect 9290 585922 9358 585978
rect 9414 585922 9482 585978
rect 9538 585922 9606 585978
rect 9662 585922 39954 585978
rect 40010 585922 40078 585978
rect 40134 585922 40202 585978
rect 40258 585922 40326 585978
rect 40382 585922 70674 585978
rect 70730 585922 70798 585978
rect 70854 585922 70922 585978
rect 70978 585922 71046 585978
rect 71102 585922 101394 585978
rect 101450 585922 101518 585978
rect 101574 585922 101642 585978
rect 101698 585922 101766 585978
rect 101822 585922 132114 585978
rect 132170 585922 132238 585978
rect 132294 585922 132362 585978
rect 132418 585922 132486 585978
rect 132542 585922 162834 585978
rect 162890 585922 162958 585978
rect 163014 585922 163082 585978
rect 163138 585922 163206 585978
rect 163262 585922 193554 585978
rect 193610 585922 193678 585978
rect 193734 585922 193802 585978
rect 193858 585922 193926 585978
rect 193982 585922 224274 585978
rect 224330 585922 224398 585978
rect 224454 585922 224522 585978
rect 224578 585922 224646 585978
rect 224702 585922 254994 585978
rect 255050 585922 255118 585978
rect 255174 585922 255242 585978
rect 255298 585922 255366 585978
rect 255422 585922 285714 585978
rect 285770 585922 285838 585978
rect 285894 585922 285962 585978
rect 286018 585922 286086 585978
rect 286142 585922 316434 585978
rect 316490 585922 316558 585978
rect 316614 585922 316682 585978
rect 316738 585922 316806 585978
rect 316862 585922 347154 585978
rect 347210 585922 347278 585978
rect 347334 585922 347402 585978
rect 347458 585922 347526 585978
rect 347582 585922 377874 585978
rect 377930 585922 377998 585978
rect 378054 585922 378122 585978
rect 378178 585922 378246 585978
rect 378302 585922 408594 585978
rect 408650 585922 408718 585978
rect 408774 585922 408842 585978
rect 408898 585922 408966 585978
rect 409022 585922 439314 585978
rect 439370 585922 439438 585978
rect 439494 585922 439562 585978
rect 439618 585922 439686 585978
rect 439742 585922 470034 585978
rect 470090 585922 470158 585978
rect 470214 585922 470282 585978
rect 470338 585922 470406 585978
rect 470462 585922 500754 585978
rect 500810 585922 500878 585978
rect 500934 585922 501002 585978
rect 501058 585922 501126 585978
rect 501182 585922 531474 585978
rect 531530 585922 531598 585978
rect 531654 585922 531722 585978
rect 531778 585922 531846 585978
rect 531902 585922 562194 585978
rect 562250 585922 562318 585978
rect 562374 585922 562442 585978
rect 562498 585922 562566 585978
rect 562622 585922 592914 585978
rect 592970 585922 593038 585978
rect 593094 585922 593162 585978
rect 593218 585922 593286 585978
rect 593342 585922 597456 585978
rect 597512 585922 597580 585978
rect 597636 585922 597704 585978
rect 597760 585922 597828 585978
rect 597884 585922 597980 585978
rect -1916 585826 597980 585922
rect -1916 580350 597980 580446
rect -1916 580294 -860 580350
rect -804 580294 -736 580350
rect -680 580294 -612 580350
rect -556 580294 -488 580350
rect -432 580294 5514 580350
rect 5570 580294 5638 580350
rect 5694 580294 5762 580350
rect 5818 580294 5886 580350
rect 5942 580294 36234 580350
rect 36290 580294 36358 580350
rect 36414 580294 36482 580350
rect 36538 580294 36606 580350
rect 36662 580294 66954 580350
rect 67010 580294 67078 580350
rect 67134 580294 67202 580350
rect 67258 580294 67326 580350
rect 67382 580294 97674 580350
rect 97730 580294 97798 580350
rect 97854 580294 97922 580350
rect 97978 580294 98046 580350
rect 98102 580294 128394 580350
rect 128450 580294 128518 580350
rect 128574 580294 128642 580350
rect 128698 580294 128766 580350
rect 128822 580294 159114 580350
rect 159170 580294 159238 580350
rect 159294 580294 159362 580350
rect 159418 580294 159486 580350
rect 159542 580294 189834 580350
rect 189890 580294 189958 580350
rect 190014 580294 190082 580350
rect 190138 580294 190206 580350
rect 190262 580294 220554 580350
rect 220610 580294 220678 580350
rect 220734 580294 220802 580350
rect 220858 580294 220926 580350
rect 220982 580294 251274 580350
rect 251330 580294 251398 580350
rect 251454 580294 251522 580350
rect 251578 580294 251646 580350
rect 251702 580294 281994 580350
rect 282050 580294 282118 580350
rect 282174 580294 282242 580350
rect 282298 580294 282366 580350
rect 282422 580294 312714 580350
rect 312770 580294 312838 580350
rect 312894 580294 312962 580350
rect 313018 580294 313086 580350
rect 313142 580294 343434 580350
rect 343490 580294 343558 580350
rect 343614 580294 343682 580350
rect 343738 580294 343806 580350
rect 343862 580294 374154 580350
rect 374210 580294 374278 580350
rect 374334 580294 374402 580350
rect 374458 580294 374526 580350
rect 374582 580294 404874 580350
rect 404930 580294 404998 580350
rect 405054 580294 405122 580350
rect 405178 580294 405246 580350
rect 405302 580294 435594 580350
rect 435650 580294 435718 580350
rect 435774 580294 435842 580350
rect 435898 580294 435966 580350
rect 436022 580294 466314 580350
rect 466370 580294 466438 580350
rect 466494 580294 466562 580350
rect 466618 580294 466686 580350
rect 466742 580294 497034 580350
rect 497090 580294 497158 580350
rect 497214 580294 497282 580350
rect 497338 580294 497406 580350
rect 497462 580294 527754 580350
rect 527810 580294 527878 580350
rect 527934 580294 528002 580350
rect 528058 580294 528126 580350
rect 528182 580294 558474 580350
rect 558530 580294 558598 580350
rect 558654 580294 558722 580350
rect 558778 580294 558846 580350
rect 558902 580294 589194 580350
rect 589250 580294 589318 580350
rect 589374 580294 589442 580350
rect 589498 580294 589566 580350
rect 589622 580294 596496 580350
rect 596552 580294 596620 580350
rect 596676 580294 596744 580350
rect 596800 580294 596868 580350
rect 596924 580294 597980 580350
rect -1916 580226 597980 580294
rect -1916 580170 -860 580226
rect -804 580170 -736 580226
rect -680 580170 -612 580226
rect -556 580170 -488 580226
rect -432 580170 5514 580226
rect 5570 580170 5638 580226
rect 5694 580170 5762 580226
rect 5818 580170 5886 580226
rect 5942 580170 36234 580226
rect 36290 580170 36358 580226
rect 36414 580170 36482 580226
rect 36538 580170 36606 580226
rect 36662 580170 66954 580226
rect 67010 580170 67078 580226
rect 67134 580170 67202 580226
rect 67258 580170 67326 580226
rect 67382 580170 97674 580226
rect 97730 580170 97798 580226
rect 97854 580170 97922 580226
rect 97978 580170 98046 580226
rect 98102 580170 128394 580226
rect 128450 580170 128518 580226
rect 128574 580170 128642 580226
rect 128698 580170 128766 580226
rect 128822 580170 159114 580226
rect 159170 580170 159238 580226
rect 159294 580170 159362 580226
rect 159418 580170 159486 580226
rect 159542 580170 189834 580226
rect 189890 580170 189958 580226
rect 190014 580170 190082 580226
rect 190138 580170 190206 580226
rect 190262 580170 220554 580226
rect 220610 580170 220678 580226
rect 220734 580170 220802 580226
rect 220858 580170 220926 580226
rect 220982 580170 251274 580226
rect 251330 580170 251398 580226
rect 251454 580170 251522 580226
rect 251578 580170 251646 580226
rect 251702 580170 281994 580226
rect 282050 580170 282118 580226
rect 282174 580170 282242 580226
rect 282298 580170 282366 580226
rect 282422 580170 312714 580226
rect 312770 580170 312838 580226
rect 312894 580170 312962 580226
rect 313018 580170 313086 580226
rect 313142 580170 343434 580226
rect 343490 580170 343558 580226
rect 343614 580170 343682 580226
rect 343738 580170 343806 580226
rect 343862 580170 374154 580226
rect 374210 580170 374278 580226
rect 374334 580170 374402 580226
rect 374458 580170 374526 580226
rect 374582 580170 404874 580226
rect 404930 580170 404998 580226
rect 405054 580170 405122 580226
rect 405178 580170 405246 580226
rect 405302 580170 435594 580226
rect 435650 580170 435718 580226
rect 435774 580170 435842 580226
rect 435898 580170 435966 580226
rect 436022 580170 466314 580226
rect 466370 580170 466438 580226
rect 466494 580170 466562 580226
rect 466618 580170 466686 580226
rect 466742 580170 497034 580226
rect 497090 580170 497158 580226
rect 497214 580170 497282 580226
rect 497338 580170 497406 580226
rect 497462 580170 527754 580226
rect 527810 580170 527878 580226
rect 527934 580170 528002 580226
rect 528058 580170 528126 580226
rect 528182 580170 558474 580226
rect 558530 580170 558598 580226
rect 558654 580170 558722 580226
rect 558778 580170 558846 580226
rect 558902 580170 589194 580226
rect 589250 580170 589318 580226
rect 589374 580170 589442 580226
rect 589498 580170 589566 580226
rect 589622 580170 596496 580226
rect 596552 580170 596620 580226
rect 596676 580170 596744 580226
rect 596800 580170 596868 580226
rect 596924 580170 597980 580226
rect -1916 580102 597980 580170
rect -1916 580046 -860 580102
rect -804 580046 -736 580102
rect -680 580046 -612 580102
rect -556 580046 -488 580102
rect -432 580046 5514 580102
rect 5570 580046 5638 580102
rect 5694 580046 5762 580102
rect 5818 580046 5886 580102
rect 5942 580046 36234 580102
rect 36290 580046 36358 580102
rect 36414 580046 36482 580102
rect 36538 580046 36606 580102
rect 36662 580046 66954 580102
rect 67010 580046 67078 580102
rect 67134 580046 67202 580102
rect 67258 580046 67326 580102
rect 67382 580046 97674 580102
rect 97730 580046 97798 580102
rect 97854 580046 97922 580102
rect 97978 580046 98046 580102
rect 98102 580046 128394 580102
rect 128450 580046 128518 580102
rect 128574 580046 128642 580102
rect 128698 580046 128766 580102
rect 128822 580046 159114 580102
rect 159170 580046 159238 580102
rect 159294 580046 159362 580102
rect 159418 580046 159486 580102
rect 159542 580046 189834 580102
rect 189890 580046 189958 580102
rect 190014 580046 190082 580102
rect 190138 580046 190206 580102
rect 190262 580046 220554 580102
rect 220610 580046 220678 580102
rect 220734 580046 220802 580102
rect 220858 580046 220926 580102
rect 220982 580046 251274 580102
rect 251330 580046 251398 580102
rect 251454 580046 251522 580102
rect 251578 580046 251646 580102
rect 251702 580046 281994 580102
rect 282050 580046 282118 580102
rect 282174 580046 282242 580102
rect 282298 580046 282366 580102
rect 282422 580046 312714 580102
rect 312770 580046 312838 580102
rect 312894 580046 312962 580102
rect 313018 580046 313086 580102
rect 313142 580046 343434 580102
rect 343490 580046 343558 580102
rect 343614 580046 343682 580102
rect 343738 580046 343806 580102
rect 343862 580046 374154 580102
rect 374210 580046 374278 580102
rect 374334 580046 374402 580102
rect 374458 580046 374526 580102
rect 374582 580046 404874 580102
rect 404930 580046 404998 580102
rect 405054 580046 405122 580102
rect 405178 580046 405246 580102
rect 405302 580046 435594 580102
rect 435650 580046 435718 580102
rect 435774 580046 435842 580102
rect 435898 580046 435966 580102
rect 436022 580046 466314 580102
rect 466370 580046 466438 580102
rect 466494 580046 466562 580102
rect 466618 580046 466686 580102
rect 466742 580046 497034 580102
rect 497090 580046 497158 580102
rect 497214 580046 497282 580102
rect 497338 580046 497406 580102
rect 497462 580046 527754 580102
rect 527810 580046 527878 580102
rect 527934 580046 528002 580102
rect 528058 580046 528126 580102
rect 528182 580046 558474 580102
rect 558530 580046 558598 580102
rect 558654 580046 558722 580102
rect 558778 580046 558846 580102
rect 558902 580046 589194 580102
rect 589250 580046 589318 580102
rect 589374 580046 589442 580102
rect 589498 580046 589566 580102
rect 589622 580046 596496 580102
rect 596552 580046 596620 580102
rect 596676 580046 596744 580102
rect 596800 580046 596868 580102
rect 596924 580046 597980 580102
rect -1916 579978 597980 580046
rect -1916 579922 -860 579978
rect -804 579922 -736 579978
rect -680 579922 -612 579978
rect -556 579922 -488 579978
rect -432 579922 5514 579978
rect 5570 579922 5638 579978
rect 5694 579922 5762 579978
rect 5818 579922 5886 579978
rect 5942 579922 36234 579978
rect 36290 579922 36358 579978
rect 36414 579922 36482 579978
rect 36538 579922 36606 579978
rect 36662 579922 66954 579978
rect 67010 579922 67078 579978
rect 67134 579922 67202 579978
rect 67258 579922 67326 579978
rect 67382 579922 97674 579978
rect 97730 579922 97798 579978
rect 97854 579922 97922 579978
rect 97978 579922 98046 579978
rect 98102 579922 128394 579978
rect 128450 579922 128518 579978
rect 128574 579922 128642 579978
rect 128698 579922 128766 579978
rect 128822 579922 159114 579978
rect 159170 579922 159238 579978
rect 159294 579922 159362 579978
rect 159418 579922 159486 579978
rect 159542 579922 189834 579978
rect 189890 579922 189958 579978
rect 190014 579922 190082 579978
rect 190138 579922 190206 579978
rect 190262 579922 220554 579978
rect 220610 579922 220678 579978
rect 220734 579922 220802 579978
rect 220858 579922 220926 579978
rect 220982 579922 251274 579978
rect 251330 579922 251398 579978
rect 251454 579922 251522 579978
rect 251578 579922 251646 579978
rect 251702 579922 281994 579978
rect 282050 579922 282118 579978
rect 282174 579922 282242 579978
rect 282298 579922 282366 579978
rect 282422 579922 312714 579978
rect 312770 579922 312838 579978
rect 312894 579922 312962 579978
rect 313018 579922 313086 579978
rect 313142 579922 343434 579978
rect 343490 579922 343558 579978
rect 343614 579922 343682 579978
rect 343738 579922 343806 579978
rect 343862 579922 374154 579978
rect 374210 579922 374278 579978
rect 374334 579922 374402 579978
rect 374458 579922 374526 579978
rect 374582 579922 404874 579978
rect 404930 579922 404998 579978
rect 405054 579922 405122 579978
rect 405178 579922 405246 579978
rect 405302 579922 435594 579978
rect 435650 579922 435718 579978
rect 435774 579922 435842 579978
rect 435898 579922 435966 579978
rect 436022 579922 466314 579978
rect 466370 579922 466438 579978
rect 466494 579922 466562 579978
rect 466618 579922 466686 579978
rect 466742 579922 497034 579978
rect 497090 579922 497158 579978
rect 497214 579922 497282 579978
rect 497338 579922 497406 579978
rect 497462 579922 527754 579978
rect 527810 579922 527878 579978
rect 527934 579922 528002 579978
rect 528058 579922 528126 579978
rect 528182 579922 558474 579978
rect 558530 579922 558598 579978
rect 558654 579922 558722 579978
rect 558778 579922 558846 579978
rect 558902 579922 589194 579978
rect 589250 579922 589318 579978
rect 589374 579922 589442 579978
rect 589498 579922 589566 579978
rect 589622 579922 596496 579978
rect 596552 579922 596620 579978
rect 596676 579922 596744 579978
rect 596800 579922 596868 579978
rect 596924 579922 597980 579978
rect -1916 579826 597980 579922
rect 200828 571258 330836 571274
rect 200828 571202 200844 571258
rect 200900 571202 330764 571258
rect 330820 571202 330836 571258
rect 200828 571186 330836 571202
rect 290428 569638 333524 569654
rect 290428 569582 290444 569638
rect 290500 569582 333452 569638
rect 333508 569582 333524 569638
rect 290428 569566 333524 569582
rect -1916 568407 597980 568446
rect -1916 568351 39954 568407
rect 40010 568351 40078 568407
rect 40134 568351 40202 568407
rect 40258 568351 40326 568407
rect 40382 568351 101394 568407
rect 101450 568351 101518 568407
rect 101574 568351 101642 568407
rect 101698 568351 101766 568407
rect 101822 568351 597980 568407
rect -1916 568350 597980 568351
rect -1916 568294 -1820 568350
rect -1764 568294 -1696 568350
rect -1640 568294 -1572 568350
rect -1516 568294 -1448 568350
rect -1392 568294 9234 568350
rect 9290 568294 9358 568350
rect 9414 568294 9482 568350
rect 9538 568294 9606 568350
rect 9662 568294 70674 568350
rect 70730 568294 70798 568350
rect 70854 568294 70922 568350
rect 70978 568294 71046 568350
rect 71102 568294 132114 568350
rect 132170 568294 132238 568350
rect 132294 568294 132362 568350
rect 132418 568294 132486 568350
rect 132542 568294 162834 568350
rect 162890 568294 162958 568350
rect 163014 568294 163082 568350
rect 163138 568294 163206 568350
rect 163262 568294 193554 568350
rect 193610 568294 193678 568350
rect 193734 568294 193802 568350
rect 193858 568294 193926 568350
rect 193982 568294 224274 568350
rect 224330 568294 224398 568350
rect 224454 568294 224522 568350
rect 224578 568294 224646 568350
rect 224702 568294 254994 568350
rect 255050 568294 255118 568350
rect 255174 568294 255242 568350
rect 255298 568294 255366 568350
rect 255422 568294 285714 568350
rect 285770 568294 285838 568350
rect 285894 568294 285962 568350
rect 286018 568294 286086 568350
rect 286142 568294 316434 568350
rect 316490 568294 316558 568350
rect 316614 568294 316682 568350
rect 316738 568294 316806 568350
rect 316862 568294 347154 568350
rect 347210 568294 347278 568350
rect 347334 568294 347402 568350
rect 347458 568294 347526 568350
rect 347582 568294 377874 568350
rect 377930 568294 377998 568350
rect 378054 568294 378122 568350
rect 378178 568294 378246 568350
rect 378302 568294 408594 568350
rect 408650 568294 408718 568350
rect 408774 568294 408842 568350
rect 408898 568294 408966 568350
rect 409022 568294 439314 568350
rect 439370 568294 439438 568350
rect 439494 568294 439562 568350
rect 439618 568294 439686 568350
rect 439742 568294 470034 568350
rect 470090 568294 470158 568350
rect 470214 568294 470282 568350
rect 470338 568294 470406 568350
rect 470462 568294 500754 568350
rect 500810 568294 500878 568350
rect 500934 568294 501002 568350
rect 501058 568294 501126 568350
rect 501182 568294 531474 568350
rect 531530 568294 531598 568350
rect 531654 568294 531722 568350
rect 531778 568294 531846 568350
rect 531902 568294 562194 568350
rect 562250 568294 562318 568350
rect 562374 568294 562442 568350
rect 562498 568294 562566 568350
rect 562622 568294 592914 568350
rect 592970 568294 593038 568350
rect 593094 568294 593162 568350
rect 593218 568294 593286 568350
rect 593342 568294 597456 568350
rect 597512 568294 597580 568350
rect 597636 568294 597704 568350
rect 597760 568294 597828 568350
rect 597884 568294 597980 568350
rect -1916 568283 597980 568294
rect -1916 568227 39954 568283
rect 40010 568227 40078 568283
rect 40134 568227 40202 568283
rect 40258 568227 40326 568283
rect 40382 568227 101394 568283
rect 101450 568227 101518 568283
rect 101574 568227 101642 568283
rect 101698 568227 101766 568283
rect 101822 568227 597980 568283
rect -1916 568226 597980 568227
rect -1916 568170 -1820 568226
rect -1764 568170 -1696 568226
rect -1640 568170 -1572 568226
rect -1516 568170 -1448 568226
rect -1392 568170 9234 568226
rect 9290 568170 9358 568226
rect 9414 568170 9482 568226
rect 9538 568170 9606 568226
rect 9662 568170 70674 568226
rect 70730 568170 70798 568226
rect 70854 568170 70922 568226
rect 70978 568170 71046 568226
rect 71102 568170 132114 568226
rect 132170 568170 132238 568226
rect 132294 568170 132362 568226
rect 132418 568170 132486 568226
rect 132542 568170 162834 568226
rect 162890 568170 162958 568226
rect 163014 568170 163082 568226
rect 163138 568170 163206 568226
rect 163262 568170 193554 568226
rect 193610 568170 193678 568226
rect 193734 568170 193802 568226
rect 193858 568170 193926 568226
rect 193982 568170 224274 568226
rect 224330 568170 224398 568226
rect 224454 568170 224522 568226
rect 224578 568170 224646 568226
rect 224702 568170 254994 568226
rect 255050 568170 255118 568226
rect 255174 568170 255242 568226
rect 255298 568170 255366 568226
rect 255422 568170 285714 568226
rect 285770 568170 285838 568226
rect 285894 568170 285962 568226
rect 286018 568170 286086 568226
rect 286142 568170 316434 568226
rect 316490 568170 316558 568226
rect 316614 568170 316682 568226
rect 316738 568170 316806 568226
rect 316862 568170 347154 568226
rect 347210 568170 347278 568226
rect 347334 568170 347402 568226
rect 347458 568170 347526 568226
rect 347582 568170 377874 568226
rect 377930 568170 377998 568226
rect 378054 568170 378122 568226
rect 378178 568170 378246 568226
rect 378302 568170 408594 568226
rect 408650 568170 408718 568226
rect 408774 568170 408842 568226
rect 408898 568170 408966 568226
rect 409022 568170 439314 568226
rect 439370 568170 439438 568226
rect 439494 568170 439562 568226
rect 439618 568170 439686 568226
rect 439742 568170 470034 568226
rect 470090 568170 470158 568226
rect 470214 568170 470282 568226
rect 470338 568170 470406 568226
rect 470462 568170 500754 568226
rect 500810 568170 500878 568226
rect 500934 568170 501002 568226
rect 501058 568170 501126 568226
rect 501182 568170 531474 568226
rect 531530 568170 531598 568226
rect 531654 568170 531722 568226
rect 531778 568170 531846 568226
rect 531902 568170 562194 568226
rect 562250 568170 562318 568226
rect 562374 568170 562442 568226
rect 562498 568170 562566 568226
rect 562622 568170 592914 568226
rect 592970 568170 593038 568226
rect 593094 568170 593162 568226
rect 593218 568170 593286 568226
rect 593342 568170 597456 568226
rect 597512 568170 597580 568226
rect 597636 568170 597704 568226
rect 597760 568170 597828 568226
rect 597884 568170 597980 568226
rect -1916 568102 597980 568170
rect -1916 568046 -1820 568102
rect -1764 568046 -1696 568102
rect -1640 568046 -1572 568102
rect -1516 568046 -1448 568102
rect -1392 568046 9234 568102
rect 9290 568046 9358 568102
rect 9414 568046 9482 568102
rect 9538 568046 9606 568102
rect 9662 568046 70674 568102
rect 70730 568046 70798 568102
rect 70854 568046 70922 568102
rect 70978 568046 71046 568102
rect 71102 568046 132114 568102
rect 132170 568046 132238 568102
rect 132294 568046 132362 568102
rect 132418 568046 132486 568102
rect 132542 568046 162834 568102
rect 162890 568046 162958 568102
rect 163014 568046 163082 568102
rect 163138 568046 163206 568102
rect 163262 568046 193554 568102
rect 193610 568046 193678 568102
rect 193734 568046 193802 568102
rect 193858 568046 193926 568102
rect 193982 568046 224274 568102
rect 224330 568046 224398 568102
rect 224454 568046 224522 568102
rect 224578 568046 224646 568102
rect 224702 568046 254994 568102
rect 255050 568046 255118 568102
rect 255174 568046 255242 568102
rect 255298 568046 255366 568102
rect 255422 568046 285714 568102
rect 285770 568046 285838 568102
rect 285894 568046 285962 568102
rect 286018 568046 286086 568102
rect 286142 568046 316434 568102
rect 316490 568046 316558 568102
rect 316614 568046 316682 568102
rect 316738 568046 316806 568102
rect 316862 568046 347154 568102
rect 347210 568046 347278 568102
rect 347334 568046 347402 568102
rect 347458 568046 347526 568102
rect 347582 568046 377874 568102
rect 377930 568046 377998 568102
rect 378054 568046 378122 568102
rect 378178 568046 378246 568102
rect 378302 568046 408594 568102
rect 408650 568046 408718 568102
rect 408774 568046 408842 568102
rect 408898 568046 408966 568102
rect 409022 568046 439314 568102
rect 439370 568046 439438 568102
rect 439494 568046 439562 568102
rect 439618 568046 439686 568102
rect 439742 568046 470034 568102
rect 470090 568046 470158 568102
rect 470214 568046 470282 568102
rect 470338 568046 470406 568102
rect 470462 568046 500754 568102
rect 500810 568046 500878 568102
rect 500934 568046 501002 568102
rect 501058 568046 501126 568102
rect 501182 568046 531474 568102
rect 531530 568046 531598 568102
rect 531654 568046 531722 568102
rect 531778 568046 531846 568102
rect 531902 568046 562194 568102
rect 562250 568046 562318 568102
rect 562374 568046 562442 568102
rect 562498 568046 562566 568102
rect 562622 568046 592914 568102
rect 592970 568046 593038 568102
rect 593094 568046 593162 568102
rect 593218 568046 593286 568102
rect 593342 568046 597456 568102
rect 597512 568046 597580 568102
rect 597636 568046 597704 568102
rect 597760 568046 597828 568102
rect 597884 568046 597980 568102
rect -1916 567978 597980 568046
rect -1916 567922 -1820 567978
rect -1764 567922 -1696 567978
rect -1640 567922 -1572 567978
rect -1516 567922 -1448 567978
rect -1392 567922 9234 567978
rect 9290 567922 9358 567978
rect 9414 567922 9482 567978
rect 9538 567922 9606 567978
rect 9662 567922 70674 567978
rect 70730 567922 70798 567978
rect 70854 567922 70922 567978
rect 70978 567922 71046 567978
rect 71102 567922 132114 567978
rect 132170 567922 132238 567978
rect 132294 567922 132362 567978
rect 132418 567922 132486 567978
rect 132542 567922 162834 567978
rect 162890 567922 162958 567978
rect 163014 567922 163082 567978
rect 163138 567922 163206 567978
rect 163262 567922 193554 567978
rect 193610 567922 193678 567978
rect 193734 567922 193802 567978
rect 193858 567922 193926 567978
rect 193982 567922 224274 567978
rect 224330 567922 224398 567978
rect 224454 567922 224522 567978
rect 224578 567922 224646 567978
rect 224702 567922 254994 567978
rect 255050 567922 255118 567978
rect 255174 567922 255242 567978
rect 255298 567922 255366 567978
rect 255422 567922 285714 567978
rect 285770 567922 285838 567978
rect 285894 567922 285962 567978
rect 286018 567922 286086 567978
rect 286142 567922 316434 567978
rect 316490 567922 316558 567978
rect 316614 567922 316682 567978
rect 316738 567922 316806 567978
rect 316862 567922 347154 567978
rect 347210 567922 347278 567978
rect 347334 567922 347402 567978
rect 347458 567922 347526 567978
rect 347582 567922 377874 567978
rect 377930 567922 377998 567978
rect 378054 567922 378122 567978
rect 378178 567922 378246 567978
rect 378302 567922 408594 567978
rect 408650 567922 408718 567978
rect 408774 567922 408842 567978
rect 408898 567922 408966 567978
rect 409022 567922 439314 567978
rect 439370 567922 439438 567978
rect 439494 567922 439562 567978
rect 439618 567922 439686 567978
rect 439742 567922 470034 567978
rect 470090 567922 470158 567978
rect 470214 567922 470282 567978
rect 470338 567922 470406 567978
rect 470462 567922 500754 567978
rect 500810 567922 500878 567978
rect 500934 567922 501002 567978
rect 501058 567922 501126 567978
rect 501182 567922 531474 567978
rect 531530 567922 531598 567978
rect 531654 567922 531722 567978
rect 531778 567922 531846 567978
rect 531902 567922 562194 567978
rect 562250 567922 562318 567978
rect 562374 567922 562442 567978
rect 562498 567922 562566 567978
rect 562622 567922 592914 567978
rect 592970 567922 593038 567978
rect 593094 567922 593162 567978
rect 593218 567922 593286 567978
rect 593342 567922 597456 567978
rect 597512 567922 597580 567978
rect 597636 567922 597704 567978
rect 597760 567922 597828 567978
rect 597884 567922 597980 567978
rect -1916 567826 597980 567922
rect 289308 566938 585524 566954
rect 289308 566882 289324 566938
rect 289380 566882 585452 566938
rect 585508 566882 585524 566938
rect 289308 566866 585524 566882
rect -1916 562350 597980 562446
rect -1916 562294 -860 562350
rect -804 562294 -736 562350
rect -680 562294 -612 562350
rect -556 562294 -488 562350
rect -432 562294 5514 562350
rect 5570 562294 5638 562350
rect 5694 562294 5762 562350
rect 5818 562294 5886 562350
rect 5942 562294 24518 562350
rect 24574 562294 24642 562350
rect 24698 562294 36234 562350
rect 36290 562294 36358 562350
rect 36414 562294 36482 562350
rect 36538 562294 36606 562350
rect 36662 562294 55238 562350
rect 55294 562294 55362 562350
rect 55418 562294 66954 562350
rect 67010 562294 67078 562350
rect 67134 562294 67202 562350
rect 67258 562294 67326 562350
rect 67382 562294 86518 562350
rect 86574 562294 86642 562350
rect 86698 562294 97674 562350
rect 97730 562294 97798 562350
rect 97854 562294 97922 562350
rect 97978 562294 98046 562350
rect 98102 562294 117238 562350
rect 117294 562294 117362 562350
rect 117418 562294 128394 562350
rect 128450 562294 128518 562350
rect 128574 562294 128642 562350
rect 128698 562294 128766 562350
rect 128822 562294 148518 562350
rect 148574 562294 148642 562350
rect 148698 562294 159114 562350
rect 159170 562294 159238 562350
rect 159294 562294 159362 562350
rect 159418 562294 159486 562350
rect 159542 562294 179238 562350
rect 179294 562294 179362 562350
rect 179418 562294 189834 562350
rect 189890 562294 189958 562350
rect 190014 562294 190082 562350
rect 190138 562294 190206 562350
rect 190262 562294 210518 562350
rect 210574 562294 210642 562350
rect 210698 562294 220554 562350
rect 220610 562294 220678 562350
rect 220734 562294 220802 562350
rect 220858 562294 220926 562350
rect 220982 562294 241238 562350
rect 241294 562294 241362 562350
rect 241418 562294 251274 562350
rect 251330 562294 251398 562350
rect 251454 562294 251522 562350
rect 251578 562294 251646 562350
rect 251702 562294 272518 562350
rect 272574 562294 272642 562350
rect 272698 562294 303238 562350
rect 303294 562294 303362 562350
rect 303418 562294 343434 562350
rect 343490 562294 343558 562350
rect 343614 562294 343682 562350
rect 343738 562294 343806 562350
rect 343862 562294 356518 562350
rect 356574 562294 356642 562350
rect 356698 562294 374154 562350
rect 374210 562294 374278 562350
rect 374334 562294 374402 562350
rect 374458 562294 374526 562350
rect 374582 562294 387238 562350
rect 387294 562294 387362 562350
rect 387418 562294 404874 562350
rect 404930 562294 404998 562350
rect 405054 562294 405122 562350
rect 405178 562294 405246 562350
rect 405302 562294 418518 562350
rect 418574 562294 418642 562350
rect 418698 562294 435594 562350
rect 435650 562294 435718 562350
rect 435774 562294 435842 562350
rect 435898 562294 435966 562350
rect 436022 562294 449238 562350
rect 449294 562294 449362 562350
rect 449418 562294 466314 562350
rect 466370 562294 466438 562350
rect 466494 562294 466562 562350
rect 466618 562294 466686 562350
rect 466742 562294 480518 562350
rect 480574 562294 480642 562350
rect 480698 562294 497034 562350
rect 497090 562294 497158 562350
rect 497214 562294 497282 562350
rect 497338 562294 497406 562350
rect 497462 562294 511238 562350
rect 511294 562294 511362 562350
rect 511418 562294 527754 562350
rect 527810 562294 527878 562350
rect 527934 562294 528002 562350
rect 528058 562294 528126 562350
rect 528182 562294 542518 562350
rect 542574 562294 542642 562350
rect 542698 562294 558474 562350
rect 558530 562294 558598 562350
rect 558654 562294 558722 562350
rect 558778 562294 558846 562350
rect 558902 562294 573238 562350
rect 573294 562294 573362 562350
rect 573418 562294 589194 562350
rect 589250 562294 589318 562350
rect 589374 562294 589442 562350
rect 589498 562294 589566 562350
rect 589622 562294 596496 562350
rect 596552 562294 596620 562350
rect 596676 562294 596744 562350
rect 596800 562294 596868 562350
rect 596924 562294 597980 562350
rect -1916 562226 597980 562294
rect -1916 562170 -860 562226
rect -804 562170 -736 562226
rect -680 562170 -612 562226
rect -556 562170 -488 562226
rect -432 562170 5514 562226
rect 5570 562170 5638 562226
rect 5694 562170 5762 562226
rect 5818 562170 5886 562226
rect 5942 562170 24518 562226
rect 24574 562170 24642 562226
rect 24698 562170 36234 562226
rect 36290 562170 36358 562226
rect 36414 562170 36482 562226
rect 36538 562170 36606 562226
rect 36662 562170 55238 562226
rect 55294 562170 55362 562226
rect 55418 562170 66954 562226
rect 67010 562170 67078 562226
rect 67134 562170 67202 562226
rect 67258 562170 67326 562226
rect 67382 562170 86518 562226
rect 86574 562170 86642 562226
rect 86698 562170 97674 562226
rect 97730 562170 97798 562226
rect 97854 562170 97922 562226
rect 97978 562170 98046 562226
rect 98102 562170 117238 562226
rect 117294 562170 117362 562226
rect 117418 562170 128394 562226
rect 128450 562170 128518 562226
rect 128574 562170 128642 562226
rect 128698 562170 128766 562226
rect 128822 562170 148518 562226
rect 148574 562170 148642 562226
rect 148698 562170 159114 562226
rect 159170 562170 159238 562226
rect 159294 562170 159362 562226
rect 159418 562170 159486 562226
rect 159542 562170 179238 562226
rect 179294 562170 179362 562226
rect 179418 562170 189834 562226
rect 189890 562170 189958 562226
rect 190014 562170 190082 562226
rect 190138 562170 190206 562226
rect 190262 562170 210518 562226
rect 210574 562170 210642 562226
rect 210698 562170 220554 562226
rect 220610 562170 220678 562226
rect 220734 562170 220802 562226
rect 220858 562170 220926 562226
rect 220982 562170 241238 562226
rect 241294 562170 241362 562226
rect 241418 562170 251274 562226
rect 251330 562170 251398 562226
rect 251454 562170 251522 562226
rect 251578 562170 251646 562226
rect 251702 562170 272518 562226
rect 272574 562170 272642 562226
rect 272698 562170 303238 562226
rect 303294 562170 303362 562226
rect 303418 562170 343434 562226
rect 343490 562170 343558 562226
rect 343614 562170 343682 562226
rect 343738 562170 343806 562226
rect 343862 562170 356518 562226
rect 356574 562170 356642 562226
rect 356698 562170 374154 562226
rect 374210 562170 374278 562226
rect 374334 562170 374402 562226
rect 374458 562170 374526 562226
rect 374582 562170 387238 562226
rect 387294 562170 387362 562226
rect 387418 562170 404874 562226
rect 404930 562170 404998 562226
rect 405054 562170 405122 562226
rect 405178 562170 405246 562226
rect 405302 562170 418518 562226
rect 418574 562170 418642 562226
rect 418698 562170 435594 562226
rect 435650 562170 435718 562226
rect 435774 562170 435842 562226
rect 435898 562170 435966 562226
rect 436022 562170 449238 562226
rect 449294 562170 449362 562226
rect 449418 562170 466314 562226
rect 466370 562170 466438 562226
rect 466494 562170 466562 562226
rect 466618 562170 466686 562226
rect 466742 562170 480518 562226
rect 480574 562170 480642 562226
rect 480698 562170 497034 562226
rect 497090 562170 497158 562226
rect 497214 562170 497282 562226
rect 497338 562170 497406 562226
rect 497462 562170 511238 562226
rect 511294 562170 511362 562226
rect 511418 562170 527754 562226
rect 527810 562170 527878 562226
rect 527934 562170 528002 562226
rect 528058 562170 528126 562226
rect 528182 562170 542518 562226
rect 542574 562170 542642 562226
rect 542698 562170 558474 562226
rect 558530 562170 558598 562226
rect 558654 562170 558722 562226
rect 558778 562170 558846 562226
rect 558902 562170 573238 562226
rect 573294 562170 573362 562226
rect 573418 562170 589194 562226
rect 589250 562170 589318 562226
rect 589374 562170 589442 562226
rect 589498 562170 589566 562226
rect 589622 562170 596496 562226
rect 596552 562170 596620 562226
rect 596676 562170 596744 562226
rect 596800 562170 596868 562226
rect 596924 562170 597980 562226
rect -1916 562102 597980 562170
rect -1916 562046 -860 562102
rect -804 562046 -736 562102
rect -680 562046 -612 562102
rect -556 562046 -488 562102
rect -432 562046 5514 562102
rect 5570 562046 5638 562102
rect 5694 562046 5762 562102
rect 5818 562046 5886 562102
rect 5942 562046 24518 562102
rect 24574 562046 24642 562102
rect 24698 562046 36234 562102
rect 36290 562046 36358 562102
rect 36414 562046 36482 562102
rect 36538 562046 36606 562102
rect 36662 562046 55238 562102
rect 55294 562046 55362 562102
rect 55418 562046 66954 562102
rect 67010 562046 67078 562102
rect 67134 562046 67202 562102
rect 67258 562046 67326 562102
rect 67382 562046 86518 562102
rect 86574 562046 86642 562102
rect 86698 562046 97674 562102
rect 97730 562046 97798 562102
rect 97854 562046 97922 562102
rect 97978 562046 98046 562102
rect 98102 562046 117238 562102
rect 117294 562046 117362 562102
rect 117418 562046 128394 562102
rect 128450 562046 128518 562102
rect 128574 562046 128642 562102
rect 128698 562046 128766 562102
rect 128822 562046 148518 562102
rect 148574 562046 148642 562102
rect 148698 562046 159114 562102
rect 159170 562046 159238 562102
rect 159294 562046 159362 562102
rect 159418 562046 159486 562102
rect 159542 562046 179238 562102
rect 179294 562046 179362 562102
rect 179418 562046 189834 562102
rect 189890 562046 189958 562102
rect 190014 562046 190082 562102
rect 190138 562046 190206 562102
rect 190262 562046 210518 562102
rect 210574 562046 210642 562102
rect 210698 562046 220554 562102
rect 220610 562046 220678 562102
rect 220734 562046 220802 562102
rect 220858 562046 220926 562102
rect 220982 562046 241238 562102
rect 241294 562046 241362 562102
rect 241418 562046 251274 562102
rect 251330 562046 251398 562102
rect 251454 562046 251522 562102
rect 251578 562046 251646 562102
rect 251702 562046 272518 562102
rect 272574 562046 272642 562102
rect 272698 562046 303238 562102
rect 303294 562046 303362 562102
rect 303418 562046 343434 562102
rect 343490 562046 343558 562102
rect 343614 562046 343682 562102
rect 343738 562046 343806 562102
rect 343862 562046 356518 562102
rect 356574 562046 356642 562102
rect 356698 562046 374154 562102
rect 374210 562046 374278 562102
rect 374334 562046 374402 562102
rect 374458 562046 374526 562102
rect 374582 562046 387238 562102
rect 387294 562046 387362 562102
rect 387418 562046 404874 562102
rect 404930 562046 404998 562102
rect 405054 562046 405122 562102
rect 405178 562046 405246 562102
rect 405302 562046 418518 562102
rect 418574 562046 418642 562102
rect 418698 562046 435594 562102
rect 435650 562046 435718 562102
rect 435774 562046 435842 562102
rect 435898 562046 435966 562102
rect 436022 562046 449238 562102
rect 449294 562046 449362 562102
rect 449418 562046 466314 562102
rect 466370 562046 466438 562102
rect 466494 562046 466562 562102
rect 466618 562046 466686 562102
rect 466742 562046 480518 562102
rect 480574 562046 480642 562102
rect 480698 562046 497034 562102
rect 497090 562046 497158 562102
rect 497214 562046 497282 562102
rect 497338 562046 497406 562102
rect 497462 562046 511238 562102
rect 511294 562046 511362 562102
rect 511418 562046 527754 562102
rect 527810 562046 527878 562102
rect 527934 562046 528002 562102
rect 528058 562046 528126 562102
rect 528182 562046 542518 562102
rect 542574 562046 542642 562102
rect 542698 562046 558474 562102
rect 558530 562046 558598 562102
rect 558654 562046 558722 562102
rect 558778 562046 558846 562102
rect 558902 562046 573238 562102
rect 573294 562046 573362 562102
rect 573418 562046 589194 562102
rect 589250 562046 589318 562102
rect 589374 562046 589442 562102
rect 589498 562046 589566 562102
rect 589622 562046 596496 562102
rect 596552 562046 596620 562102
rect 596676 562046 596744 562102
rect 596800 562046 596868 562102
rect 596924 562046 597980 562102
rect -1916 561978 597980 562046
rect -1916 561922 -860 561978
rect -804 561922 -736 561978
rect -680 561922 -612 561978
rect -556 561922 -488 561978
rect -432 561922 5514 561978
rect 5570 561922 5638 561978
rect 5694 561922 5762 561978
rect 5818 561922 5886 561978
rect 5942 561922 24518 561978
rect 24574 561922 24642 561978
rect 24698 561922 36234 561978
rect 36290 561922 36358 561978
rect 36414 561922 36482 561978
rect 36538 561922 36606 561978
rect 36662 561922 55238 561978
rect 55294 561922 55362 561978
rect 55418 561922 66954 561978
rect 67010 561922 67078 561978
rect 67134 561922 67202 561978
rect 67258 561922 67326 561978
rect 67382 561922 86518 561978
rect 86574 561922 86642 561978
rect 86698 561922 97674 561978
rect 97730 561922 97798 561978
rect 97854 561922 97922 561978
rect 97978 561922 98046 561978
rect 98102 561922 117238 561978
rect 117294 561922 117362 561978
rect 117418 561922 128394 561978
rect 128450 561922 128518 561978
rect 128574 561922 128642 561978
rect 128698 561922 128766 561978
rect 128822 561922 148518 561978
rect 148574 561922 148642 561978
rect 148698 561922 159114 561978
rect 159170 561922 159238 561978
rect 159294 561922 159362 561978
rect 159418 561922 159486 561978
rect 159542 561922 179238 561978
rect 179294 561922 179362 561978
rect 179418 561922 189834 561978
rect 189890 561922 189958 561978
rect 190014 561922 190082 561978
rect 190138 561922 190206 561978
rect 190262 561922 210518 561978
rect 210574 561922 210642 561978
rect 210698 561922 220554 561978
rect 220610 561922 220678 561978
rect 220734 561922 220802 561978
rect 220858 561922 220926 561978
rect 220982 561922 241238 561978
rect 241294 561922 241362 561978
rect 241418 561922 251274 561978
rect 251330 561922 251398 561978
rect 251454 561922 251522 561978
rect 251578 561922 251646 561978
rect 251702 561922 272518 561978
rect 272574 561922 272642 561978
rect 272698 561922 303238 561978
rect 303294 561922 303362 561978
rect 303418 561922 343434 561978
rect 343490 561922 343558 561978
rect 343614 561922 343682 561978
rect 343738 561922 343806 561978
rect 343862 561922 356518 561978
rect 356574 561922 356642 561978
rect 356698 561922 374154 561978
rect 374210 561922 374278 561978
rect 374334 561922 374402 561978
rect 374458 561922 374526 561978
rect 374582 561922 387238 561978
rect 387294 561922 387362 561978
rect 387418 561922 404874 561978
rect 404930 561922 404998 561978
rect 405054 561922 405122 561978
rect 405178 561922 405246 561978
rect 405302 561922 418518 561978
rect 418574 561922 418642 561978
rect 418698 561922 435594 561978
rect 435650 561922 435718 561978
rect 435774 561922 435842 561978
rect 435898 561922 435966 561978
rect 436022 561922 449238 561978
rect 449294 561922 449362 561978
rect 449418 561922 466314 561978
rect 466370 561922 466438 561978
rect 466494 561922 466562 561978
rect 466618 561922 466686 561978
rect 466742 561922 480518 561978
rect 480574 561922 480642 561978
rect 480698 561922 497034 561978
rect 497090 561922 497158 561978
rect 497214 561922 497282 561978
rect 497338 561922 497406 561978
rect 497462 561922 511238 561978
rect 511294 561922 511362 561978
rect 511418 561922 527754 561978
rect 527810 561922 527878 561978
rect 527934 561922 528002 561978
rect 528058 561922 528126 561978
rect 528182 561922 542518 561978
rect 542574 561922 542642 561978
rect 542698 561922 558474 561978
rect 558530 561922 558598 561978
rect 558654 561922 558722 561978
rect 558778 561922 558846 561978
rect 558902 561922 573238 561978
rect 573294 561922 573362 561978
rect 573418 561922 589194 561978
rect 589250 561922 589318 561978
rect 589374 561922 589442 561978
rect 589498 561922 589566 561978
rect 589622 561922 596496 561978
rect 596552 561922 596620 561978
rect 596676 561922 596744 561978
rect 596800 561922 596868 561978
rect 596924 561922 597980 561978
rect -1916 561826 597980 561922
rect 144044 555238 201700 555254
rect 144044 555182 144060 555238
rect 144116 555182 201628 555238
rect 201684 555182 201700 555238
rect 144044 555166 201700 555182
rect 352700 555238 473748 555254
rect 352700 555182 352716 555238
rect 352772 555182 414652 555238
rect 414708 555182 473676 555238
rect 473732 555182 473748 555238
rect 352700 555166 473748 555182
rect 476012 554698 478844 554714
rect 476012 554642 476028 554698
rect 476084 554642 478844 554698
rect 476012 554626 478844 554642
rect 478756 554534 478844 554626
rect 18380 554518 141108 554534
rect 18380 554462 18396 554518
rect 18452 554462 82684 554518
rect 82740 554462 141036 554518
rect 141092 554462 141108 554518
rect 18380 554446 141108 554462
rect 478756 554518 519108 554534
rect 478756 554462 519036 554518
rect 519092 554462 519108 554518
rect 478756 554446 519108 554462
rect -1916 550350 597980 550446
rect -1916 550294 -1820 550350
rect -1764 550294 -1696 550350
rect -1640 550294 -1572 550350
rect -1516 550294 -1448 550350
rect -1392 550294 9234 550350
rect 9290 550294 9358 550350
rect 9414 550294 9482 550350
rect 9538 550294 9606 550350
rect 9662 550294 39878 550350
rect 39934 550294 40002 550350
rect 40058 550294 70674 550350
rect 70730 550294 70798 550350
rect 70854 550294 70922 550350
rect 70978 550294 71046 550350
rect 71102 550294 101878 550350
rect 101934 550294 102002 550350
rect 102058 550294 132114 550350
rect 132170 550294 132238 550350
rect 132294 550294 132362 550350
rect 132418 550294 132486 550350
rect 132542 550294 163878 550350
rect 163934 550294 164002 550350
rect 164058 550294 193554 550350
rect 193610 550294 193678 550350
rect 193734 550294 193802 550350
rect 193858 550294 193926 550350
rect 193982 550294 225878 550350
rect 225934 550294 226002 550350
rect 226058 550294 254994 550350
rect 255050 550294 255118 550350
rect 255174 550294 255242 550350
rect 255298 550294 255366 550350
rect 255422 550294 287878 550350
rect 287934 550294 288002 550350
rect 288058 550294 318598 550350
rect 318654 550294 318722 550350
rect 318778 550294 347154 550350
rect 347210 550294 347278 550350
rect 347334 550294 347402 550350
rect 347458 550294 347526 550350
rect 347582 550294 371878 550350
rect 371934 550294 372002 550350
rect 372058 550294 377874 550350
rect 377930 550294 377998 550350
rect 378054 550294 378122 550350
rect 378178 550294 378246 550350
rect 378302 550294 408594 550350
rect 408650 550294 408718 550350
rect 408774 550294 408842 550350
rect 408898 550294 408966 550350
rect 409022 550294 433878 550350
rect 433934 550294 434002 550350
rect 434058 550294 470034 550350
rect 470090 550294 470158 550350
rect 470214 550294 470282 550350
rect 470338 550294 470406 550350
rect 470462 550294 495878 550350
rect 495934 550294 496002 550350
rect 496058 550294 500754 550350
rect 500810 550294 500878 550350
rect 500934 550294 501002 550350
rect 501058 550294 501126 550350
rect 501182 550294 531474 550350
rect 531530 550294 531598 550350
rect 531654 550294 531722 550350
rect 531778 550294 531846 550350
rect 531902 550294 557878 550350
rect 557934 550294 558002 550350
rect 558058 550294 562194 550350
rect 562250 550294 562318 550350
rect 562374 550294 562442 550350
rect 562498 550294 562566 550350
rect 562622 550294 592914 550350
rect 592970 550294 593038 550350
rect 593094 550294 593162 550350
rect 593218 550294 593286 550350
rect 593342 550294 597456 550350
rect 597512 550294 597580 550350
rect 597636 550294 597704 550350
rect 597760 550294 597828 550350
rect 597884 550294 597980 550350
rect -1916 550226 597980 550294
rect -1916 550170 -1820 550226
rect -1764 550170 -1696 550226
rect -1640 550170 -1572 550226
rect -1516 550170 -1448 550226
rect -1392 550170 9234 550226
rect 9290 550170 9358 550226
rect 9414 550170 9482 550226
rect 9538 550170 9606 550226
rect 9662 550170 39878 550226
rect 39934 550170 40002 550226
rect 40058 550170 70674 550226
rect 70730 550170 70798 550226
rect 70854 550170 70922 550226
rect 70978 550170 71046 550226
rect 71102 550170 101878 550226
rect 101934 550170 102002 550226
rect 102058 550170 132114 550226
rect 132170 550170 132238 550226
rect 132294 550170 132362 550226
rect 132418 550170 132486 550226
rect 132542 550170 163878 550226
rect 163934 550170 164002 550226
rect 164058 550170 193554 550226
rect 193610 550170 193678 550226
rect 193734 550170 193802 550226
rect 193858 550170 193926 550226
rect 193982 550170 225878 550226
rect 225934 550170 226002 550226
rect 226058 550170 254994 550226
rect 255050 550170 255118 550226
rect 255174 550170 255242 550226
rect 255298 550170 255366 550226
rect 255422 550170 287878 550226
rect 287934 550170 288002 550226
rect 288058 550170 318598 550226
rect 318654 550170 318722 550226
rect 318778 550170 347154 550226
rect 347210 550170 347278 550226
rect 347334 550170 347402 550226
rect 347458 550170 347526 550226
rect 347582 550170 371878 550226
rect 371934 550170 372002 550226
rect 372058 550170 377874 550226
rect 377930 550170 377998 550226
rect 378054 550170 378122 550226
rect 378178 550170 378246 550226
rect 378302 550170 408594 550226
rect 408650 550170 408718 550226
rect 408774 550170 408842 550226
rect 408898 550170 408966 550226
rect 409022 550170 433878 550226
rect 433934 550170 434002 550226
rect 434058 550170 470034 550226
rect 470090 550170 470158 550226
rect 470214 550170 470282 550226
rect 470338 550170 470406 550226
rect 470462 550170 495878 550226
rect 495934 550170 496002 550226
rect 496058 550170 500754 550226
rect 500810 550170 500878 550226
rect 500934 550170 501002 550226
rect 501058 550170 501126 550226
rect 501182 550170 531474 550226
rect 531530 550170 531598 550226
rect 531654 550170 531722 550226
rect 531778 550170 531846 550226
rect 531902 550170 557878 550226
rect 557934 550170 558002 550226
rect 558058 550170 562194 550226
rect 562250 550170 562318 550226
rect 562374 550170 562442 550226
rect 562498 550170 562566 550226
rect 562622 550170 592914 550226
rect 592970 550170 593038 550226
rect 593094 550170 593162 550226
rect 593218 550170 593286 550226
rect 593342 550170 597456 550226
rect 597512 550170 597580 550226
rect 597636 550170 597704 550226
rect 597760 550170 597828 550226
rect 597884 550170 597980 550226
rect -1916 550102 597980 550170
rect -1916 550046 -1820 550102
rect -1764 550046 -1696 550102
rect -1640 550046 -1572 550102
rect -1516 550046 -1448 550102
rect -1392 550046 9234 550102
rect 9290 550046 9358 550102
rect 9414 550046 9482 550102
rect 9538 550046 9606 550102
rect 9662 550046 39878 550102
rect 39934 550046 40002 550102
rect 40058 550046 70674 550102
rect 70730 550046 70798 550102
rect 70854 550046 70922 550102
rect 70978 550046 71046 550102
rect 71102 550046 101878 550102
rect 101934 550046 102002 550102
rect 102058 550046 132114 550102
rect 132170 550046 132238 550102
rect 132294 550046 132362 550102
rect 132418 550046 132486 550102
rect 132542 550046 163878 550102
rect 163934 550046 164002 550102
rect 164058 550046 193554 550102
rect 193610 550046 193678 550102
rect 193734 550046 193802 550102
rect 193858 550046 193926 550102
rect 193982 550046 225878 550102
rect 225934 550046 226002 550102
rect 226058 550046 254994 550102
rect 255050 550046 255118 550102
rect 255174 550046 255242 550102
rect 255298 550046 255366 550102
rect 255422 550046 287878 550102
rect 287934 550046 288002 550102
rect 288058 550046 318598 550102
rect 318654 550046 318722 550102
rect 318778 550046 347154 550102
rect 347210 550046 347278 550102
rect 347334 550046 347402 550102
rect 347458 550046 347526 550102
rect 347582 550046 371878 550102
rect 371934 550046 372002 550102
rect 372058 550046 377874 550102
rect 377930 550046 377998 550102
rect 378054 550046 378122 550102
rect 378178 550046 378246 550102
rect 378302 550046 408594 550102
rect 408650 550046 408718 550102
rect 408774 550046 408842 550102
rect 408898 550046 408966 550102
rect 409022 550046 433878 550102
rect 433934 550046 434002 550102
rect 434058 550046 470034 550102
rect 470090 550046 470158 550102
rect 470214 550046 470282 550102
rect 470338 550046 470406 550102
rect 470462 550046 495878 550102
rect 495934 550046 496002 550102
rect 496058 550046 500754 550102
rect 500810 550046 500878 550102
rect 500934 550046 501002 550102
rect 501058 550046 501126 550102
rect 501182 550046 531474 550102
rect 531530 550046 531598 550102
rect 531654 550046 531722 550102
rect 531778 550046 531846 550102
rect 531902 550046 557878 550102
rect 557934 550046 558002 550102
rect 558058 550046 562194 550102
rect 562250 550046 562318 550102
rect 562374 550046 562442 550102
rect 562498 550046 562566 550102
rect 562622 550046 592914 550102
rect 592970 550046 593038 550102
rect 593094 550046 593162 550102
rect 593218 550046 593286 550102
rect 593342 550046 597456 550102
rect 597512 550046 597580 550102
rect 597636 550046 597704 550102
rect 597760 550046 597828 550102
rect 597884 550046 597980 550102
rect -1916 549978 597980 550046
rect -1916 549922 -1820 549978
rect -1764 549922 -1696 549978
rect -1640 549922 -1572 549978
rect -1516 549922 -1448 549978
rect -1392 549922 9234 549978
rect 9290 549922 9358 549978
rect 9414 549922 9482 549978
rect 9538 549922 9606 549978
rect 9662 549922 39878 549978
rect 39934 549922 40002 549978
rect 40058 549922 70674 549978
rect 70730 549922 70798 549978
rect 70854 549922 70922 549978
rect 70978 549922 71046 549978
rect 71102 549922 101878 549978
rect 101934 549922 102002 549978
rect 102058 549922 132114 549978
rect 132170 549922 132238 549978
rect 132294 549922 132362 549978
rect 132418 549922 132486 549978
rect 132542 549922 163878 549978
rect 163934 549922 164002 549978
rect 164058 549922 193554 549978
rect 193610 549922 193678 549978
rect 193734 549922 193802 549978
rect 193858 549922 193926 549978
rect 193982 549922 225878 549978
rect 225934 549922 226002 549978
rect 226058 549922 254994 549978
rect 255050 549922 255118 549978
rect 255174 549922 255242 549978
rect 255298 549922 255366 549978
rect 255422 549922 287878 549978
rect 287934 549922 288002 549978
rect 288058 549922 318598 549978
rect 318654 549922 318722 549978
rect 318778 549922 347154 549978
rect 347210 549922 347278 549978
rect 347334 549922 347402 549978
rect 347458 549922 347526 549978
rect 347582 549922 371878 549978
rect 371934 549922 372002 549978
rect 372058 549922 377874 549978
rect 377930 549922 377998 549978
rect 378054 549922 378122 549978
rect 378178 549922 378246 549978
rect 378302 549922 408594 549978
rect 408650 549922 408718 549978
rect 408774 549922 408842 549978
rect 408898 549922 408966 549978
rect 409022 549922 433878 549978
rect 433934 549922 434002 549978
rect 434058 549922 470034 549978
rect 470090 549922 470158 549978
rect 470214 549922 470282 549978
rect 470338 549922 470406 549978
rect 470462 549922 495878 549978
rect 495934 549922 496002 549978
rect 496058 549922 500754 549978
rect 500810 549922 500878 549978
rect 500934 549922 501002 549978
rect 501058 549922 501126 549978
rect 501182 549922 531474 549978
rect 531530 549922 531598 549978
rect 531654 549922 531722 549978
rect 531778 549922 531846 549978
rect 531902 549922 557878 549978
rect 557934 549922 558002 549978
rect 558058 549922 562194 549978
rect 562250 549922 562318 549978
rect 562374 549922 562442 549978
rect 562498 549922 562566 549978
rect 562622 549922 592914 549978
rect 592970 549922 593038 549978
rect 593094 549922 593162 549978
rect 593218 549922 593286 549978
rect 593342 549922 597456 549978
rect 597512 549922 597580 549978
rect 597636 549922 597704 549978
rect 597760 549922 597828 549978
rect 597884 549922 597980 549978
rect -1916 549826 597980 549922
rect -1916 544350 597980 544446
rect -1916 544294 -860 544350
rect -804 544294 -736 544350
rect -680 544294 -612 544350
rect -556 544294 -488 544350
rect -432 544294 5514 544350
rect 5570 544294 5638 544350
rect 5694 544294 5762 544350
rect 5818 544294 5886 544350
rect 5942 544294 24518 544350
rect 24574 544294 24642 544350
rect 24698 544294 36234 544350
rect 36290 544294 36358 544350
rect 36414 544294 36482 544350
rect 36538 544294 36606 544350
rect 36662 544294 55238 544350
rect 55294 544294 55362 544350
rect 55418 544294 66954 544350
rect 67010 544294 67078 544350
rect 67134 544294 67202 544350
rect 67258 544294 67326 544350
rect 67382 544294 86518 544350
rect 86574 544294 86642 544350
rect 86698 544294 97674 544350
rect 97730 544294 97798 544350
rect 97854 544294 97922 544350
rect 97978 544294 98046 544350
rect 98102 544294 117238 544350
rect 117294 544294 117362 544350
rect 117418 544294 128394 544350
rect 128450 544294 128518 544350
rect 128574 544294 128642 544350
rect 128698 544294 128766 544350
rect 128822 544294 148518 544350
rect 148574 544294 148642 544350
rect 148698 544294 159114 544350
rect 159170 544294 159238 544350
rect 159294 544294 159362 544350
rect 159418 544294 159486 544350
rect 159542 544294 179238 544350
rect 179294 544294 179362 544350
rect 179418 544294 189834 544350
rect 189890 544294 189958 544350
rect 190014 544294 190082 544350
rect 190138 544294 190206 544350
rect 190262 544294 210518 544350
rect 210574 544294 210642 544350
rect 210698 544294 220554 544350
rect 220610 544294 220678 544350
rect 220734 544294 220802 544350
rect 220858 544294 220926 544350
rect 220982 544294 241238 544350
rect 241294 544294 241362 544350
rect 241418 544294 251274 544350
rect 251330 544294 251398 544350
rect 251454 544294 251522 544350
rect 251578 544294 251646 544350
rect 251702 544294 272518 544350
rect 272574 544294 272642 544350
rect 272698 544294 303238 544350
rect 303294 544294 303362 544350
rect 303418 544294 343434 544350
rect 343490 544294 343558 544350
rect 343614 544294 343682 544350
rect 343738 544294 343806 544350
rect 343862 544294 356518 544350
rect 356574 544294 356642 544350
rect 356698 544294 374154 544350
rect 374210 544294 374278 544350
rect 374334 544294 374402 544350
rect 374458 544294 374526 544350
rect 374582 544294 387238 544350
rect 387294 544294 387362 544350
rect 387418 544294 404874 544350
rect 404930 544294 404998 544350
rect 405054 544294 405122 544350
rect 405178 544294 405246 544350
rect 405302 544294 418518 544350
rect 418574 544294 418642 544350
rect 418698 544294 449238 544350
rect 449294 544294 449362 544350
rect 449418 544294 466314 544350
rect 466370 544294 466438 544350
rect 466494 544294 466562 544350
rect 466618 544294 466686 544350
rect 466742 544294 480518 544350
rect 480574 544294 480642 544350
rect 480698 544294 497034 544350
rect 497090 544294 497158 544350
rect 497214 544294 497282 544350
rect 497338 544294 497406 544350
rect 497462 544294 511238 544350
rect 511294 544294 511362 544350
rect 511418 544294 527754 544350
rect 527810 544294 527878 544350
rect 527934 544294 528002 544350
rect 528058 544294 528126 544350
rect 528182 544294 542518 544350
rect 542574 544294 542642 544350
rect 542698 544294 558474 544350
rect 558530 544294 558598 544350
rect 558654 544294 558722 544350
rect 558778 544294 558846 544350
rect 558902 544294 573238 544350
rect 573294 544294 573362 544350
rect 573418 544294 589194 544350
rect 589250 544294 589318 544350
rect 589374 544294 589442 544350
rect 589498 544294 589566 544350
rect 589622 544294 596496 544350
rect 596552 544294 596620 544350
rect 596676 544294 596744 544350
rect 596800 544294 596868 544350
rect 596924 544294 597980 544350
rect -1916 544226 597980 544294
rect -1916 544170 -860 544226
rect -804 544170 -736 544226
rect -680 544170 -612 544226
rect -556 544170 -488 544226
rect -432 544170 5514 544226
rect 5570 544170 5638 544226
rect 5694 544170 5762 544226
rect 5818 544170 5886 544226
rect 5942 544170 24518 544226
rect 24574 544170 24642 544226
rect 24698 544170 36234 544226
rect 36290 544170 36358 544226
rect 36414 544170 36482 544226
rect 36538 544170 36606 544226
rect 36662 544170 55238 544226
rect 55294 544170 55362 544226
rect 55418 544170 66954 544226
rect 67010 544170 67078 544226
rect 67134 544170 67202 544226
rect 67258 544170 67326 544226
rect 67382 544170 86518 544226
rect 86574 544170 86642 544226
rect 86698 544170 97674 544226
rect 97730 544170 97798 544226
rect 97854 544170 97922 544226
rect 97978 544170 98046 544226
rect 98102 544170 117238 544226
rect 117294 544170 117362 544226
rect 117418 544170 128394 544226
rect 128450 544170 128518 544226
rect 128574 544170 128642 544226
rect 128698 544170 128766 544226
rect 128822 544170 148518 544226
rect 148574 544170 148642 544226
rect 148698 544170 159114 544226
rect 159170 544170 159238 544226
rect 159294 544170 159362 544226
rect 159418 544170 159486 544226
rect 159542 544170 179238 544226
rect 179294 544170 179362 544226
rect 179418 544170 189834 544226
rect 189890 544170 189958 544226
rect 190014 544170 190082 544226
rect 190138 544170 190206 544226
rect 190262 544170 210518 544226
rect 210574 544170 210642 544226
rect 210698 544170 220554 544226
rect 220610 544170 220678 544226
rect 220734 544170 220802 544226
rect 220858 544170 220926 544226
rect 220982 544170 241238 544226
rect 241294 544170 241362 544226
rect 241418 544170 251274 544226
rect 251330 544170 251398 544226
rect 251454 544170 251522 544226
rect 251578 544170 251646 544226
rect 251702 544170 272518 544226
rect 272574 544170 272642 544226
rect 272698 544170 303238 544226
rect 303294 544170 303362 544226
rect 303418 544170 343434 544226
rect 343490 544170 343558 544226
rect 343614 544170 343682 544226
rect 343738 544170 343806 544226
rect 343862 544170 356518 544226
rect 356574 544170 356642 544226
rect 356698 544170 374154 544226
rect 374210 544170 374278 544226
rect 374334 544170 374402 544226
rect 374458 544170 374526 544226
rect 374582 544170 387238 544226
rect 387294 544170 387362 544226
rect 387418 544170 404874 544226
rect 404930 544170 404998 544226
rect 405054 544170 405122 544226
rect 405178 544170 405246 544226
rect 405302 544170 418518 544226
rect 418574 544170 418642 544226
rect 418698 544170 449238 544226
rect 449294 544170 449362 544226
rect 449418 544170 466314 544226
rect 466370 544170 466438 544226
rect 466494 544170 466562 544226
rect 466618 544170 466686 544226
rect 466742 544170 480518 544226
rect 480574 544170 480642 544226
rect 480698 544170 497034 544226
rect 497090 544170 497158 544226
rect 497214 544170 497282 544226
rect 497338 544170 497406 544226
rect 497462 544170 511238 544226
rect 511294 544170 511362 544226
rect 511418 544170 527754 544226
rect 527810 544170 527878 544226
rect 527934 544170 528002 544226
rect 528058 544170 528126 544226
rect 528182 544170 542518 544226
rect 542574 544170 542642 544226
rect 542698 544170 558474 544226
rect 558530 544170 558598 544226
rect 558654 544170 558722 544226
rect 558778 544170 558846 544226
rect 558902 544170 573238 544226
rect 573294 544170 573362 544226
rect 573418 544170 589194 544226
rect 589250 544170 589318 544226
rect 589374 544170 589442 544226
rect 589498 544170 589566 544226
rect 589622 544170 596496 544226
rect 596552 544170 596620 544226
rect 596676 544170 596744 544226
rect 596800 544170 596868 544226
rect 596924 544170 597980 544226
rect -1916 544102 597980 544170
rect -1916 544046 -860 544102
rect -804 544046 -736 544102
rect -680 544046 -612 544102
rect -556 544046 -488 544102
rect -432 544046 5514 544102
rect 5570 544046 5638 544102
rect 5694 544046 5762 544102
rect 5818 544046 5886 544102
rect 5942 544046 24518 544102
rect 24574 544046 24642 544102
rect 24698 544046 36234 544102
rect 36290 544046 36358 544102
rect 36414 544046 36482 544102
rect 36538 544046 36606 544102
rect 36662 544046 55238 544102
rect 55294 544046 55362 544102
rect 55418 544046 66954 544102
rect 67010 544046 67078 544102
rect 67134 544046 67202 544102
rect 67258 544046 67326 544102
rect 67382 544046 86518 544102
rect 86574 544046 86642 544102
rect 86698 544046 97674 544102
rect 97730 544046 97798 544102
rect 97854 544046 97922 544102
rect 97978 544046 98046 544102
rect 98102 544046 117238 544102
rect 117294 544046 117362 544102
rect 117418 544046 128394 544102
rect 128450 544046 128518 544102
rect 128574 544046 128642 544102
rect 128698 544046 128766 544102
rect 128822 544046 148518 544102
rect 148574 544046 148642 544102
rect 148698 544046 159114 544102
rect 159170 544046 159238 544102
rect 159294 544046 159362 544102
rect 159418 544046 159486 544102
rect 159542 544046 179238 544102
rect 179294 544046 179362 544102
rect 179418 544046 189834 544102
rect 189890 544046 189958 544102
rect 190014 544046 190082 544102
rect 190138 544046 190206 544102
rect 190262 544046 210518 544102
rect 210574 544046 210642 544102
rect 210698 544046 220554 544102
rect 220610 544046 220678 544102
rect 220734 544046 220802 544102
rect 220858 544046 220926 544102
rect 220982 544046 241238 544102
rect 241294 544046 241362 544102
rect 241418 544046 251274 544102
rect 251330 544046 251398 544102
rect 251454 544046 251522 544102
rect 251578 544046 251646 544102
rect 251702 544046 272518 544102
rect 272574 544046 272642 544102
rect 272698 544046 303238 544102
rect 303294 544046 303362 544102
rect 303418 544046 343434 544102
rect 343490 544046 343558 544102
rect 343614 544046 343682 544102
rect 343738 544046 343806 544102
rect 343862 544046 356518 544102
rect 356574 544046 356642 544102
rect 356698 544046 374154 544102
rect 374210 544046 374278 544102
rect 374334 544046 374402 544102
rect 374458 544046 374526 544102
rect 374582 544046 387238 544102
rect 387294 544046 387362 544102
rect 387418 544046 404874 544102
rect 404930 544046 404998 544102
rect 405054 544046 405122 544102
rect 405178 544046 405246 544102
rect 405302 544046 418518 544102
rect 418574 544046 418642 544102
rect 418698 544046 449238 544102
rect 449294 544046 449362 544102
rect 449418 544046 466314 544102
rect 466370 544046 466438 544102
rect 466494 544046 466562 544102
rect 466618 544046 466686 544102
rect 466742 544046 480518 544102
rect 480574 544046 480642 544102
rect 480698 544046 497034 544102
rect 497090 544046 497158 544102
rect 497214 544046 497282 544102
rect 497338 544046 497406 544102
rect 497462 544046 511238 544102
rect 511294 544046 511362 544102
rect 511418 544046 527754 544102
rect 527810 544046 527878 544102
rect 527934 544046 528002 544102
rect 528058 544046 528126 544102
rect 528182 544046 542518 544102
rect 542574 544046 542642 544102
rect 542698 544046 558474 544102
rect 558530 544046 558598 544102
rect 558654 544046 558722 544102
rect 558778 544046 558846 544102
rect 558902 544046 573238 544102
rect 573294 544046 573362 544102
rect 573418 544046 589194 544102
rect 589250 544046 589318 544102
rect 589374 544046 589442 544102
rect 589498 544046 589566 544102
rect 589622 544046 596496 544102
rect 596552 544046 596620 544102
rect 596676 544046 596744 544102
rect 596800 544046 596868 544102
rect 596924 544046 597980 544102
rect -1916 543978 597980 544046
rect -1916 543922 -860 543978
rect -804 543922 -736 543978
rect -680 543922 -612 543978
rect -556 543922 -488 543978
rect -432 543922 5514 543978
rect 5570 543922 5638 543978
rect 5694 543922 5762 543978
rect 5818 543922 5886 543978
rect 5942 543922 24518 543978
rect 24574 543922 24642 543978
rect 24698 543922 36234 543978
rect 36290 543922 36358 543978
rect 36414 543922 36482 543978
rect 36538 543922 36606 543978
rect 36662 543922 55238 543978
rect 55294 543922 55362 543978
rect 55418 543922 66954 543978
rect 67010 543922 67078 543978
rect 67134 543922 67202 543978
rect 67258 543922 67326 543978
rect 67382 543922 86518 543978
rect 86574 543922 86642 543978
rect 86698 543922 97674 543978
rect 97730 543922 97798 543978
rect 97854 543922 97922 543978
rect 97978 543922 98046 543978
rect 98102 543922 117238 543978
rect 117294 543922 117362 543978
rect 117418 543922 128394 543978
rect 128450 543922 128518 543978
rect 128574 543922 128642 543978
rect 128698 543922 128766 543978
rect 128822 543922 148518 543978
rect 148574 543922 148642 543978
rect 148698 543922 159114 543978
rect 159170 543922 159238 543978
rect 159294 543922 159362 543978
rect 159418 543922 159486 543978
rect 159542 543922 179238 543978
rect 179294 543922 179362 543978
rect 179418 543922 189834 543978
rect 189890 543922 189958 543978
rect 190014 543922 190082 543978
rect 190138 543922 190206 543978
rect 190262 543922 210518 543978
rect 210574 543922 210642 543978
rect 210698 543922 220554 543978
rect 220610 543922 220678 543978
rect 220734 543922 220802 543978
rect 220858 543922 220926 543978
rect 220982 543922 241238 543978
rect 241294 543922 241362 543978
rect 241418 543922 251274 543978
rect 251330 543922 251398 543978
rect 251454 543922 251522 543978
rect 251578 543922 251646 543978
rect 251702 543922 272518 543978
rect 272574 543922 272642 543978
rect 272698 543922 303238 543978
rect 303294 543922 303362 543978
rect 303418 543922 343434 543978
rect 343490 543922 343558 543978
rect 343614 543922 343682 543978
rect 343738 543922 343806 543978
rect 343862 543922 356518 543978
rect 356574 543922 356642 543978
rect 356698 543922 374154 543978
rect 374210 543922 374278 543978
rect 374334 543922 374402 543978
rect 374458 543922 374526 543978
rect 374582 543922 387238 543978
rect 387294 543922 387362 543978
rect 387418 543922 404874 543978
rect 404930 543922 404998 543978
rect 405054 543922 405122 543978
rect 405178 543922 405246 543978
rect 405302 543922 418518 543978
rect 418574 543922 418642 543978
rect 418698 543922 449238 543978
rect 449294 543922 449362 543978
rect 449418 543922 466314 543978
rect 466370 543922 466438 543978
rect 466494 543922 466562 543978
rect 466618 543922 466686 543978
rect 466742 543922 480518 543978
rect 480574 543922 480642 543978
rect 480698 543922 497034 543978
rect 497090 543922 497158 543978
rect 497214 543922 497282 543978
rect 497338 543922 497406 543978
rect 497462 543922 511238 543978
rect 511294 543922 511362 543978
rect 511418 543922 527754 543978
rect 527810 543922 527878 543978
rect 527934 543922 528002 543978
rect 528058 543922 528126 543978
rect 528182 543922 542518 543978
rect 542574 543922 542642 543978
rect 542698 543922 558474 543978
rect 558530 543922 558598 543978
rect 558654 543922 558722 543978
rect 558778 543922 558846 543978
rect 558902 543922 573238 543978
rect 573294 543922 573362 543978
rect 573418 543922 589194 543978
rect 589250 543922 589318 543978
rect 589374 543922 589442 543978
rect 589498 543922 589566 543978
rect 589622 543922 596496 543978
rect 596552 543922 596620 543978
rect 596676 543922 596744 543978
rect 596800 543922 596868 543978
rect 596924 543922 597980 543978
rect -1916 543826 597980 543922
rect 204860 533458 263860 533474
rect 204860 533402 204876 533458
rect 204932 533402 263788 533458
rect 263844 533402 263860 533458
rect 204860 533386 263860 533402
rect -1916 532350 597980 532446
rect -1916 532294 -1820 532350
rect -1764 532294 -1696 532350
rect -1640 532294 -1572 532350
rect -1516 532294 -1448 532350
rect -1392 532294 9234 532350
rect 9290 532294 9358 532350
rect 9414 532294 9482 532350
rect 9538 532294 9606 532350
rect 9662 532294 39878 532350
rect 39934 532294 40002 532350
rect 40058 532294 70674 532350
rect 70730 532294 70798 532350
rect 70854 532294 70922 532350
rect 70978 532294 71046 532350
rect 71102 532294 101878 532350
rect 101934 532294 102002 532350
rect 102058 532294 132114 532350
rect 132170 532294 132238 532350
rect 132294 532294 132362 532350
rect 132418 532294 132486 532350
rect 132542 532294 162834 532350
rect 162890 532294 162958 532350
rect 163014 532294 163082 532350
rect 163138 532294 163206 532350
rect 163262 532294 163878 532350
rect 163934 532294 164002 532350
rect 164058 532294 193554 532350
rect 193610 532294 193678 532350
rect 193734 532294 193802 532350
rect 193858 532294 193926 532350
rect 193982 532294 224274 532350
rect 224330 532294 224398 532350
rect 224454 532294 224522 532350
rect 224578 532294 224646 532350
rect 224702 532294 225878 532350
rect 225934 532294 226002 532350
rect 226058 532294 254994 532350
rect 255050 532294 255118 532350
rect 255174 532294 255242 532350
rect 255298 532294 255366 532350
rect 255422 532294 287878 532350
rect 287934 532294 288002 532350
rect 288058 532294 318598 532350
rect 318654 532294 318722 532350
rect 318778 532294 347154 532350
rect 347210 532294 347278 532350
rect 347334 532294 347402 532350
rect 347458 532294 347526 532350
rect 347582 532294 371878 532350
rect 371934 532294 372002 532350
rect 372058 532294 377874 532350
rect 377930 532294 377998 532350
rect 378054 532294 378122 532350
rect 378178 532294 378246 532350
rect 378302 532294 408594 532350
rect 408650 532294 408718 532350
rect 408774 532294 408842 532350
rect 408898 532294 408966 532350
rect 409022 532294 433878 532350
rect 433934 532294 434002 532350
rect 434058 532294 439314 532350
rect 439370 532294 439438 532350
rect 439494 532294 439562 532350
rect 439618 532294 439686 532350
rect 439742 532294 470034 532350
rect 470090 532294 470158 532350
rect 470214 532294 470282 532350
rect 470338 532294 470406 532350
rect 470462 532294 495878 532350
rect 495934 532294 496002 532350
rect 496058 532294 500754 532350
rect 500810 532294 500878 532350
rect 500934 532294 501002 532350
rect 501058 532294 501126 532350
rect 501182 532294 531474 532350
rect 531530 532294 531598 532350
rect 531654 532294 531722 532350
rect 531778 532294 531846 532350
rect 531902 532294 557878 532350
rect 557934 532294 558002 532350
rect 558058 532294 562194 532350
rect 562250 532294 562318 532350
rect 562374 532294 562442 532350
rect 562498 532294 562566 532350
rect 562622 532294 592914 532350
rect 592970 532294 593038 532350
rect 593094 532294 593162 532350
rect 593218 532294 593286 532350
rect 593342 532294 597456 532350
rect 597512 532294 597580 532350
rect 597636 532294 597704 532350
rect 597760 532294 597828 532350
rect 597884 532294 597980 532350
rect -1916 532226 597980 532294
rect -1916 532170 -1820 532226
rect -1764 532170 -1696 532226
rect -1640 532170 -1572 532226
rect -1516 532170 -1448 532226
rect -1392 532170 9234 532226
rect 9290 532170 9358 532226
rect 9414 532170 9482 532226
rect 9538 532170 9606 532226
rect 9662 532170 39878 532226
rect 39934 532170 40002 532226
rect 40058 532170 70674 532226
rect 70730 532170 70798 532226
rect 70854 532170 70922 532226
rect 70978 532170 71046 532226
rect 71102 532170 101878 532226
rect 101934 532170 102002 532226
rect 102058 532170 132114 532226
rect 132170 532170 132238 532226
rect 132294 532170 132362 532226
rect 132418 532170 132486 532226
rect 132542 532170 162834 532226
rect 162890 532170 162958 532226
rect 163014 532170 163082 532226
rect 163138 532170 163206 532226
rect 163262 532170 163878 532226
rect 163934 532170 164002 532226
rect 164058 532170 193554 532226
rect 193610 532170 193678 532226
rect 193734 532170 193802 532226
rect 193858 532170 193926 532226
rect 193982 532170 224274 532226
rect 224330 532170 224398 532226
rect 224454 532170 224522 532226
rect 224578 532170 224646 532226
rect 224702 532170 225878 532226
rect 225934 532170 226002 532226
rect 226058 532170 254994 532226
rect 255050 532170 255118 532226
rect 255174 532170 255242 532226
rect 255298 532170 255366 532226
rect 255422 532170 287878 532226
rect 287934 532170 288002 532226
rect 288058 532170 318598 532226
rect 318654 532170 318722 532226
rect 318778 532170 347154 532226
rect 347210 532170 347278 532226
rect 347334 532170 347402 532226
rect 347458 532170 347526 532226
rect 347582 532170 371878 532226
rect 371934 532170 372002 532226
rect 372058 532170 377874 532226
rect 377930 532170 377998 532226
rect 378054 532170 378122 532226
rect 378178 532170 378246 532226
rect 378302 532170 408594 532226
rect 408650 532170 408718 532226
rect 408774 532170 408842 532226
rect 408898 532170 408966 532226
rect 409022 532170 433878 532226
rect 433934 532170 434002 532226
rect 434058 532170 439314 532226
rect 439370 532170 439438 532226
rect 439494 532170 439562 532226
rect 439618 532170 439686 532226
rect 439742 532170 470034 532226
rect 470090 532170 470158 532226
rect 470214 532170 470282 532226
rect 470338 532170 470406 532226
rect 470462 532170 495878 532226
rect 495934 532170 496002 532226
rect 496058 532170 500754 532226
rect 500810 532170 500878 532226
rect 500934 532170 501002 532226
rect 501058 532170 501126 532226
rect 501182 532170 531474 532226
rect 531530 532170 531598 532226
rect 531654 532170 531722 532226
rect 531778 532170 531846 532226
rect 531902 532170 557878 532226
rect 557934 532170 558002 532226
rect 558058 532170 562194 532226
rect 562250 532170 562318 532226
rect 562374 532170 562442 532226
rect 562498 532170 562566 532226
rect 562622 532170 592914 532226
rect 592970 532170 593038 532226
rect 593094 532170 593162 532226
rect 593218 532170 593286 532226
rect 593342 532170 597456 532226
rect 597512 532170 597580 532226
rect 597636 532170 597704 532226
rect 597760 532170 597828 532226
rect 597884 532170 597980 532226
rect -1916 532102 597980 532170
rect -1916 532046 -1820 532102
rect -1764 532046 -1696 532102
rect -1640 532046 -1572 532102
rect -1516 532046 -1448 532102
rect -1392 532046 9234 532102
rect 9290 532046 9358 532102
rect 9414 532046 9482 532102
rect 9538 532046 9606 532102
rect 9662 532046 39878 532102
rect 39934 532046 40002 532102
rect 40058 532046 70674 532102
rect 70730 532046 70798 532102
rect 70854 532046 70922 532102
rect 70978 532046 71046 532102
rect 71102 532046 101878 532102
rect 101934 532046 102002 532102
rect 102058 532046 132114 532102
rect 132170 532046 132238 532102
rect 132294 532046 132362 532102
rect 132418 532046 132486 532102
rect 132542 532046 162834 532102
rect 162890 532046 162958 532102
rect 163014 532046 163082 532102
rect 163138 532046 163206 532102
rect 163262 532046 163878 532102
rect 163934 532046 164002 532102
rect 164058 532046 193554 532102
rect 193610 532046 193678 532102
rect 193734 532046 193802 532102
rect 193858 532046 193926 532102
rect 193982 532046 224274 532102
rect 224330 532046 224398 532102
rect 224454 532046 224522 532102
rect 224578 532046 224646 532102
rect 224702 532046 225878 532102
rect 225934 532046 226002 532102
rect 226058 532046 254994 532102
rect 255050 532046 255118 532102
rect 255174 532046 255242 532102
rect 255298 532046 255366 532102
rect 255422 532046 287878 532102
rect 287934 532046 288002 532102
rect 288058 532046 318598 532102
rect 318654 532046 318722 532102
rect 318778 532046 347154 532102
rect 347210 532046 347278 532102
rect 347334 532046 347402 532102
rect 347458 532046 347526 532102
rect 347582 532046 371878 532102
rect 371934 532046 372002 532102
rect 372058 532046 377874 532102
rect 377930 532046 377998 532102
rect 378054 532046 378122 532102
rect 378178 532046 378246 532102
rect 378302 532046 408594 532102
rect 408650 532046 408718 532102
rect 408774 532046 408842 532102
rect 408898 532046 408966 532102
rect 409022 532046 433878 532102
rect 433934 532046 434002 532102
rect 434058 532046 439314 532102
rect 439370 532046 439438 532102
rect 439494 532046 439562 532102
rect 439618 532046 439686 532102
rect 439742 532046 470034 532102
rect 470090 532046 470158 532102
rect 470214 532046 470282 532102
rect 470338 532046 470406 532102
rect 470462 532046 495878 532102
rect 495934 532046 496002 532102
rect 496058 532046 500754 532102
rect 500810 532046 500878 532102
rect 500934 532046 501002 532102
rect 501058 532046 501126 532102
rect 501182 532046 531474 532102
rect 531530 532046 531598 532102
rect 531654 532046 531722 532102
rect 531778 532046 531846 532102
rect 531902 532046 557878 532102
rect 557934 532046 558002 532102
rect 558058 532046 562194 532102
rect 562250 532046 562318 532102
rect 562374 532046 562442 532102
rect 562498 532046 562566 532102
rect 562622 532046 592914 532102
rect 592970 532046 593038 532102
rect 593094 532046 593162 532102
rect 593218 532046 593286 532102
rect 593342 532046 597456 532102
rect 597512 532046 597580 532102
rect 597636 532046 597704 532102
rect 597760 532046 597828 532102
rect 597884 532046 597980 532102
rect -1916 531978 597980 532046
rect -1916 531922 -1820 531978
rect -1764 531922 -1696 531978
rect -1640 531922 -1572 531978
rect -1516 531922 -1448 531978
rect -1392 531922 9234 531978
rect 9290 531922 9358 531978
rect 9414 531922 9482 531978
rect 9538 531922 9606 531978
rect 9662 531922 39878 531978
rect 39934 531922 40002 531978
rect 40058 531922 70674 531978
rect 70730 531922 70798 531978
rect 70854 531922 70922 531978
rect 70978 531922 71046 531978
rect 71102 531922 101878 531978
rect 101934 531922 102002 531978
rect 102058 531922 132114 531978
rect 132170 531922 132238 531978
rect 132294 531922 132362 531978
rect 132418 531922 132486 531978
rect 132542 531922 162834 531978
rect 162890 531922 162958 531978
rect 163014 531922 163082 531978
rect 163138 531922 163206 531978
rect 163262 531922 163878 531978
rect 163934 531922 164002 531978
rect 164058 531922 193554 531978
rect 193610 531922 193678 531978
rect 193734 531922 193802 531978
rect 193858 531922 193926 531978
rect 193982 531922 224274 531978
rect 224330 531922 224398 531978
rect 224454 531922 224522 531978
rect 224578 531922 224646 531978
rect 224702 531922 225878 531978
rect 225934 531922 226002 531978
rect 226058 531922 254994 531978
rect 255050 531922 255118 531978
rect 255174 531922 255242 531978
rect 255298 531922 255366 531978
rect 255422 531922 287878 531978
rect 287934 531922 288002 531978
rect 288058 531922 318598 531978
rect 318654 531922 318722 531978
rect 318778 531922 347154 531978
rect 347210 531922 347278 531978
rect 347334 531922 347402 531978
rect 347458 531922 347526 531978
rect 347582 531922 371878 531978
rect 371934 531922 372002 531978
rect 372058 531922 377874 531978
rect 377930 531922 377998 531978
rect 378054 531922 378122 531978
rect 378178 531922 378246 531978
rect 378302 531922 408594 531978
rect 408650 531922 408718 531978
rect 408774 531922 408842 531978
rect 408898 531922 408966 531978
rect 409022 531922 433878 531978
rect 433934 531922 434002 531978
rect 434058 531922 439314 531978
rect 439370 531922 439438 531978
rect 439494 531922 439562 531978
rect 439618 531922 439686 531978
rect 439742 531922 470034 531978
rect 470090 531922 470158 531978
rect 470214 531922 470282 531978
rect 470338 531922 470406 531978
rect 470462 531922 495878 531978
rect 495934 531922 496002 531978
rect 496058 531922 500754 531978
rect 500810 531922 500878 531978
rect 500934 531922 501002 531978
rect 501058 531922 501126 531978
rect 501182 531922 531474 531978
rect 531530 531922 531598 531978
rect 531654 531922 531722 531978
rect 531778 531922 531846 531978
rect 531902 531922 557878 531978
rect 557934 531922 558002 531978
rect 558058 531922 562194 531978
rect 562250 531922 562318 531978
rect 562374 531922 562442 531978
rect 562498 531922 562566 531978
rect 562622 531922 592914 531978
rect 592970 531922 593038 531978
rect 593094 531922 593162 531978
rect 593218 531922 593286 531978
rect 593342 531922 597456 531978
rect 597512 531922 597580 531978
rect 597636 531922 597704 531978
rect 597760 531922 597828 531978
rect 597884 531922 597980 531978
rect -1916 531826 597980 531922
rect -1916 526350 597980 526446
rect -1916 526294 -860 526350
rect -804 526294 -736 526350
rect -680 526294 -612 526350
rect -556 526294 -488 526350
rect -432 526294 5514 526350
rect 5570 526294 5638 526350
rect 5694 526294 5762 526350
rect 5818 526294 5886 526350
rect 5942 526294 36234 526350
rect 36290 526294 36358 526350
rect 36414 526294 36482 526350
rect 36538 526294 36606 526350
rect 36662 526294 66954 526350
rect 67010 526294 67078 526350
rect 67134 526294 67202 526350
rect 67258 526294 67326 526350
rect 67382 526294 97674 526350
rect 97730 526294 97798 526350
rect 97854 526294 97922 526350
rect 97978 526294 98046 526350
rect 98102 526294 128394 526350
rect 128450 526294 128518 526350
rect 128574 526294 128642 526350
rect 128698 526294 128766 526350
rect 128822 526294 159114 526350
rect 159170 526294 159238 526350
rect 159294 526294 159362 526350
rect 159418 526294 159486 526350
rect 159542 526294 189834 526350
rect 189890 526294 189958 526350
rect 190014 526294 190082 526350
rect 190138 526294 190206 526350
rect 190262 526294 220554 526350
rect 220610 526294 220678 526350
rect 220734 526294 220802 526350
rect 220858 526294 220926 526350
rect 220982 526294 251274 526350
rect 251330 526294 251398 526350
rect 251454 526294 251522 526350
rect 251578 526294 251646 526350
rect 251702 526294 272518 526350
rect 272574 526294 272642 526350
rect 272698 526294 303238 526350
rect 303294 526294 303362 526350
rect 303418 526294 343434 526350
rect 343490 526294 343558 526350
rect 343614 526294 343682 526350
rect 343738 526294 343806 526350
rect 343862 526294 374154 526350
rect 374210 526294 374278 526350
rect 374334 526294 374402 526350
rect 374458 526294 374526 526350
rect 374582 526294 404874 526350
rect 404930 526294 404998 526350
rect 405054 526294 405122 526350
rect 405178 526294 405246 526350
rect 405302 526294 435594 526350
rect 435650 526294 435718 526350
rect 435774 526294 435842 526350
rect 435898 526294 435966 526350
rect 436022 526294 466314 526350
rect 466370 526294 466438 526350
rect 466494 526294 466562 526350
rect 466618 526294 466686 526350
rect 466742 526294 497034 526350
rect 497090 526294 497158 526350
rect 497214 526294 497282 526350
rect 497338 526294 497406 526350
rect 497462 526294 527754 526350
rect 527810 526294 527878 526350
rect 527934 526294 528002 526350
rect 528058 526294 528126 526350
rect 528182 526294 558474 526350
rect 558530 526294 558598 526350
rect 558654 526294 558722 526350
rect 558778 526294 558846 526350
rect 558902 526294 589194 526350
rect 589250 526294 589318 526350
rect 589374 526294 589442 526350
rect 589498 526294 589566 526350
rect 589622 526294 596496 526350
rect 596552 526294 596620 526350
rect 596676 526294 596744 526350
rect 596800 526294 596868 526350
rect 596924 526294 597980 526350
rect -1916 526226 597980 526294
rect -1916 526170 -860 526226
rect -804 526170 -736 526226
rect -680 526170 -612 526226
rect -556 526170 -488 526226
rect -432 526170 5514 526226
rect 5570 526170 5638 526226
rect 5694 526170 5762 526226
rect 5818 526170 5886 526226
rect 5942 526170 36234 526226
rect 36290 526170 36358 526226
rect 36414 526170 36482 526226
rect 36538 526170 36606 526226
rect 36662 526170 66954 526226
rect 67010 526170 67078 526226
rect 67134 526170 67202 526226
rect 67258 526170 67326 526226
rect 67382 526170 97674 526226
rect 97730 526170 97798 526226
rect 97854 526170 97922 526226
rect 97978 526170 98046 526226
rect 98102 526170 128394 526226
rect 128450 526170 128518 526226
rect 128574 526170 128642 526226
rect 128698 526170 128766 526226
rect 128822 526170 159114 526226
rect 159170 526170 159238 526226
rect 159294 526170 159362 526226
rect 159418 526170 159486 526226
rect 159542 526170 189834 526226
rect 189890 526170 189958 526226
rect 190014 526170 190082 526226
rect 190138 526170 190206 526226
rect 190262 526170 220554 526226
rect 220610 526170 220678 526226
rect 220734 526170 220802 526226
rect 220858 526170 220926 526226
rect 220982 526170 251274 526226
rect 251330 526170 251398 526226
rect 251454 526170 251522 526226
rect 251578 526170 251646 526226
rect 251702 526170 272518 526226
rect 272574 526170 272642 526226
rect 272698 526170 303238 526226
rect 303294 526170 303362 526226
rect 303418 526170 343434 526226
rect 343490 526170 343558 526226
rect 343614 526170 343682 526226
rect 343738 526170 343806 526226
rect 343862 526170 374154 526226
rect 374210 526170 374278 526226
rect 374334 526170 374402 526226
rect 374458 526170 374526 526226
rect 374582 526170 404874 526226
rect 404930 526170 404998 526226
rect 405054 526170 405122 526226
rect 405178 526170 405246 526226
rect 405302 526170 435594 526226
rect 435650 526170 435718 526226
rect 435774 526170 435842 526226
rect 435898 526170 435966 526226
rect 436022 526170 466314 526226
rect 466370 526170 466438 526226
rect 466494 526170 466562 526226
rect 466618 526170 466686 526226
rect 466742 526170 497034 526226
rect 497090 526170 497158 526226
rect 497214 526170 497282 526226
rect 497338 526170 497406 526226
rect 497462 526170 527754 526226
rect 527810 526170 527878 526226
rect 527934 526170 528002 526226
rect 528058 526170 528126 526226
rect 528182 526170 558474 526226
rect 558530 526170 558598 526226
rect 558654 526170 558722 526226
rect 558778 526170 558846 526226
rect 558902 526170 589194 526226
rect 589250 526170 589318 526226
rect 589374 526170 589442 526226
rect 589498 526170 589566 526226
rect 589622 526170 596496 526226
rect 596552 526170 596620 526226
rect 596676 526170 596744 526226
rect 596800 526170 596868 526226
rect 596924 526170 597980 526226
rect -1916 526102 597980 526170
rect -1916 526046 -860 526102
rect -804 526046 -736 526102
rect -680 526046 -612 526102
rect -556 526046 -488 526102
rect -432 526046 5514 526102
rect 5570 526046 5638 526102
rect 5694 526046 5762 526102
rect 5818 526046 5886 526102
rect 5942 526046 36234 526102
rect 36290 526046 36358 526102
rect 36414 526046 36482 526102
rect 36538 526046 36606 526102
rect 36662 526046 66954 526102
rect 67010 526046 67078 526102
rect 67134 526046 67202 526102
rect 67258 526046 67326 526102
rect 67382 526046 97674 526102
rect 97730 526046 97798 526102
rect 97854 526046 97922 526102
rect 97978 526046 98046 526102
rect 98102 526046 128394 526102
rect 128450 526046 128518 526102
rect 128574 526046 128642 526102
rect 128698 526046 128766 526102
rect 128822 526046 159114 526102
rect 159170 526046 159238 526102
rect 159294 526046 159362 526102
rect 159418 526046 159486 526102
rect 159542 526046 189834 526102
rect 189890 526046 189958 526102
rect 190014 526046 190082 526102
rect 190138 526046 190206 526102
rect 190262 526046 220554 526102
rect 220610 526046 220678 526102
rect 220734 526046 220802 526102
rect 220858 526046 220926 526102
rect 220982 526046 251274 526102
rect 251330 526046 251398 526102
rect 251454 526046 251522 526102
rect 251578 526046 251646 526102
rect 251702 526046 272518 526102
rect 272574 526046 272642 526102
rect 272698 526046 303238 526102
rect 303294 526046 303362 526102
rect 303418 526046 343434 526102
rect 343490 526046 343558 526102
rect 343614 526046 343682 526102
rect 343738 526046 343806 526102
rect 343862 526046 374154 526102
rect 374210 526046 374278 526102
rect 374334 526046 374402 526102
rect 374458 526046 374526 526102
rect 374582 526046 404874 526102
rect 404930 526046 404998 526102
rect 405054 526046 405122 526102
rect 405178 526046 405246 526102
rect 405302 526046 435594 526102
rect 435650 526046 435718 526102
rect 435774 526046 435842 526102
rect 435898 526046 435966 526102
rect 436022 526046 466314 526102
rect 466370 526046 466438 526102
rect 466494 526046 466562 526102
rect 466618 526046 466686 526102
rect 466742 526046 497034 526102
rect 497090 526046 497158 526102
rect 497214 526046 497282 526102
rect 497338 526046 497406 526102
rect 497462 526046 527754 526102
rect 527810 526046 527878 526102
rect 527934 526046 528002 526102
rect 528058 526046 528126 526102
rect 528182 526046 558474 526102
rect 558530 526046 558598 526102
rect 558654 526046 558722 526102
rect 558778 526046 558846 526102
rect 558902 526046 589194 526102
rect 589250 526046 589318 526102
rect 589374 526046 589442 526102
rect 589498 526046 589566 526102
rect 589622 526046 596496 526102
rect 596552 526046 596620 526102
rect 596676 526046 596744 526102
rect 596800 526046 596868 526102
rect 596924 526046 597980 526102
rect -1916 525978 597980 526046
rect -1916 525922 -860 525978
rect -804 525922 -736 525978
rect -680 525922 -612 525978
rect -556 525922 -488 525978
rect -432 525922 5514 525978
rect 5570 525922 5638 525978
rect 5694 525922 5762 525978
rect 5818 525922 5886 525978
rect 5942 525922 36234 525978
rect 36290 525922 36358 525978
rect 36414 525922 36482 525978
rect 36538 525922 36606 525978
rect 36662 525922 66954 525978
rect 67010 525922 67078 525978
rect 67134 525922 67202 525978
rect 67258 525922 67326 525978
rect 67382 525922 97674 525978
rect 97730 525922 97798 525978
rect 97854 525922 97922 525978
rect 97978 525922 98046 525978
rect 98102 525922 128394 525978
rect 128450 525922 128518 525978
rect 128574 525922 128642 525978
rect 128698 525922 128766 525978
rect 128822 525922 159114 525978
rect 159170 525922 159238 525978
rect 159294 525922 159362 525978
rect 159418 525922 159486 525978
rect 159542 525922 189834 525978
rect 189890 525922 189958 525978
rect 190014 525922 190082 525978
rect 190138 525922 190206 525978
rect 190262 525922 220554 525978
rect 220610 525922 220678 525978
rect 220734 525922 220802 525978
rect 220858 525922 220926 525978
rect 220982 525922 251274 525978
rect 251330 525922 251398 525978
rect 251454 525922 251522 525978
rect 251578 525922 251646 525978
rect 251702 525922 272518 525978
rect 272574 525922 272642 525978
rect 272698 525922 303238 525978
rect 303294 525922 303362 525978
rect 303418 525922 343434 525978
rect 343490 525922 343558 525978
rect 343614 525922 343682 525978
rect 343738 525922 343806 525978
rect 343862 525922 374154 525978
rect 374210 525922 374278 525978
rect 374334 525922 374402 525978
rect 374458 525922 374526 525978
rect 374582 525922 404874 525978
rect 404930 525922 404998 525978
rect 405054 525922 405122 525978
rect 405178 525922 405246 525978
rect 405302 525922 435594 525978
rect 435650 525922 435718 525978
rect 435774 525922 435842 525978
rect 435898 525922 435966 525978
rect 436022 525922 466314 525978
rect 466370 525922 466438 525978
rect 466494 525922 466562 525978
rect 466618 525922 466686 525978
rect 466742 525922 497034 525978
rect 497090 525922 497158 525978
rect 497214 525922 497282 525978
rect 497338 525922 497406 525978
rect 497462 525922 527754 525978
rect 527810 525922 527878 525978
rect 527934 525922 528002 525978
rect 528058 525922 528126 525978
rect 528182 525922 558474 525978
rect 558530 525922 558598 525978
rect 558654 525922 558722 525978
rect 558778 525922 558846 525978
rect 558902 525922 589194 525978
rect 589250 525922 589318 525978
rect 589374 525922 589442 525978
rect 589498 525922 589566 525978
rect 589622 525922 596496 525978
rect 596552 525922 596620 525978
rect 596676 525922 596744 525978
rect 596800 525922 596868 525978
rect 596924 525922 597980 525978
rect -1916 525826 597980 525922
rect -1916 514350 597980 514446
rect -1916 514294 -1820 514350
rect -1764 514294 -1696 514350
rect -1640 514294 -1572 514350
rect -1516 514294 -1448 514350
rect -1392 514294 9234 514350
rect 9290 514294 9358 514350
rect 9414 514294 9482 514350
rect 9538 514294 9606 514350
rect 9662 514294 70674 514350
rect 70730 514294 70798 514350
rect 70854 514294 70922 514350
rect 70978 514294 71046 514350
rect 71102 514294 132114 514350
rect 132170 514294 132238 514350
rect 132294 514294 132362 514350
rect 132418 514294 132486 514350
rect 132542 514294 162834 514350
rect 162890 514294 162958 514350
rect 163014 514294 163082 514350
rect 163138 514294 163206 514350
rect 163262 514294 193554 514350
rect 193610 514294 193678 514350
rect 193734 514294 193802 514350
rect 193858 514294 193926 514350
rect 193982 514294 224274 514350
rect 224330 514294 224398 514350
rect 224454 514294 224522 514350
rect 224578 514294 224646 514350
rect 224702 514294 254994 514350
rect 255050 514294 255118 514350
rect 255174 514294 255242 514350
rect 255298 514294 255366 514350
rect 255422 514294 287878 514350
rect 287934 514294 288002 514350
rect 288058 514294 318598 514350
rect 318654 514294 318722 514350
rect 318778 514294 347154 514350
rect 347210 514294 347278 514350
rect 347334 514294 347402 514350
rect 347458 514294 347526 514350
rect 347582 514294 377874 514350
rect 377930 514294 377998 514350
rect 378054 514294 378122 514350
rect 378178 514294 378246 514350
rect 378302 514294 408594 514350
rect 408650 514294 408718 514350
rect 408774 514294 408842 514350
rect 408898 514294 408966 514350
rect 409022 514294 439314 514350
rect 439370 514294 439438 514350
rect 439494 514294 439562 514350
rect 439618 514294 439686 514350
rect 439742 514294 470034 514350
rect 470090 514294 470158 514350
rect 470214 514294 470282 514350
rect 470338 514294 470406 514350
rect 470462 514294 500754 514350
rect 500810 514294 500878 514350
rect 500934 514294 501002 514350
rect 501058 514294 501126 514350
rect 501182 514294 531474 514350
rect 531530 514294 531598 514350
rect 531654 514294 531722 514350
rect 531778 514294 531846 514350
rect 531902 514294 562194 514350
rect 562250 514294 562318 514350
rect 562374 514294 562442 514350
rect 562498 514294 562566 514350
rect 562622 514294 592914 514350
rect 592970 514294 593038 514350
rect 593094 514294 593162 514350
rect 593218 514294 593286 514350
rect 593342 514294 597456 514350
rect 597512 514294 597580 514350
rect 597636 514294 597704 514350
rect 597760 514294 597828 514350
rect 597884 514294 597980 514350
rect -1916 514226 597980 514294
rect -1916 514170 -1820 514226
rect -1764 514170 -1696 514226
rect -1640 514170 -1572 514226
rect -1516 514170 -1448 514226
rect -1392 514170 9234 514226
rect 9290 514170 9358 514226
rect 9414 514170 9482 514226
rect 9538 514170 9606 514226
rect 9662 514170 70674 514226
rect 70730 514170 70798 514226
rect 70854 514170 70922 514226
rect 70978 514170 71046 514226
rect 71102 514170 132114 514226
rect 132170 514170 132238 514226
rect 132294 514170 132362 514226
rect 132418 514170 132486 514226
rect 132542 514170 162834 514226
rect 162890 514170 162958 514226
rect 163014 514170 163082 514226
rect 163138 514170 163206 514226
rect 163262 514170 193554 514226
rect 193610 514170 193678 514226
rect 193734 514170 193802 514226
rect 193858 514170 193926 514226
rect 193982 514170 224274 514226
rect 224330 514170 224398 514226
rect 224454 514170 224522 514226
rect 224578 514170 224646 514226
rect 224702 514170 254994 514226
rect 255050 514170 255118 514226
rect 255174 514170 255242 514226
rect 255298 514170 255366 514226
rect 255422 514170 287878 514226
rect 287934 514170 288002 514226
rect 288058 514170 318598 514226
rect 318654 514170 318722 514226
rect 318778 514170 347154 514226
rect 347210 514170 347278 514226
rect 347334 514170 347402 514226
rect 347458 514170 347526 514226
rect 347582 514170 377874 514226
rect 377930 514170 377998 514226
rect 378054 514170 378122 514226
rect 378178 514170 378246 514226
rect 378302 514170 408594 514226
rect 408650 514170 408718 514226
rect 408774 514170 408842 514226
rect 408898 514170 408966 514226
rect 409022 514170 439314 514226
rect 439370 514170 439438 514226
rect 439494 514170 439562 514226
rect 439618 514170 439686 514226
rect 439742 514170 470034 514226
rect 470090 514170 470158 514226
rect 470214 514170 470282 514226
rect 470338 514170 470406 514226
rect 470462 514170 500754 514226
rect 500810 514170 500878 514226
rect 500934 514170 501002 514226
rect 501058 514170 501126 514226
rect 501182 514170 531474 514226
rect 531530 514170 531598 514226
rect 531654 514170 531722 514226
rect 531778 514170 531846 514226
rect 531902 514170 562194 514226
rect 562250 514170 562318 514226
rect 562374 514170 562442 514226
rect 562498 514170 562566 514226
rect 562622 514170 592914 514226
rect 592970 514170 593038 514226
rect 593094 514170 593162 514226
rect 593218 514170 593286 514226
rect 593342 514170 597456 514226
rect 597512 514170 597580 514226
rect 597636 514170 597704 514226
rect 597760 514170 597828 514226
rect 597884 514170 597980 514226
rect -1916 514102 597980 514170
rect -1916 514046 -1820 514102
rect -1764 514046 -1696 514102
rect -1640 514046 -1572 514102
rect -1516 514046 -1448 514102
rect -1392 514046 9234 514102
rect 9290 514046 9358 514102
rect 9414 514046 9482 514102
rect 9538 514046 9606 514102
rect 9662 514046 70674 514102
rect 70730 514046 70798 514102
rect 70854 514046 70922 514102
rect 70978 514046 71046 514102
rect 71102 514046 132114 514102
rect 132170 514046 132238 514102
rect 132294 514046 132362 514102
rect 132418 514046 132486 514102
rect 132542 514046 162834 514102
rect 162890 514046 162958 514102
rect 163014 514046 163082 514102
rect 163138 514046 163206 514102
rect 163262 514046 193554 514102
rect 193610 514046 193678 514102
rect 193734 514046 193802 514102
rect 193858 514046 193926 514102
rect 193982 514046 224274 514102
rect 224330 514046 224398 514102
rect 224454 514046 224522 514102
rect 224578 514046 224646 514102
rect 224702 514046 254994 514102
rect 255050 514046 255118 514102
rect 255174 514046 255242 514102
rect 255298 514046 255366 514102
rect 255422 514046 287878 514102
rect 287934 514046 288002 514102
rect 288058 514046 318598 514102
rect 318654 514046 318722 514102
rect 318778 514046 347154 514102
rect 347210 514046 347278 514102
rect 347334 514046 347402 514102
rect 347458 514046 347526 514102
rect 347582 514046 377874 514102
rect 377930 514046 377998 514102
rect 378054 514046 378122 514102
rect 378178 514046 378246 514102
rect 378302 514046 408594 514102
rect 408650 514046 408718 514102
rect 408774 514046 408842 514102
rect 408898 514046 408966 514102
rect 409022 514046 439314 514102
rect 439370 514046 439438 514102
rect 439494 514046 439562 514102
rect 439618 514046 439686 514102
rect 439742 514046 470034 514102
rect 470090 514046 470158 514102
rect 470214 514046 470282 514102
rect 470338 514046 470406 514102
rect 470462 514046 500754 514102
rect 500810 514046 500878 514102
rect 500934 514046 501002 514102
rect 501058 514046 501126 514102
rect 501182 514046 531474 514102
rect 531530 514046 531598 514102
rect 531654 514046 531722 514102
rect 531778 514046 531846 514102
rect 531902 514046 562194 514102
rect 562250 514046 562318 514102
rect 562374 514046 562442 514102
rect 562498 514046 562566 514102
rect 562622 514046 592914 514102
rect 592970 514046 593038 514102
rect 593094 514046 593162 514102
rect 593218 514046 593286 514102
rect 593342 514046 597456 514102
rect 597512 514046 597580 514102
rect 597636 514046 597704 514102
rect 597760 514046 597828 514102
rect 597884 514046 597980 514102
rect -1916 513978 597980 514046
rect -1916 513922 -1820 513978
rect -1764 513922 -1696 513978
rect -1640 513922 -1572 513978
rect -1516 513922 -1448 513978
rect -1392 513922 9234 513978
rect 9290 513922 9358 513978
rect 9414 513922 9482 513978
rect 9538 513922 9606 513978
rect 9662 513922 70674 513978
rect 70730 513922 70798 513978
rect 70854 513922 70922 513978
rect 70978 513922 71046 513978
rect 71102 513922 132114 513978
rect 132170 513922 132238 513978
rect 132294 513922 132362 513978
rect 132418 513922 132486 513978
rect 132542 513922 162834 513978
rect 162890 513922 162958 513978
rect 163014 513922 163082 513978
rect 163138 513922 163206 513978
rect 163262 513922 193554 513978
rect 193610 513922 193678 513978
rect 193734 513922 193802 513978
rect 193858 513922 193926 513978
rect 193982 513922 224274 513978
rect 224330 513922 224398 513978
rect 224454 513922 224522 513978
rect 224578 513922 224646 513978
rect 224702 513922 254994 513978
rect 255050 513922 255118 513978
rect 255174 513922 255242 513978
rect 255298 513922 255366 513978
rect 255422 513922 287878 513978
rect 287934 513922 288002 513978
rect 288058 513922 318598 513978
rect 318654 513922 318722 513978
rect 318778 513922 347154 513978
rect 347210 513922 347278 513978
rect 347334 513922 347402 513978
rect 347458 513922 347526 513978
rect 347582 513922 377874 513978
rect 377930 513922 377998 513978
rect 378054 513922 378122 513978
rect 378178 513922 378246 513978
rect 378302 513922 408594 513978
rect 408650 513922 408718 513978
rect 408774 513922 408842 513978
rect 408898 513922 408966 513978
rect 409022 513922 439314 513978
rect 439370 513922 439438 513978
rect 439494 513922 439562 513978
rect 439618 513922 439686 513978
rect 439742 513922 470034 513978
rect 470090 513922 470158 513978
rect 470214 513922 470282 513978
rect 470338 513922 470406 513978
rect 470462 513922 500754 513978
rect 500810 513922 500878 513978
rect 500934 513922 501002 513978
rect 501058 513922 501126 513978
rect 501182 513922 531474 513978
rect 531530 513922 531598 513978
rect 531654 513922 531722 513978
rect 531778 513922 531846 513978
rect 531902 513922 562194 513978
rect 562250 513922 562318 513978
rect 562374 513922 562442 513978
rect 562498 513922 562566 513978
rect 562622 513922 592914 513978
rect 592970 513922 593038 513978
rect 593094 513922 593162 513978
rect 593218 513922 593286 513978
rect 593342 513922 597456 513978
rect 597512 513922 597580 513978
rect 597636 513922 597704 513978
rect 597760 513922 597828 513978
rect 597884 513922 597980 513978
rect -1916 513826 597980 513922
rect -1916 508350 597980 508446
rect -1916 508294 -860 508350
rect -804 508294 -736 508350
rect -680 508294 -612 508350
rect -556 508294 -488 508350
rect -432 508294 5514 508350
rect 5570 508294 5638 508350
rect 5694 508294 5762 508350
rect 5818 508294 5886 508350
rect 5942 508294 36234 508350
rect 36290 508294 36358 508350
rect 36414 508294 36482 508350
rect 36538 508294 36606 508350
rect 36662 508294 66954 508350
rect 67010 508294 67078 508350
rect 67134 508294 67202 508350
rect 67258 508294 67326 508350
rect 67382 508294 97674 508350
rect 97730 508294 97798 508350
rect 97854 508294 97922 508350
rect 97978 508294 98046 508350
rect 98102 508294 128394 508350
rect 128450 508294 128518 508350
rect 128574 508294 128642 508350
rect 128698 508294 128766 508350
rect 128822 508294 159114 508350
rect 159170 508294 159238 508350
rect 159294 508294 159362 508350
rect 159418 508294 159486 508350
rect 159542 508294 189834 508350
rect 189890 508294 189958 508350
rect 190014 508294 190082 508350
rect 190138 508294 190206 508350
rect 190262 508294 220554 508350
rect 220610 508294 220678 508350
rect 220734 508294 220802 508350
rect 220858 508294 220926 508350
rect 220982 508294 251274 508350
rect 251330 508294 251398 508350
rect 251454 508294 251522 508350
rect 251578 508294 251646 508350
rect 251702 508294 272518 508350
rect 272574 508294 272642 508350
rect 272698 508294 303238 508350
rect 303294 508294 303362 508350
rect 303418 508294 343434 508350
rect 343490 508294 343558 508350
rect 343614 508294 343682 508350
rect 343738 508294 343806 508350
rect 343862 508294 374154 508350
rect 374210 508294 374278 508350
rect 374334 508294 374402 508350
rect 374458 508294 374526 508350
rect 374582 508294 404874 508350
rect 404930 508294 404998 508350
rect 405054 508294 405122 508350
rect 405178 508294 405246 508350
rect 405302 508294 435594 508350
rect 435650 508294 435718 508350
rect 435774 508294 435842 508350
rect 435898 508294 435966 508350
rect 436022 508294 466314 508350
rect 466370 508294 466438 508350
rect 466494 508294 466562 508350
rect 466618 508294 466686 508350
rect 466742 508294 497034 508350
rect 497090 508294 497158 508350
rect 497214 508294 497282 508350
rect 497338 508294 497406 508350
rect 497462 508294 527754 508350
rect 527810 508294 527878 508350
rect 527934 508294 528002 508350
rect 528058 508294 528126 508350
rect 528182 508294 558474 508350
rect 558530 508294 558598 508350
rect 558654 508294 558722 508350
rect 558778 508294 558846 508350
rect 558902 508294 589194 508350
rect 589250 508294 589318 508350
rect 589374 508294 589442 508350
rect 589498 508294 589566 508350
rect 589622 508294 596496 508350
rect 596552 508294 596620 508350
rect 596676 508294 596744 508350
rect 596800 508294 596868 508350
rect 596924 508294 597980 508350
rect -1916 508226 597980 508294
rect -1916 508170 -860 508226
rect -804 508170 -736 508226
rect -680 508170 -612 508226
rect -556 508170 -488 508226
rect -432 508170 5514 508226
rect 5570 508170 5638 508226
rect 5694 508170 5762 508226
rect 5818 508170 5886 508226
rect 5942 508170 36234 508226
rect 36290 508170 36358 508226
rect 36414 508170 36482 508226
rect 36538 508170 36606 508226
rect 36662 508170 66954 508226
rect 67010 508170 67078 508226
rect 67134 508170 67202 508226
rect 67258 508170 67326 508226
rect 67382 508170 97674 508226
rect 97730 508170 97798 508226
rect 97854 508170 97922 508226
rect 97978 508170 98046 508226
rect 98102 508170 128394 508226
rect 128450 508170 128518 508226
rect 128574 508170 128642 508226
rect 128698 508170 128766 508226
rect 128822 508170 159114 508226
rect 159170 508170 159238 508226
rect 159294 508170 159362 508226
rect 159418 508170 159486 508226
rect 159542 508170 189834 508226
rect 189890 508170 189958 508226
rect 190014 508170 190082 508226
rect 190138 508170 190206 508226
rect 190262 508170 220554 508226
rect 220610 508170 220678 508226
rect 220734 508170 220802 508226
rect 220858 508170 220926 508226
rect 220982 508170 251274 508226
rect 251330 508170 251398 508226
rect 251454 508170 251522 508226
rect 251578 508170 251646 508226
rect 251702 508170 272518 508226
rect 272574 508170 272642 508226
rect 272698 508170 303238 508226
rect 303294 508170 303362 508226
rect 303418 508170 343434 508226
rect 343490 508170 343558 508226
rect 343614 508170 343682 508226
rect 343738 508170 343806 508226
rect 343862 508170 374154 508226
rect 374210 508170 374278 508226
rect 374334 508170 374402 508226
rect 374458 508170 374526 508226
rect 374582 508170 404874 508226
rect 404930 508170 404998 508226
rect 405054 508170 405122 508226
rect 405178 508170 405246 508226
rect 405302 508170 435594 508226
rect 435650 508170 435718 508226
rect 435774 508170 435842 508226
rect 435898 508170 435966 508226
rect 436022 508170 466314 508226
rect 466370 508170 466438 508226
rect 466494 508170 466562 508226
rect 466618 508170 466686 508226
rect 466742 508170 497034 508226
rect 497090 508170 497158 508226
rect 497214 508170 497282 508226
rect 497338 508170 497406 508226
rect 497462 508170 527754 508226
rect 527810 508170 527878 508226
rect 527934 508170 528002 508226
rect 528058 508170 528126 508226
rect 528182 508170 558474 508226
rect 558530 508170 558598 508226
rect 558654 508170 558722 508226
rect 558778 508170 558846 508226
rect 558902 508170 589194 508226
rect 589250 508170 589318 508226
rect 589374 508170 589442 508226
rect 589498 508170 589566 508226
rect 589622 508170 596496 508226
rect 596552 508170 596620 508226
rect 596676 508170 596744 508226
rect 596800 508170 596868 508226
rect 596924 508170 597980 508226
rect -1916 508102 597980 508170
rect -1916 508046 -860 508102
rect -804 508046 -736 508102
rect -680 508046 -612 508102
rect -556 508046 -488 508102
rect -432 508046 5514 508102
rect 5570 508046 5638 508102
rect 5694 508046 5762 508102
rect 5818 508046 5886 508102
rect 5942 508046 36234 508102
rect 36290 508046 36358 508102
rect 36414 508046 36482 508102
rect 36538 508046 36606 508102
rect 36662 508046 66954 508102
rect 67010 508046 67078 508102
rect 67134 508046 67202 508102
rect 67258 508046 67326 508102
rect 67382 508046 97674 508102
rect 97730 508046 97798 508102
rect 97854 508046 97922 508102
rect 97978 508046 98046 508102
rect 98102 508046 128394 508102
rect 128450 508046 128518 508102
rect 128574 508046 128642 508102
rect 128698 508046 128766 508102
rect 128822 508046 159114 508102
rect 159170 508046 159238 508102
rect 159294 508046 159362 508102
rect 159418 508046 159486 508102
rect 159542 508046 189834 508102
rect 189890 508046 189958 508102
rect 190014 508046 190082 508102
rect 190138 508046 190206 508102
rect 190262 508046 220554 508102
rect 220610 508046 220678 508102
rect 220734 508046 220802 508102
rect 220858 508046 220926 508102
rect 220982 508046 251274 508102
rect 251330 508046 251398 508102
rect 251454 508046 251522 508102
rect 251578 508046 251646 508102
rect 251702 508046 272518 508102
rect 272574 508046 272642 508102
rect 272698 508046 303238 508102
rect 303294 508046 303362 508102
rect 303418 508046 343434 508102
rect 343490 508046 343558 508102
rect 343614 508046 343682 508102
rect 343738 508046 343806 508102
rect 343862 508046 374154 508102
rect 374210 508046 374278 508102
rect 374334 508046 374402 508102
rect 374458 508046 374526 508102
rect 374582 508046 404874 508102
rect 404930 508046 404998 508102
rect 405054 508046 405122 508102
rect 405178 508046 405246 508102
rect 405302 508046 435594 508102
rect 435650 508046 435718 508102
rect 435774 508046 435842 508102
rect 435898 508046 435966 508102
rect 436022 508046 466314 508102
rect 466370 508046 466438 508102
rect 466494 508046 466562 508102
rect 466618 508046 466686 508102
rect 466742 508046 497034 508102
rect 497090 508046 497158 508102
rect 497214 508046 497282 508102
rect 497338 508046 497406 508102
rect 497462 508046 527754 508102
rect 527810 508046 527878 508102
rect 527934 508046 528002 508102
rect 528058 508046 528126 508102
rect 528182 508046 558474 508102
rect 558530 508046 558598 508102
rect 558654 508046 558722 508102
rect 558778 508046 558846 508102
rect 558902 508046 589194 508102
rect 589250 508046 589318 508102
rect 589374 508046 589442 508102
rect 589498 508046 589566 508102
rect 589622 508046 596496 508102
rect 596552 508046 596620 508102
rect 596676 508046 596744 508102
rect 596800 508046 596868 508102
rect 596924 508046 597980 508102
rect -1916 507978 597980 508046
rect -1916 507922 -860 507978
rect -804 507922 -736 507978
rect -680 507922 -612 507978
rect -556 507922 -488 507978
rect -432 507922 5514 507978
rect 5570 507922 5638 507978
rect 5694 507922 5762 507978
rect 5818 507922 5886 507978
rect 5942 507922 36234 507978
rect 36290 507922 36358 507978
rect 36414 507922 36482 507978
rect 36538 507922 36606 507978
rect 36662 507922 66954 507978
rect 67010 507922 67078 507978
rect 67134 507922 67202 507978
rect 67258 507922 67326 507978
rect 67382 507922 97674 507978
rect 97730 507922 97798 507978
rect 97854 507922 97922 507978
rect 97978 507922 98046 507978
rect 98102 507922 128394 507978
rect 128450 507922 128518 507978
rect 128574 507922 128642 507978
rect 128698 507922 128766 507978
rect 128822 507922 159114 507978
rect 159170 507922 159238 507978
rect 159294 507922 159362 507978
rect 159418 507922 159486 507978
rect 159542 507922 189834 507978
rect 189890 507922 189958 507978
rect 190014 507922 190082 507978
rect 190138 507922 190206 507978
rect 190262 507922 220554 507978
rect 220610 507922 220678 507978
rect 220734 507922 220802 507978
rect 220858 507922 220926 507978
rect 220982 507922 251274 507978
rect 251330 507922 251398 507978
rect 251454 507922 251522 507978
rect 251578 507922 251646 507978
rect 251702 507922 272518 507978
rect 272574 507922 272642 507978
rect 272698 507922 303238 507978
rect 303294 507922 303362 507978
rect 303418 507922 343434 507978
rect 343490 507922 343558 507978
rect 343614 507922 343682 507978
rect 343738 507922 343806 507978
rect 343862 507922 374154 507978
rect 374210 507922 374278 507978
rect 374334 507922 374402 507978
rect 374458 507922 374526 507978
rect 374582 507922 404874 507978
rect 404930 507922 404998 507978
rect 405054 507922 405122 507978
rect 405178 507922 405246 507978
rect 405302 507922 435594 507978
rect 435650 507922 435718 507978
rect 435774 507922 435842 507978
rect 435898 507922 435966 507978
rect 436022 507922 466314 507978
rect 466370 507922 466438 507978
rect 466494 507922 466562 507978
rect 466618 507922 466686 507978
rect 466742 507922 497034 507978
rect 497090 507922 497158 507978
rect 497214 507922 497282 507978
rect 497338 507922 497406 507978
rect 497462 507922 527754 507978
rect 527810 507922 527878 507978
rect 527934 507922 528002 507978
rect 528058 507922 528126 507978
rect 528182 507922 558474 507978
rect 558530 507922 558598 507978
rect 558654 507922 558722 507978
rect 558778 507922 558846 507978
rect 558902 507922 589194 507978
rect 589250 507922 589318 507978
rect 589374 507922 589442 507978
rect 589498 507922 589566 507978
rect 589622 507922 596496 507978
rect 596552 507922 596620 507978
rect 596676 507922 596744 507978
rect 596800 507922 596868 507978
rect 596924 507922 597980 507978
rect -1916 507826 597980 507922
rect -1916 496350 597980 496446
rect -1916 496294 -1820 496350
rect -1764 496294 -1696 496350
rect -1640 496294 -1572 496350
rect -1516 496294 -1448 496350
rect -1392 496294 9234 496350
rect 9290 496294 9358 496350
rect 9414 496294 9482 496350
rect 9538 496294 9606 496350
rect 9662 496294 70674 496350
rect 70730 496294 70798 496350
rect 70854 496294 70922 496350
rect 70978 496294 71046 496350
rect 71102 496294 132114 496350
rect 132170 496294 132238 496350
rect 132294 496294 132362 496350
rect 132418 496294 132486 496350
rect 132542 496294 162834 496350
rect 162890 496294 162958 496350
rect 163014 496294 163082 496350
rect 163138 496294 163206 496350
rect 163262 496294 193554 496350
rect 193610 496294 193678 496350
rect 193734 496294 193802 496350
rect 193858 496294 193926 496350
rect 193982 496294 224274 496350
rect 224330 496294 224398 496350
rect 224454 496294 224522 496350
rect 224578 496294 224646 496350
rect 224702 496294 254994 496350
rect 255050 496294 255118 496350
rect 255174 496294 255242 496350
rect 255298 496294 255366 496350
rect 255422 496294 287878 496350
rect 287934 496294 288002 496350
rect 288058 496294 318598 496350
rect 318654 496294 318722 496350
rect 318778 496294 347154 496350
rect 347210 496294 347278 496350
rect 347334 496294 347402 496350
rect 347458 496294 347526 496350
rect 347582 496294 377874 496350
rect 377930 496294 377998 496350
rect 378054 496294 378122 496350
rect 378178 496294 378246 496350
rect 378302 496294 408594 496350
rect 408650 496294 408718 496350
rect 408774 496294 408842 496350
rect 408898 496294 408966 496350
rect 409022 496294 439314 496350
rect 439370 496294 439438 496350
rect 439494 496294 439562 496350
rect 439618 496294 439686 496350
rect 439742 496294 470034 496350
rect 470090 496294 470158 496350
rect 470214 496294 470282 496350
rect 470338 496294 470406 496350
rect 470462 496294 500754 496350
rect 500810 496294 500878 496350
rect 500934 496294 501002 496350
rect 501058 496294 501126 496350
rect 501182 496294 531474 496350
rect 531530 496294 531598 496350
rect 531654 496294 531722 496350
rect 531778 496294 531846 496350
rect 531902 496294 562194 496350
rect 562250 496294 562318 496350
rect 562374 496294 562442 496350
rect 562498 496294 562566 496350
rect 562622 496294 592914 496350
rect 592970 496294 593038 496350
rect 593094 496294 593162 496350
rect 593218 496294 593286 496350
rect 593342 496294 597456 496350
rect 597512 496294 597580 496350
rect 597636 496294 597704 496350
rect 597760 496294 597828 496350
rect 597884 496294 597980 496350
rect -1916 496226 597980 496294
rect -1916 496170 -1820 496226
rect -1764 496170 -1696 496226
rect -1640 496170 -1572 496226
rect -1516 496170 -1448 496226
rect -1392 496170 9234 496226
rect 9290 496170 9358 496226
rect 9414 496170 9482 496226
rect 9538 496170 9606 496226
rect 9662 496170 70674 496226
rect 70730 496170 70798 496226
rect 70854 496170 70922 496226
rect 70978 496170 71046 496226
rect 71102 496170 132114 496226
rect 132170 496170 132238 496226
rect 132294 496170 132362 496226
rect 132418 496170 132486 496226
rect 132542 496170 162834 496226
rect 162890 496170 162958 496226
rect 163014 496170 163082 496226
rect 163138 496170 163206 496226
rect 163262 496170 193554 496226
rect 193610 496170 193678 496226
rect 193734 496170 193802 496226
rect 193858 496170 193926 496226
rect 193982 496170 224274 496226
rect 224330 496170 224398 496226
rect 224454 496170 224522 496226
rect 224578 496170 224646 496226
rect 224702 496170 254994 496226
rect 255050 496170 255118 496226
rect 255174 496170 255242 496226
rect 255298 496170 255366 496226
rect 255422 496170 287878 496226
rect 287934 496170 288002 496226
rect 288058 496170 318598 496226
rect 318654 496170 318722 496226
rect 318778 496170 347154 496226
rect 347210 496170 347278 496226
rect 347334 496170 347402 496226
rect 347458 496170 347526 496226
rect 347582 496170 377874 496226
rect 377930 496170 377998 496226
rect 378054 496170 378122 496226
rect 378178 496170 378246 496226
rect 378302 496170 408594 496226
rect 408650 496170 408718 496226
rect 408774 496170 408842 496226
rect 408898 496170 408966 496226
rect 409022 496170 439314 496226
rect 439370 496170 439438 496226
rect 439494 496170 439562 496226
rect 439618 496170 439686 496226
rect 439742 496170 470034 496226
rect 470090 496170 470158 496226
rect 470214 496170 470282 496226
rect 470338 496170 470406 496226
rect 470462 496170 500754 496226
rect 500810 496170 500878 496226
rect 500934 496170 501002 496226
rect 501058 496170 501126 496226
rect 501182 496170 531474 496226
rect 531530 496170 531598 496226
rect 531654 496170 531722 496226
rect 531778 496170 531846 496226
rect 531902 496170 562194 496226
rect 562250 496170 562318 496226
rect 562374 496170 562442 496226
rect 562498 496170 562566 496226
rect 562622 496170 592914 496226
rect 592970 496170 593038 496226
rect 593094 496170 593162 496226
rect 593218 496170 593286 496226
rect 593342 496170 597456 496226
rect 597512 496170 597580 496226
rect 597636 496170 597704 496226
rect 597760 496170 597828 496226
rect 597884 496170 597980 496226
rect -1916 496102 597980 496170
rect -1916 496046 -1820 496102
rect -1764 496046 -1696 496102
rect -1640 496046 -1572 496102
rect -1516 496046 -1448 496102
rect -1392 496046 9234 496102
rect 9290 496046 9358 496102
rect 9414 496046 9482 496102
rect 9538 496046 9606 496102
rect 9662 496046 70674 496102
rect 70730 496046 70798 496102
rect 70854 496046 70922 496102
rect 70978 496046 71046 496102
rect 71102 496046 132114 496102
rect 132170 496046 132238 496102
rect 132294 496046 132362 496102
rect 132418 496046 132486 496102
rect 132542 496046 162834 496102
rect 162890 496046 162958 496102
rect 163014 496046 163082 496102
rect 163138 496046 163206 496102
rect 163262 496046 193554 496102
rect 193610 496046 193678 496102
rect 193734 496046 193802 496102
rect 193858 496046 193926 496102
rect 193982 496046 224274 496102
rect 224330 496046 224398 496102
rect 224454 496046 224522 496102
rect 224578 496046 224646 496102
rect 224702 496046 254994 496102
rect 255050 496046 255118 496102
rect 255174 496046 255242 496102
rect 255298 496046 255366 496102
rect 255422 496046 287878 496102
rect 287934 496046 288002 496102
rect 288058 496046 318598 496102
rect 318654 496046 318722 496102
rect 318778 496046 347154 496102
rect 347210 496046 347278 496102
rect 347334 496046 347402 496102
rect 347458 496046 347526 496102
rect 347582 496046 377874 496102
rect 377930 496046 377998 496102
rect 378054 496046 378122 496102
rect 378178 496046 378246 496102
rect 378302 496046 408594 496102
rect 408650 496046 408718 496102
rect 408774 496046 408842 496102
rect 408898 496046 408966 496102
rect 409022 496046 439314 496102
rect 439370 496046 439438 496102
rect 439494 496046 439562 496102
rect 439618 496046 439686 496102
rect 439742 496046 470034 496102
rect 470090 496046 470158 496102
rect 470214 496046 470282 496102
rect 470338 496046 470406 496102
rect 470462 496046 500754 496102
rect 500810 496046 500878 496102
rect 500934 496046 501002 496102
rect 501058 496046 501126 496102
rect 501182 496046 531474 496102
rect 531530 496046 531598 496102
rect 531654 496046 531722 496102
rect 531778 496046 531846 496102
rect 531902 496046 562194 496102
rect 562250 496046 562318 496102
rect 562374 496046 562442 496102
rect 562498 496046 562566 496102
rect 562622 496046 592914 496102
rect 592970 496046 593038 496102
rect 593094 496046 593162 496102
rect 593218 496046 593286 496102
rect 593342 496046 597456 496102
rect 597512 496046 597580 496102
rect 597636 496046 597704 496102
rect 597760 496046 597828 496102
rect 597884 496046 597980 496102
rect -1916 495978 597980 496046
rect -1916 495922 -1820 495978
rect -1764 495922 -1696 495978
rect -1640 495922 -1572 495978
rect -1516 495922 -1448 495978
rect -1392 495922 9234 495978
rect 9290 495922 9358 495978
rect 9414 495922 9482 495978
rect 9538 495922 9606 495978
rect 9662 495922 70674 495978
rect 70730 495922 70798 495978
rect 70854 495922 70922 495978
rect 70978 495922 71046 495978
rect 71102 495922 132114 495978
rect 132170 495922 132238 495978
rect 132294 495922 132362 495978
rect 132418 495922 132486 495978
rect 132542 495922 162834 495978
rect 162890 495922 162958 495978
rect 163014 495922 163082 495978
rect 163138 495922 163206 495978
rect 163262 495922 193554 495978
rect 193610 495922 193678 495978
rect 193734 495922 193802 495978
rect 193858 495922 193926 495978
rect 193982 495922 224274 495978
rect 224330 495922 224398 495978
rect 224454 495922 224522 495978
rect 224578 495922 224646 495978
rect 224702 495922 254994 495978
rect 255050 495922 255118 495978
rect 255174 495922 255242 495978
rect 255298 495922 255366 495978
rect 255422 495922 287878 495978
rect 287934 495922 288002 495978
rect 288058 495922 318598 495978
rect 318654 495922 318722 495978
rect 318778 495922 347154 495978
rect 347210 495922 347278 495978
rect 347334 495922 347402 495978
rect 347458 495922 347526 495978
rect 347582 495922 377874 495978
rect 377930 495922 377998 495978
rect 378054 495922 378122 495978
rect 378178 495922 378246 495978
rect 378302 495922 408594 495978
rect 408650 495922 408718 495978
rect 408774 495922 408842 495978
rect 408898 495922 408966 495978
rect 409022 495922 439314 495978
rect 439370 495922 439438 495978
rect 439494 495922 439562 495978
rect 439618 495922 439686 495978
rect 439742 495922 470034 495978
rect 470090 495922 470158 495978
rect 470214 495922 470282 495978
rect 470338 495922 470406 495978
rect 470462 495922 500754 495978
rect 500810 495922 500878 495978
rect 500934 495922 501002 495978
rect 501058 495922 501126 495978
rect 501182 495922 531474 495978
rect 531530 495922 531598 495978
rect 531654 495922 531722 495978
rect 531778 495922 531846 495978
rect 531902 495922 562194 495978
rect 562250 495922 562318 495978
rect 562374 495922 562442 495978
rect 562498 495922 562566 495978
rect 562622 495922 592914 495978
rect 592970 495922 593038 495978
rect 593094 495922 593162 495978
rect 593218 495922 593286 495978
rect 593342 495922 597456 495978
rect 597512 495922 597580 495978
rect 597636 495922 597704 495978
rect 597760 495922 597828 495978
rect 597884 495922 597980 495978
rect -1916 495826 597980 495922
rect -1916 490350 597980 490446
rect -1916 490294 -860 490350
rect -804 490294 -736 490350
rect -680 490294 -612 490350
rect -556 490294 -488 490350
rect -432 490294 5514 490350
rect 5570 490294 5638 490350
rect 5694 490294 5762 490350
rect 5818 490294 5886 490350
rect 5942 490294 24518 490350
rect 24574 490294 24642 490350
rect 24698 490294 36234 490350
rect 36290 490294 36358 490350
rect 36414 490294 36482 490350
rect 36538 490294 36606 490350
rect 36662 490294 55238 490350
rect 55294 490294 55362 490350
rect 55418 490294 66954 490350
rect 67010 490294 67078 490350
rect 67134 490294 67202 490350
rect 67258 490294 67326 490350
rect 67382 490294 86518 490350
rect 86574 490294 86642 490350
rect 86698 490294 97674 490350
rect 97730 490294 97798 490350
rect 97854 490294 97922 490350
rect 97978 490294 98046 490350
rect 98102 490294 117238 490350
rect 117294 490294 117362 490350
rect 117418 490294 128394 490350
rect 128450 490294 128518 490350
rect 128574 490294 128642 490350
rect 128698 490294 128766 490350
rect 128822 490294 148518 490350
rect 148574 490294 148642 490350
rect 148698 490294 159114 490350
rect 159170 490294 159238 490350
rect 159294 490294 159362 490350
rect 159418 490294 159486 490350
rect 159542 490294 179238 490350
rect 179294 490294 179362 490350
rect 179418 490294 189834 490350
rect 189890 490294 189958 490350
rect 190014 490294 190082 490350
rect 190138 490294 190206 490350
rect 190262 490294 210518 490350
rect 210574 490294 210642 490350
rect 210698 490294 220554 490350
rect 220610 490294 220678 490350
rect 220734 490294 220802 490350
rect 220858 490294 220926 490350
rect 220982 490294 241238 490350
rect 241294 490294 241362 490350
rect 241418 490294 251274 490350
rect 251330 490294 251398 490350
rect 251454 490294 251522 490350
rect 251578 490294 251646 490350
rect 251702 490294 272518 490350
rect 272574 490294 272642 490350
rect 272698 490294 303238 490350
rect 303294 490294 303362 490350
rect 303418 490294 343434 490350
rect 343490 490294 343558 490350
rect 343614 490294 343682 490350
rect 343738 490294 343806 490350
rect 343862 490294 356518 490350
rect 356574 490294 356642 490350
rect 356698 490294 374154 490350
rect 374210 490294 374278 490350
rect 374334 490294 374402 490350
rect 374458 490294 374526 490350
rect 374582 490294 387238 490350
rect 387294 490294 387362 490350
rect 387418 490294 404874 490350
rect 404930 490294 404998 490350
rect 405054 490294 405122 490350
rect 405178 490294 405246 490350
rect 405302 490294 418518 490350
rect 418574 490294 418642 490350
rect 418698 490294 435594 490350
rect 435650 490294 435718 490350
rect 435774 490294 435842 490350
rect 435898 490294 435966 490350
rect 436022 490294 449238 490350
rect 449294 490294 449362 490350
rect 449418 490294 466314 490350
rect 466370 490294 466438 490350
rect 466494 490294 466562 490350
rect 466618 490294 466686 490350
rect 466742 490294 480518 490350
rect 480574 490294 480642 490350
rect 480698 490294 497034 490350
rect 497090 490294 497158 490350
rect 497214 490294 497282 490350
rect 497338 490294 497406 490350
rect 497462 490294 511238 490350
rect 511294 490294 511362 490350
rect 511418 490294 527754 490350
rect 527810 490294 527878 490350
rect 527934 490294 528002 490350
rect 528058 490294 528126 490350
rect 528182 490294 542518 490350
rect 542574 490294 542642 490350
rect 542698 490294 558474 490350
rect 558530 490294 558598 490350
rect 558654 490294 558722 490350
rect 558778 490294 558846 490350
rect 558902 490294 573238 490350
rect 573294 490294 573362 490350
rect 573418 490294 589194 490350
rect 589250 490294 589318 490350
rect 589374 490294 589442 490350
rect 589498 490294 589566 490350
rect 589622 490294 596496 490350
rect 596552 490294 596620 490350
rect 596676 490294 596744 490350
rect 596800 490294 596868 490350
rect 596924 490294 597980 490350
rect -1916 490226 597980 490294
rect -1916 490170 -860 490226
rect -804 490170 -736 490226
rect -680 490170 -612 490226
rect -556 490170 -488 490226
rect -432 490170 5514 490226
rect 5570 490170 5638 490226
rect 5694 490170 5762 490226
rect 5818 490170 5886 490226
rect 5942 490170 24518 490226
rect 24574 490170 24642 490226
rect 24698 490170 36234 490226
rect 36290 490170 36358 490226
rect 36414 490170 36482 490226
rect 36538 490170 36606 490226
rect 36662 490170 55238 490226
rect 55294 490170 55362 490226
rect 55418 490170 66954 490226
rect 67010 490170 67078 490226
rect 67134 490170 67202 490226
rect 67258 490170 67326 490226
rect 67382 490170 86518 490226
rect 86574 490170 86642 490226
rect 86698 490170 97674 490226
rect 97730 490170 97798 490226
rect 97854 490170 97922 490226
rect 97978 490170 98046 490226
rect 98102 490170 117238 490226
rect 117294 490170 117362 490226
rect 117418 490170 128394 490226
rect 128450 490170 128518 490226
rect 128574 490170 128642 490226
rect 128698 490170 128766 490226
rect 128822 490170 148518 490226
rect 148574 490170 148642 490226
rect 148698 490170 159114 490226
rect 159170 490170 159238 490226
rect 159294 490170 159362 490226
rect 159418 490170 159486 490226
rect 159542 490170 179238 490226
rect 179294 490170 179362 490226
rect 179418 490170 189834 490226
rect 189890 490170 189958 490226
rect 190014 490170 190082 490226
rect 190138 490170 190206 490226
rect 190262 490170 210518 490226
rect 210574 490170 210642 490226
rect 210698 490170 220554 490226
rect 220610 490170 220678 490226
rect 220734 490170 220802 490226
rect 220858 490170 220926 490226
rect 220982 490170 241238 490226
rect 241294 490170 241362 490226
rect 241418 490170 251274 490226
rect 251330 490170 251398 490226
rect 251454 490170 251522 490226
rect 251578 490170 251646 490226
rect 251702 490170 272518 490226
rect 272574 490170 272642 490226
rect 272698 490170 303238 490226
rect 303294 490170 303362 490226
rect 303418 490170 343434 490226
rect 343490 490170 343558 490226
rect 343614 490170 343682 490226
rect 343738 490170 343806 490226
rect 343862 490170 356518 490226
rect 356574 490170 356642 490226
rect 356698 490170 374154 490226
rect 374210 490170 374278 490226
rect 374334 490170 374402 490226
rect 374458 490170 374526 490226
rect 374582 490170 387238 490226
rect 387294 490170 387362 490226
rect 387418 490170 404874 490226
rect 404930 490170 404998 490226
rect 405054 490170 405122 490226
rect 405178 490170 405246 490226
rect 405302 490170 418518 490226
rect 418574 490170 418642 490226
rect 418698 490170 435594 490226
rect 435650 490170 435718 490226
rect 435774 490170 435842 490226
rect 435898 490170 435966 490226
rect 436022 490170 449238 490226
rect 449294 490170 449362 490226
rect 449418 490170 466314 490226
rect 466370 490170 466438 490226
rect 466494 490170 466562 490226
rect 466618 490170 466686 490226
rect 466742 490170 480518 490226
rect 480574 490170 480642 490226
rect 480698 490170 497034 490226
rect 497090 490170 497158 490226
rect 497214 490170 497282 490226
rect 497338 490170 497406 490226
rect 497462 490170 511238 490226
rect 511294 490170 511362 490226
rect 511418 490170 527754 490226
rect 527810 490170 527878 490226
rect 527934 490170 528002 490226
rect 528058 490170 528126 490226
rect 528182 490170 542518 490226
rect 542574 490170 542642 490226
rect 542698 490170 558474 490226
rect 558530 490170 558598 490226
rect 558654 490170 558722 490226
rect 558778 490170 558846 490226
rect 558902 490170 573238 490226
rect 573294 490170 573362 490226
rect 573418 490170 589194 490226
rect 589250 490170 589318 490226
rect 589374 490170 589442 490226
rect 589498 490170 589566 490226
rect 589622 490170 596496 490226
rect 596552 490170 596620 490226
rect 596676 490170 596744 490226
rect 596800 490170 596868 490226
rect 596924 490170 597980 490226
rect -1916 490102 597980 490170
rect -1916 490046 -860 490102
rect -804 490046 -736 490102
rect -680 490046 -612 490102
rect -556 490046 -488 490102
rect -432 490046 5514 490102
rect 5570 490046 5638 490102
rect 5694 490046 5762 490102
rect 5818 490046 5886 490102
rect 5942 490046 24518 490102
rect 24574 490046 24642 490102
rect 24698 490046 36234 490102
rect 36290 490046 36358 490102
rect 36414 490046 36482 490102
rect 36538 490046 36606 490102
rect 36662 490046 55238 490102
rect 55294 490046 55362 490102
rect 55418 490046 66954 490102
rect 67010 490046 67078 490102
rect 67134 490046 67202 490102
rect 67258 490046 67326 490102
rect 67382 490046 86518 490102
rect 86574 490046 86642 490102
rect 86698 490046 97674 490102
rect 97730 490046 97798 490102
rect 97854 490046 97922 490102
rect 97978 490046 98046 490102
rect 98102 490046 117238 490102
rect 117294 490046 117362 490102
rect 117418 490046 128394 490102
rect 128450 490046 128518 490102
rect 128574 490046 128642 490102
rect 128698 490046 128766 490102
rect 128822 490046 148518 490102
rect 148574 490046 148642 490102
rect 148698 490046 159114 490102
rect 159170 490046 159238 490102
rect 159294 490046 159362 490102
rect 159418 490046 159486 490102
rect 159542 490046 179238 490102
rect 179294 490046 179362 490102
rect 179418 490046 189834 490102
rect 189890 490046 189958 490102
rect 190014 490046 190082 490102
rect 190138 490046 190206 490102
rect 190262 490046 210518 490102
rect 210574 490046 210642 490102
rect 210698 490046 220554 490102
rect 220610 490046 220678 490102
rect 220734 490046 220802 490102
rect 220858 490046 220926 490102
rect 220982 490046 241238 490102
rect 241294 490046 241362 490102
rect 241418 490046 251274 490102
rect 251330 490046 251398 490102
rect 251454 490046 251522 490102
rect 251578 490046 251646 490102
rect 251702 490046 272518 490102
rect 272574 490046 272642 490102
rect 272698 490046 303238 490102
rect 303294 490046 303362 490102
rect 303418 490046 343434 490102
rect 343490 490046 343558 490102
rect 343614 490046 343682 490102
rect 343738 490046 343806 490102
rect 343862 490046 356518 490102
rect 356574 490046 356642 490102
rect 356698 490046 374154 490102
rect 374210 490046 374278 490102
rect 374334 490046 374402 490102
rect 374458 490046 374526 490102
rect 374582 490046 387238 490102
rect 387294 490046 387362 490102
rect 387418 490046 404874 490102
rect 404930 490046 404998 490102
rect 405054 490046 405122 490102
rect 405178 490046 405246 490102
rect 405302 490046 418518 490102
rect 418574 490046 418642 490102
rect 418698 490046 435594 490102
rect 435650 490046 435718 490102
rect 435774 490046 435842 490102
rect 435898 490046 435966 490102
rect 436022 490046 449238 490102
rect 449294 490046 449362 490102
rect 449418 490046 466314 490102
rect 466370 490046 466438 490102
rect 466494 490046 466562 490102
rect 466618 490046 466686 490102
rect 466742 490046 480518 490102
rect 480574 490046 480642 490102
rect 480698 490046 497034 490102
rect 497090 490046 497158 490102
rect 497214 490046 497282 490102
rect 497338 490046 497406 490102
rect 497462 490046 511238 490102
rect 511294 490046 511362 490102
rect 511418 490046 527754 490102
rect 527810 490046 527878 490102
rect 527934 490046 528002 490102
rect 528058 490046 528126 490102
rect 528182 490046 542518 490102
rect 542574 490046 542642 490102
rect 542698 490046 558474 490102
rect 558530 490046 558598 490102
rect 558654 490046 558722 490102
rect 558778 490046 558846 490102
rect 558902 490046 573238 490102
rect 573294 490046 573362 490102
rect 573418 490046 589194 490102
rect 589250 490046 589318 490102
rect 589374 490046 589442 490102
rect 589498 490046 589566 490102
rect 589622 490046 596496 490102
rect 596552 490046 596620 490102
rect 596676 490046 596744 490102
rect 596800 490046 596868 490102
rect 596924 490046 597980 490102
rect -1916 489978 597980 490046
rect -1916 489922 -860 489978
rect -804 489922 -736 489978
rect -680 489922 -612 489978
rect -556 489922 -488 489978
rect -432 489922 5514 489978
rect 5570 489922 5638 489978
rect 5694 489922 5762 489978
rect 5818 489922 5886 489978
rect 5942 489922 24518 489978
rect 24574 489922 24642 489978
rect 24698 489922 36234 489978
rect 36290 489922 36358 489978
rect 36414 489922 36482 489978
rect 36538 489922 36606 489978
rect 36662 489922 55238 489978
rect 55294 489922 55362 489978
rect 55418 489922 66954 489978
rect 67010 489922 67078 489978
rect 67134 489922 67202 489978
rect 67258 489922 67326 489978
rect 67382 489922 86518 489978
rect 86574 489922 86642 489978
rect 86698 489922 97674 489978
rect 97730 489922 97798 489978
rect 97854 489922 97922 489978
rect 97978 489922 98046 489978
rect 98102 489922 117238 489978
rect 117294 489922 117362 489978
rect 117418 489922 128394 489978
rect 128450 489922 128518 489978
rect 128574 489922 128642 489978
rect 128698 489922 128766 489978
rect 128822 489922 148518 489978
rect 148574 489922 148642 489978
rect 148698 489922 159114 489978
rect 159170 489922 159238 489978
rect 159294 489922 159362 489978
rect 159418 489922 159486 489978
rect 159542 489922 179238 489978
rect 179294 489922 179362 489978
rect 179418 489922 189834 489978
rect 189890 489922 189958 489978
rect 190014 489922 190082 489978
rect 190138 489922 190206 489978
rect 190262 489922 210518 489978
rect 210574 489922 210642 489978
rect 210698 489922 220554 489978
rect 220610 489922 220678 489978
rect 220734 489922 220802 489978
rect 220858 489922 220926 489978
rect 220982 489922 241238 489978
rect 241294 489922 241362 489978
rect 241418 489922 251274 489978
rect 251330 489922 251398 489978
rect 251454 489922 251522 489978
rect 251578 489922 251646 489978
rect 251702 489922 272518 489978
rect 272574 489922 272642 489978
rect 272698 489922 303238 489978
rect 303294 489922 303362 489978
rect 303418 489922 343434 489978
rect 343490 489922 343558 489978
rect 343614 489922 343682 489978
rect 343738 489922 343806 489978
rect 343862 489922 356518 489978
rect 356574 489922 356642 489978
rect 356698 489922 374154 489978
rect 374210 489922 374278 489978
rect 374334 489922 374402 489978
rect 374458 489922 374526 489978
rect 374582 489922 387238 489978
rect 387294 489922 387362 489978
rect 387418 489922 404874 489978
rect 404930 489922 404998 489978
rect 405054 489922 405122 489978
rect 405178 489922 405246 489978
rect 405302 489922 418518 489978
rect 418574 489922 418642 489978
rect 418698 489922 435594 489978
rect 435650 489922 435718 489978
rect 435774 489922 435842 489978
rect 435898 489922 435966 489978
rect 436022 489922 449238 489978
rect 449294 489922 449362 489978
rect 449418 489922 466314 489978
rect 466370 489922 466438 489978
rect 466494 489922 466562 489978
rect 466618 489922 466686 489978
rect 466742 489922 480518 489978
rect 480574 489922 480642 489978
rect 480698 489922 497034 489978
rect 497090 489922 497158 489978
rect 497214 489922 497282 489978
rect 497338 489922 497406 489978
rect 497462 489922 511238 489978
rect 511294 489922 511362 489978
rect 511418 489922 527754 489978
rect 527810 489922 527878 489978
rect 527934 489922 528002 489978
rect 528058 489922 528126 489978
rect 528182 489922 542518 489978
rect 542574 489922 542642 489978
rect 542698 489922 558474 489978
rect 558530 489922 558598 489978
rect 558654 489922 558722 489978
rect 558778 489922 558846 489978
rect 558902 489922 573238 489978
rect 573294 489922 573362 489978
rect 573418 489922 589194 489978
rect 589250 489922 589318 489978
rect 589374 489922 589442 489978
rect 589498 489922 589566 489978
rect 589622 489922 596496 489978
rect 596552 489922 596620 489978
rect 596676 489922 596744 489978
rect 596800 489922 596868 489978
rect 596924 489922 597980 489978
rect -1916 489826 597980 489922
rect 476012 484678 534340 484694
rect 476012 484622 476028 484678
rect 476084 484622 534268 484678
rect 534324 484622 534340 484678
rect 476012 484606 534340 484622
rect 411500 483958 473748 483974
rect 411500 483902 414652 483958
rect 414708 483902 473676 483958
rect 473732 483902 473748 483958
rect 411500 483886 473748 483902
rect 411500 483074 411588 483886
rect 78916 483058 201700 483074
rect 78916 483002 82684 483058
rect 82740 483002 141036 483058
rect 141092 483002 201628 483058
rect 201684 483002 201700 483058
rect 78916 482986 201700 483002
rect 352700 483058 411588 483074
rect 352700 483002 352716 483058
rect 352772 483002 411588 483058
rect 352700 482986 411588 483002
rect 20060 482878 20204 482894
rect 20060 482822 20076 482878
rect 20132 482822 20204 482878
rect 20060 482806 20204 482822
rect 20116 482354 20204 482806
rect 78916 482354 79004 482986
rect 20116 482266 79004 482354
rect 206652 482338 248068 482354
rect 206652 482282 206668 482338
rect 206724 482282 247996 482338
rect 248052 482282 248068 482338
rect 206652 482266 248068 482282
rect 339372 480538 472292 480554
rect 339372 480482 339388 480538
rect 339444 480482 472220 480538
rect 472276 480482 472292 480538
rect 339372 480466 472292 480482
rect 554300 480538 579700 480554
rect 554300 480482 554316 480538
rect 554372 480482 579628 480538
rect 579684 480482 579700 480538
rect 554300 480466 579700 480482
rect -1916 478350 597980 478446
rect -1916 478294 -1820 478350
rect -1764 478294 -1696 478350
rect -1640 478294 -1572 478350
rect -1516 478294 -1448 478350
rect -1392 478294 9234 478350
rect 9290 478294 9358 478350
rect 9414 478294 9482 478350
rect 9538 478294 9606 478350
rect 9662 478294 39878 478350
rect 39934 478294 40002 478350
rect 40058 478294 70674 478350
rect 70730 478294 70798 478350
rect 70854 478294 70922 478350
rect 70978 478294 71046 478350
rect 71102 478294 101878 478350
rect 101934 478294 102002 478350
rect 102058 478294 132114 478350
rect 132170 478294 132238 478350
rect 132294 478294 132362 478350
rect 132418 478294 132486 478350
rect 132542 478294 162834 478350
rect 162890 478294 162958 478350
rect 163014 478294 163082 478350
rect 163138 478294 163206 478350
rect 163262 478294 163878 478350
rect 163934 478294 164002 478350
rect 164058 478294 193554 478350
rect 193610 478294 193678 478350
rect 193734 478294 193802 478350
rect 193858 478294 193926 478350
rect 193982 478294 225878 478350
rect 225934 478294 226002 478350
rect 226058 478294 254994 478350
rect 255050 478294 255118 478350
rect 255174 478294 255242 478350
rect 255298 478294 255366 478350
rect 255422 478294 287878 478350
rect 287934 478294 288002 478350
rect 288058 478294 318598 478350
rect 318654 478294 318722 478350
rect 318778 478294 347154 478350
rect 347210 478294 347278 478350
rect 347334 478294 347402 478350
rect 347458 478294 347526 478350
rect 347582 478294 371878 478350
rect 371934 478294 372002 478350
rect 372058 478294 377874 478350
rect 377930 478294 377998 478350
rect 378054 478294 378122 478350
rect 378178 478294 378246 478350
rect 378302 478294 408594 478350
rect 408650 478294 408718 478350
rect 408774 478294 408842 478350
rect 408898 478294 408966 478350
rect 409022 478294 433878 478350
rect 433934 478294 434002 478350
rect 434058 478294 439314 478350
rect 439370 478294 439438 478350
rect 439494 478294 439562 478350
rect 439618 478294 439686 478350
rect 439742 478294 470034 478350
rect 470090 478294 470158 478350
rect 470214 478294 470282 478350
rect 470338 478294 470406 478350
rect 470462 478294 495878 478350
rect 495934 478294 496002 478350
rect 496058 478294 500754 478350
rect 500810 478294 500878 478350
rect 500934 478294 501002 478350
rect 501058 478294 501126 478350
rect 501182 478294 531474 478350
rect 531530 478294 531598 478350
rect 531654 478294 531722 478350
rect 531778 478294 531846 478350
rect 531902 478294 557878 478350
rect 557934 478294 558002 478350
rect 558058 478294 562194 478350
rect 562250 478294 562318 478350
rect 562374 478294 562442 478350
rect 562498 478294 562566 478350
rect 562622 478294 592914 478350
rect 592970 478294 593038 478350
rect 593094 478294 593162 478350
rect 593218 478294 593286 478350
rect 593342 478294 597456 478350
rect 597512 478294 597580 478350
rect 597636 478294 597704 478350
rect 597760 478294 597828 478350
rect 597884 478294 597980 478350
rect -1916 478226 597980 478294
rect -1916 478170 -1820 478226
rect -1764 478170 -1696 478226
rect -1640 478170 -1572 478226
rect -1516 478170 -1448 478226
rect -1392 478170 9234 478226
rect 9290 478170 9358 478226
rect 9414 478170 9482 478226
rect 9538 478170 9606 478226
rect 9662 478170 39878 478226
rect 39934 478170 40002 478226
rect 40058 478170 70674 478226
rect 70730 478170 70798 478226
rect 70854 478170 70922 478226
rect 70978 478170 71046 478226
rect 71102 478170 101878 478226
rect 101934 478170 102002 478226
rect 102058 478170 132114 478226
rect 132170 478170 132238 478226
rect 132294 478170 132362 478226
rect 132418 478170 132486 478226
rect 132542 478170 162834 478226
rect 162890 478170 162958 478226
rect 163014 478170 163082 478226
rect 163138 478170 163206 478226
rect 163262 478170 163878 478226
rect 163934 478170 164002 478226
rect 164058 478170 193554 478226
rect 193610 478170 193678 478226
rect 193734 478170 193802 478226
rect 193858 478170 193926 478226
rect 193982 478170 225878 478226
rect 225934 478170 226002 478226
rect 226058 478170 254994 478226
rect 255050 478170 255118 478226
rect 255174 478170 255242 478226
rect 255298 478170 255366 478226
rect 255422 478170 287878 478226
rect 287934 478170 288002 478226
rect 288058 478170 318598 478226
rect 318654 478170 318722 478226
rect 318778 478170 347154 478226
rect 347210 478170 347278 478226
rect 347334 478170 347402 478226
rect 347458 478170 347526 478226
rect 347582 478170 371878 478226
rect 371934 478170 372002 478226
rect 372058 478170 377874 478226
rect 377930 478170 377998 478226
rect 378054 478170 378122 478226
rect 378178 478170 378246 478226
rect 378302 478170 408594 478226
rect 408650 478170 408718 478226
rect 408774 478170 408842 478226
rect 408898 478170 408966 478226
rect 409022 478170 433878 478226
rect 433934 478170 434002 478226
rect 434058 478170 439314 478226
rect 439370 478170 439438 478226
rect 439494 478170 439562 478226
rect 439618 478170 439686 478226
rect 439742 478170 470034 478226
rect 470090 478170 470158 478226
rect 470214 478170 470282 478226
rect 470338 478170 470406 478226
rect 470462 478170 495878 478226
rect 495934 478170 496002 478226
rect 496058 478170 500754 478226
rect 500810 478170 500878 478226
rect 500934 478170 501002 478226
rect 501058 478170 501126 478226
rect 501182 478170 531474 478226
rect 531530 478170 531598 478226
rect 531654 478170 531722 478226
rect 531778 478170 531846 478226
rect 531902 478170 557878 478226
rect 557934 478170 558002 478226
rect 558058 478170 562194 478226
rect 562250 478170 562318 478226
rect 562374 478170 562442 478226
rect 562498 478170 562566 478226
rect 562622 478170 592914 478226
rect 592970 478170 593038 478226
rect 593094 478170 593162 478226
rect 593218 478170 593286 478226
rect 593342 478170 597456 478226
rect 597512 478170 597580 478226
rect 597636 478170 597704 478226
rect 597760 478170 597828 478226
rect 597884 478170 597980 478226
rect -1916 478102 597980 478170
rect -1916 478046 -1820 478102
rect -1764 478046 -1696 478102
rect -1640 478046 -1572 478102
rect -1516 478046 -1448 478102
rect -1392 478046 9234 478102
rect 9290 478046 9358 478102
rect 9414 478046 9482 478102
rect 9538 478046 9606 478102
rect 9662 478046 39878 478102
rect 39934 478046 40002 478102
rect 40058 478046 70674 478102
rect 70730 478046 70798 478102
rect 70854 478046 70922 478102
rect 70978 478046 71046 478102
rect 71102 478046 101878 478102
rect 101934 478046 102002 478102
rect 102058 478046 132114 478102
rect 132170 478046 132238 478102
rect 132294 478046 132362 478102
rect 132418 478046 132486 478102
rect 132542 478046 162834 478102
rect 162890 478046 162958 478102
rect 163014 478046 163082 478102
rect 163138 478046 163206 478102
rect 163262 478046 163878 478102
rect 163934 478046 164002 478102
rect 164058 478046 193554 478102
rect 193610 478046 193678 478102
rect 193734 478046 193802 478102
rect 193858 478046 193926 478102
rect 193982 478046 225878 478102
rect 225934 478046 226002 478102
rect 226058 478046 254994 478102
rect 255050 478046 255118 478102
rect 255174 478046 255242 478102
rect 255298 478046 255366 478102
rect 255422 478046 287878 478102
rect 287934 478046 288002 478102
rect 288058 478046 318598 478102
rect 318654 478046 318722 478102
rect 318778 478046 347154 478102
rect 347210 478046 347278 478102
rect 347334 478046 347402 478102
rect 347458 478046 347526 478102
rect 347582 478046 371878 478102
rect 371934 478046 372002 478102
rect 372058 478046 377874 478102
rect 377930 478046 377998 478102
rect 378054 478046 378122 478102
rect 378178 478046 378246 478102
rect 378302 478046 408594 478102
rect 408650 478046 408718 478102
rect 408774 478046 408842 478102
rect 408898 478046 408966 478102
rect 409022 478046 433878 478102
rect 433934 478046 434002 478102
rect 434058 478046 439314 478102
rect 439370 478046 439438 478102
rect 439494 478046 439562 478102
rect 439618 478046 439686 478102
rect 439742 478046 470034 478102
rect 470090 478046 470158 478102
rect 470214 478046 470282 478102
rect 470338 478046 470406 478102
rect 470462 478046 495878 478102
rect 495934 478046 496002 478102
rect 496058 478046 500754 478102
rect 500810 478046 500878 478102
rect 500934 478046 501002 478102
rect 501058 478046 501126 478102
rect 501182 478046 531474 478102
rect 531530 478046 531598 478102
rect 531654 478046 531722 478102
rect 531778 478046 531846 478102
rect 531902 478046 557878 478102
rect 557934 478046 558002 478102
rect 558058 478046 562194 478102
rect 562250 478046 562318 478102
rect 562374 478046 562442 478102
rect 562498 478046 562566 478102
rect 562622 478046 592914 478102
rect 592970 478046 593038 478102
rect 593094 478046 593162 478102
rect 593218 478046 593286 478102
rect 593342 478046 597456 478102
rect 597512 478046 597580 478102
rect 597636 478046 597704 478102
rect 597760 478046 597828 478102
rect 597884 478046 597980 478102
rect -1916 477978 597980 478046
rect -1916 477922 -1820 477978
rect -1764 477922 -1696 477978
rect -1640 477922 -1572 477978
rect -1516 477922 -1448 477978
rect -1392 477922 9234 477978
rect 9290 477922 9358 477978
rect 9414 477922 9482 477978
rect 9538 477922 9606 477978
rect 9662 477922 39878 477978
rect 39934 477922 40002 477978
rect 40058 477922 70674 477978
rect 70730 477922 70798 477978
rect 70854 477922 70922 477978
rect 70978 477922 71046 477978
rect 71102 477922 101878 477978
rect 101934 477922 102002 477978
rect 102058 477922 132114 477978
rect 132170 477922 132238 477978
rect 132294 477922 132362 477978
rect 132418 477922 132486 477978
rect 132542 477922 162834 477978
rect 162890 477922 162958 477978
rect 163014 477922 163082 477978
rect 163138 477922 163206 477978
rect 163262 477922 163878 477978
rect 163934 477922 164002 477978
rect 164058 477922 193554 477978
rect 193610 477922 193678 477978
rect 193734 477922 193802 477978
rect 193858 477922 193926 477978
rect 193982 477922 225878 477978
rect 225934 477922 226002 477978
rect 226058 477922 254994 477978
rect 255050 477922 255118 477978
rect 255174 477922 255242 477978
rect 255298 477922 255366 477978
rect 255422 477922 287878 477978
rect 287934 477922 288002 477978
rect 288058 477922 318598 477978
rect 318654 477922 318722 477978
rect 318778 477922 347154 477978
rect 347210 477922 347278 477978
rect 347334 477922 347402 477978
rect 347458 477922 347526 477978
rect 347582 477922 371878 477978
rect 371934 477922 372002 477978
rect 372058 477922 377874 477978
rect 377930 477922 377998 477978
rect 378054 477922 378122 477978
rect 378178 477922 378246 477978
rect 378302 477922 408594 477978
rect 408650 477922 408718 477978
rect 408774 477922 408842 477978
rect 408898 477922 408966 477978
rect 409022 477922 433878 477978
rect 433934 477922 434002 477978
rect 434058 477922 439314 477978
rect 439370 477922 439438 477978
rect 439494 477922 439562 477978
rect 439618 477922 439686 477978
rect 439742 477922 470034 477978
rect 470090 477922 470158 477978
rect 470214 477922 470282 477978
rect 470338 477922 470406 477978
rect 470462 477922 495878 477978
rect 495934 477922 496002 477978
rect 496058 477922 500754 477978
rect 500810 477922 500878 477978
rect 500934 477922 501002 477978
rect 501058 477922 501126 477978
rect 501182 477922 531474 477978
rect 531530 477922 531598 477978
rect 531654 477922 531722 477978
rect 531778 477922 531846 477978
rect 531902 477922 557878 477978
rect 557934 477922 558002 477978
rect 558058 477922 562194 477978
rect 562250 477922 562318 477978
rect 562374 477922 562442 477978
rect 562498 477922 562566 477978
rect 562622 477922 592914 477978
rect 592970 477922 593038 477978
rect 593094 477922 593162 477978
rect 593218 477922 593286 477978
rect 593342 477922 597456 477978
rect 597512 477922 597580 477978
rect 597636 477922 597704 477978
rect 597760 477922 597828 477978
rect 597884 477922 597980 477978
rect -1916 477826 597980 477922
rect 189516 475498 223428 475514
rect 189516 475442 189532 475498
rect 189588 475442 223428 475498
rect 189516 475426 223428 475442
rect 223340 475334 223428 475426
rect 223340 475246 231884 475334
rect 231796 474614 231884 475246
rect 206540 474598 223428 474614
rect 206540 474542 206556 474598
rect 206612 474542 223356 474598
rect 223412 474542 223428 474598
rect 206540 474526 223428 474542
rect 231796 474598 264756 474614
rect 231796 474542 264684 474598
rect 264740 474542 264756 474598
rect 231796 474526 264756 474542
rect 189516 473878 249524 473894
rect 189516 473822 189532 473878
rect 189588 473822 249452 473878
rect 249508 473822 249524 473878
rect 189516 473806 249524 473822
rect 223340 473698 263860 473714
rect 223340 473642 223356 473698
rect 223412 473642 263788 473698
rect 263844 473642 263860 473698
rect 223340 473626 263860 473642
rect 334444 473698 554388 473714
rect 334444 473642 334460 473698
rect 334516 473642 554316 473698
rect 554372 473642 554388 473698
rect 334444 473626 554388 473642
rect -1916 472350 597980 472446
rect -1916 472294 -860 472350
rect -804 472294 -736 472350
rect -680 472294 -612 472350
rect -556 472294 -488 472350
rect -432 472294 5514 472350
rect 5570 472294 5638 472350
rect 5694 472294 5762 472350
rect 5818 472294 5886 472350
rect 5942 472294 24518 472350
rect 24574 472294 24642 472350
rect 24698 472294 36234 472350
rect 36290 472294 36358 472350
rect 36414 472294 36482 472350
rect 36538 472294 36606 472350
rect 36662 472294 55238 472350
rect 55294 472294 55362 472350
rect 55418 472294 66954 472350
rect 67010 472294 67078 472350
rect 67134 472294 67202 472350
rect 67258 472294 67326 472350
rect 67382 472294 86518 472350
rect 86574 472294 86642 472350
rect 86698 472294 97674 472350
rect 97730 472294 97798 472350
rect 97854 472294 97922 472350
rect 97978 472294 98046 472350
rect 98102 472294 117238 472350
rect 117294 472294 117362 472350
rect 117418 472294 128394 472350
rect 128450 472294 128518 472350
rect 128574 472294 128642 472350
rect 128698 472294 128766 472350
rect 128822 472294 148518 472350
rect 148574 472294 148642 472350
rect 148698 472294 159114 472350
rect 159170 472294 159238 472350
rect 159294 472294 159362 472350
rect 159418 472294 159486 472350
rect 159542 472294 179238 472350
rect 179294 472294 179362 472350
rect 179418 472294 189834 472350
rect 189890 472294 189958 472350
rect 190014 472294 190082 472350
rect 190138 472294 190206 472350
rect 190262 472294 210518 472350
rect 210574 472294 210642 472350
rect 210698 472294 220554 472350
rect 220610 472294 220678 472350
rect 220734 472294 220802 472350
rect 220858 472294 220926 472350
rect 220982 472294 241238 472350
rect 241294 472294 241362 472350
rect 241418 472294 251274 472350
rect 251330 472294 251398 472350
rect 251454 472294 251522 472350
rect 251578 472294 251646 472350
rect 251702 472294 272518 472350
rect 272574 472294 272642 472350
rect 272698 472294 303238 472350
rect 303294 472294 303362 472350
rect 303418 472294 343434 472350
rect 343490 472294 343558 472350
rect 343614 472294 343682 472350
rect 343738 472294 343806 472350
rect 343862 472294 356518 472350
rect 356574 472294 356642 472350
rect 356698 472294 374154 472350
rect 374210 472294 374278 472350
rect 374334 472294 374402 472350
rect 374458 472294 374526 472350
rect 374582 472294 387238 472350
rect 387294 472294 387362 472350
rect 387418 472294 404874 472350
rect 404930 472294 404998 472350
rect 405054 472294 405122 472350
rect 405178 472294 405246 472350
rect 405302 472294 418518 472350
rect 418574 472294 418642 472350
rect 418698 472294 449238 472350
rect 449294 472294 449362 472350
rect 449418 472294 466314 472350
rect 466370 472294 466438 472350
rect 466494 472294 466562 472350
rect 466618 472294 466686 472350
rect 466742 472294 480518 472350
rect 480574 472294 480642 472350
rect 480698 472294 511238 472350
rect 511294 472294 511362 472350
rect 511418 472294 527754 472350
rect 527810 472294 527878 472350
rect 527934 472294 528002 472350
rect 528058 472294 528126 472350
rect 528182 472294 542518 472350
rect 542574 472294 542642 472350
rect 542698 472294 573238 472350
rect 573294 472294 573362 472350
rect 573418 472294 589194 472350
rect 589250 472294 589318 472350
rect 589374 472294 589442 472350
rect 589498 472294 589566 472350
rect 589622 472294 596496 472350
rect 596552 472294 596620 472350
rect 596676 472294 596744 472350
rect 596800 472294 596868 472350
rect 596924 472294 597980 472350
rect -1916 472226 597980 472294
rect -1916 472170 -860 472226
rect -804 472170 -736 472226
rect -680 472170 -612 472226
rect -556 472170 -488 472226
rect -432 472170 5514 472226
rect 5570 472170 5638 472226
rect 5694 472170 5762 472226
rect 5818 472170 5886 472226
rect 5942 472170 24518 472226
rect 24574 472170 24642 472226
rect 24698 472170 36234 472226
rect 36290 472170 36358 472226
rect 36414 472170 36482 472226
rect 36538 472170 36606 472226
rect 36662 472170 55238 472226
rect 55294 472170 55362 472226
rect 55418 472170 66954 472226
rect 67010 472170 67078 472226
rect 67134 472170 67202 472226
rect 67258 472170 67326 472226
rect 67382 472170 86518 472226
rect 86574 472170 86642 472226
rect 86698 472170 97674 472226
rect 97730 472170 97798 472226
rect 97854 472170 97922 472226
rect 97978 472170 98046 472226
rect 98102 472170 117238 472226
rect 117294 472170 117362 472226
rect 117418 472170 128394 472226
rect 128450 472170 128518 472226
rect 128574 472170 128642 472226
rect 128698 472170 128766 472226
rect 128822 472170 148518 472226
rect 148574 472170 148642 472226
rect 148698 472170 159114 472226
rect 159170 472170 159238 472226
rect 159294 472170 159362 472226
rect 159418 472170 159486 472226
rect 159542 472170 179238 472226
rect 179294 472170 179362 472226
rect 179418 472170 189834 472226
rect 189890 472170 189958 472226
rect 190014 472170 190082 472226
rect 190138 472170 190206 472226
rect 190262 472170 210518 472226
rect 210574 472170 210642 472226
rect 210698 472170 220554 472226
rect 220610 472170 220678 472226
rect 220734 472170 220802 472226
rect 220858 472170 220926 472226
rect 220982 472170 241238 472226
rect 241294 472170 241362 472226
rect 241418 472170 251274 472226
rect 251330 472170 251398 472226
rect 251454 472170 251522 472226
rect 251578 472170 251646 472226
rect 251702 472170 272518 472226
rect 272574 472170 272642 472226
rect 272698 472170 303238 472226
rect 303294 472170 303362 472226
rect 303418 472170 343434 472226
rect 343490 472170 343558 472226
rect 343614 472170 343682 472226
rect 343738 472170 343806 472226
rect 343862 472170 356518 472226
rect 356574 472170 356642 472226
rect 356698 472170 374154 472226
rect 374210 472170 374278 472226
rect 374334 472170 374402 472226
rect 374458 472170 374526 472226
rect 374582 472170 387238 472226
rect 387294 472170 387362 472226
rect 387418 472170 404874 472226
rect 404930 472170 404998 472226
rect 405054 472170 405122 472226
rect 405178 472170 405246 472226
rect 405302 472170 418518 472226
rect 418574 472170 418642 472226
rect 418698 472170 449238 472226
rect 449294 472170 449362 472226
rect 449418 472170 466314 472226
rect 466370 472170 466438 472226
rect 466494 472170 466562 472226
rect 466618 472170 466686 472226
rect 466742 472170 480518 472226
rect 480574 472170 480642 472226
rect 480698 472170 511238 472226
rect 511294 472170 511362 472226
rect 511418 472170 527754 472226
rect 527810 472170 527878 472226
rect 527934 472170 528002 472226
rect 528058 472170 528126 472226
rect 528182 472170 542518 472226
rect 542574 472170 542642 472226
rect 542698 472170 573238 472226
rect 573294 472170 573362 472226
rect 573418 472170 589194 472226
rect 589250 472170 589318 472226
rect 589374 472170 589442 472226
rect 589498 472170 589566 472226
rect 589622 472170 596496 472226
rect 596552 472170 596620 472226
rect 596676 472170 596744 472226
rect 596800 472170 596868 472226
rect 596924 472170 597980 472226
rect -1916 472102 597980 472170
rect -1916 472046 -860 472102
rect -804 472046 -736 472102
rect -680 472046 -612 472102
rect -556 472046 -488 472102
rect -432 472046 5514 472102
rect 5570 472046 5638 472102
rect 5694 472046 5762 472102
rect 5818 472046 5886 472102
rect 5942 472046 24518 472102
rect 24574 472046 24642 472102
rect 24698 472046 36234 472102
rect 36290 472046 36358 472102
rect 36414 472046 36482 472102
rect 36538 472046 36606 472102
rect 36662 472046 55238 472102
rect 55294 472046 55362 472102
rect 55418 472046 66954 472102
rect 67010 472046 67078 472102
rect 67134 472046 67202 472102
rect 67258 472046 67326 472102
rect 67382 472046 86518 472102
rect 86574 472046 86642 472102
rect 86698 472046 97674 472102
rect 97730 472046 97798 472102
rect 97854 472046 97922 472102
rect 97978 472046 98046 472102
rect 98102 472046 117238 472102
rect 117294 472046 117362 472102
rect 117418 472046 128394 472102
rect 128450 472046 128518 472102
rect 128574 472046 128642 472102
rect 128698 472046 128766 472102
rect 128822 472046 148518 472102
rect 148574 472046 148642 472102
rect 148698 472046 159114 472102
rect 159170 472046 159238 472102
rect 159294 472046 159362 472102
rect 159418 472046 159486 472102
rect 159542 472046 179238 472102
rect 179294 472046 179362 472102
rect 179418 472046 189834 472102
rect 189890 472046 189958 472102
rect 190014 472046 190082 472102
rect 190138 472046 190206 472102
rect 190262 472046 210518 472102
rect 210574 472046 210642 472102
rect 210698 472046 220554 472102
rect 220610 472046 220678 472102
rect 220734 472046 220802 472102
rect 220858 472046 220926 472102
rect 220982 472046 241238 472102
rect 241294 472046 241362 472102
rect 241418 472046 251274 472102
rect 251330 472046 251398 472102
rect 251454 472046 251522 472102
rect 251578 472046 251646 472102
rect 251702 472046 272518 472102
rect 272574 472046 272642 472102
rect 272698 472046 303238 472102
rect 303294 472046 303362 472102
rect 303418 472046 343434 472102
rect 343490 472046 343558 472102
rect 343614 472046 343682 472102
rect 343738 472046 343806 472102
rect 343862 472046 356518 472102
rect 356574 472046 356642 472102
rect 356698 472046 374154 472102
rect 374210 472046 374278 472102
rect 374334 472046 374402 472102
rect 374458 472046 374526 472102
rect 374582 472046 387238 472102
rect 387294 472046 387362 472102
rect 387418 472046 404874 472102
rect 404930 472046 404998 472102
rect 405054 472046 405122 472102
rect 405178 472046 405246 472102
rect 405302 472046 418518 472102
rect 418574 472046 418642 472102
rect 418698 472060 449238 472102
rect 418698 472046 435594 472060
rect -1916 472004 435594 472046
rect 435650 472004 435718 472060
rect 435774 472004 435842 472060
rect 435898 472004 435966 472060
rect 436022 472046 449238 472060
rect 449294 472046 449362 472102
rect 449418 472046 466314 472102
rect 466370 472046 466438 472102
rect 466494 472046 466562 472102
rect 466618 472046 466686 472102
rect 466742 472046 480518 472102
rect 480574 472046 480642 472102
rect 480698 472046 511238 472102
rect 511294 472046 511362 472102
rect 511418 472046 527754 472102
rect 527810 472046 527878 472102
rect 527934 472046 528002 472102
rect 528058 472046 528126 472102
rect 528182 472046 542518 472102
rect 542574 472046 542642 472102
rect 542698 472046 573238 472102
rect 573294 472046 573362 472102
rect 573418 472046 589194 472102
rect 589250 472046 589318 472102
rect 589374 472046 589442 472102
rect 589498 472046 589566 472102
rect 589622 472046 596496 472102
rect 596552 472046 596620 472102
rect 596676 472046 596744 472102
rect 596800 472046 596868 472102
rect 596924 472046 597980 472102
rect 436022 472004 597980 472046
rect -1916 471978 597980 472004
rect -1916 471922 -860 471978
rect -804 471922 -736 471978
rect -680 471922 -612 471978
rect -556 471922 -488 471978
rect -432 471922 5514 471978
rect 5570 471922 5638 471978
rect 5694 471922 5762 471978
rect 5818 471922 5886 471978
rect 5942 471922 24518 471978
rect 24574 471922 24642 471978
rect 24698 471922 36234 471978
rect 36290 471922 36358 471978
rect 36414 471922 36482 471978
rect 36538 471922 36606 471978
rect 36662 471922 55238 471978
rect 55294 471922 55362 471978
rect 55418 471922 66954 471978
rect 67010 471922 67078 471978
rect 67134 471922 67202 471978
rect 67258 471922 67326 471978
rect 67382 471922 86518 471978
rect 86574 471922 86642 471978
rect 86698 471922 97674 471978
rect 97730 471922 97798 471978
rect 97854 471922 97922 471978
rect 97978 471922 98046 471978
rect 98102 471922 117238 471978
rect 117294 471922 117362 471978
rect 117418 471922 128394 471978
rect 128450 471922 128518 471978
rect 128574 471922 128642 471978
rect 128698 471922 128766 471978
rect 128822 471922 148518 471978
rect 148574 471922 148642 471978
rect 148698 471922 159114 471978
rect 159170 471922 159238 471978
rect 159294 471922 159362 471978
rect 159418 471922 159486 471978
rect 159542 471922 179238 471978
rect 179294 471922 179362 471978
rect 179418 471922 189834 471978
rect 189890 471922 189958 471978
rect 190014 471922 190082 471978
rect 190138 471922 190206 471978
rect 190262 471922 210518 471978
rect 210574 471922 210642 471978
rect 210698 471922 220554 471978
rect 220610 471922 220678 471978
rect 220734 471922 220802 471978
rect 220858 471922 220926 471978
rect 220982 471922 241238 471978
rect 241294 471922 241362 471978
rect 241418 471922 251274 471978
rect 251330 471922 251398 471978
rect 251454 471922 251522 471978
rect 251578 471922 251646 471978
rect 251702 471922 272518 471978
rect 272574 471922 272642 471978
rect 272698 471922 303238 471978
rect 303294 471922 303362 471978
rect 303418 471922 343434 471978
rect 343490 471922 343558 471978
rect 343614 471922 343682 471978
rect 343738 471922 343806 471978
rect 343862 471922 356518 471978
rect 356574 471922 356642 471978
rect 356698 471922 374154 471978
rect 374210 471922 374278 471978
rect 374334 471922 374402 471978
rect 374458 471922 374526 471978
rect 374582 471922 387238 471978
rect 387294 471922 387362 471978
rect 387418 471922 404874 471978
rect 404930 471922 404998 471978
rect 405054 471922 405122 471978
rect 405178 471922 405246 471978
rect 405302 471922 418518 471978
rect 418574 471922 418642 471978
rect 418698 471936 449238 471978
rect 418698 471922 435594 471936
rect -1916 471880 435594 471922
rect 435650 471880 435718 471936
rect 435774 471880 435842 471936
rect 435898 471880 435966 471936
rect 436022 471922 449238 471936
rect 449294 471922 449362 471978
rect 449418 471922 466314 471978
rect 466370 471922 466438 471978
rect 466494 471922 466562 471978
rect 466618 471922 466686 471978
rect 466742 471922 480518 471978
rect 480574 471922 480642 471978
rect 480698 471922 511238 471978
rect 511294 471922 511362 471978
rect 511418 471922 527754 471978
rect 527810 471922 527878 471978
rect 527934 471922 528002 471978
rect 528058 471922 528126 471978
rect 528182 471922 542518 471978
rect 542574 471922 542642 471978
rect 542698 471922 573238 471978
rect 573294 471922 573362 471978
rect 573418 471922 589194 471978
rect 589250 471922 589318 471978
rect 589374 471922 589442 471978
rect 589498 471922 589566 471978
rect 589622 471922 596496 471978
rect 596552 471922 596620 471978
rect 596676 471922 596744 471978
rect 596800 471922 596868 471978
rect 596924 471922 597980 471978
rect 436022 471880 597980 471922
rect -1916 471826 597980 471880
rect 334444 470638 554388 470654
rect 334444 470582 334460 470638
rect 334516 470582 554388 470638
rect 334444 470566 554388 470582
rect 334444 470458 554164 470474
rect 334444 470402 334460 470458
rect 334516 470402 554092 470458
rect 554148 470402 554164 470458
rect 334444 470386 554164 470402
rect 554300 470294 554388 470566
rect 554300 470278 583060 470294
rect 554300 470222 582988 470278
rect 583044 470222 583060 470278
rect 554300 470206 583060 470222
rect 572836 469918 579364 469934
rect 572836 469862 579292 469918
rect 579348 469862 579364 469918
rect 572836 469846 579364 469862
rect 572836 469574 572924 469846
rect 144380 469558 193188 469574
rect 144380 469502 144396 469558
rect 144452 469502 193116 469558
rect 193172 469502 193188 469558
rect 144380 469486 193188 469502
rect 197356 469558 264196 469574
rect 197356 469502 197372 469558
rect 197428 469502 264124 469558
rect 264180 469502 264196 469558
rect 197356 469486 264196 469502
rect 334444 469558 572924 469574
rect 334444 469502 334460 469558
rect 334516 469502 572924 469558
rect 334444 469486 572924 469502
rect 351020 468658 579476 468674
rect 351020 468602 351036 468658
rect 351092 468602 579404 468658
rect 579460 468602 579476 468658
rect 351020 468586 579476 468602
rect 579612 468658 579700 468674
rect 579612 468602 579628 468658
rect 579684 468602 579700 468658
rect 579612 468494 579700 468602
rect 554076 468478 579700 468494
rect 554076 468422 554092 468478
rect 554148 468422 579700 468478
rect 554076 468406 579700 468422
rect 194892 467938 264084 467954
rect 194892 467882 194908 467938
rect 194964 467882 264012 467938
rect 264068 467882 264084 467938
rect 194892 467866 264084 467882
rect 140908 466138 249636 466154
rect 140908 466082 140924 466138
rect 140980 466082 249564 466138
rect 249620 466082 249636 466138
rect 140908 466066 249636 466082
rect 334444 466138 521124 466154
rect 334444 466082 334460 466138
rect 334516 466082 521052 466138
rect 521108 466082 521124 466138
rect 334444 466066 521124 466082
rect 193100 465238 263860 465254
rect 193100 465182 193116 465238
rect 193172 465182 263788 465238
rect 263844 465182 263860 465238
rect 193100 465166 263860 465182
rect 334444 465238 473188 465254
rect 334444 465182 334460 465238
rect 334516 465182 473116 465238
rect 473172 465182 473188 465238
rect 334444 465166 473188 465182
rect 199036 463618 263860 463634
rect 199036 463562 199052 463618
rect 199108 463562 263788 463618
rect 263844 463562 263860 463618
rect 199036 463546 263860 463562
rect 334444 462898 462884 462914
rect 334444 462842 334460 462898
rect 334516 462842 462812 462898
rect 462868 462842 462884 462898
rect 334444 462826 462884 462842
rect -1916 460350 597980 460446
rect -1916 460294 -1820 460350
rect -1764 460294 -1696 460350
rect -1640 460294 -1572 460350
rect -1516 460294 -1448 460350
rect -1392 460294 9234 460350
rect 9290 460294 9358 460350
rect 9414 460294 9482 460350
rect 9538 460294 9606 460350
rect 9662 460294 39878 460350
rect 39934 460294 40002 460350
rect 40058 460294 70674 460350
rect 70730 460294 70798 460350
rect 70854 460294 70922 460350
rect 70978 460294 71046 460350
rect 71102 460294 101878 460350
rect 101934 460294 102002 460350
rect 102058 460294 132114 460350
rect 132170 460294 132238 460350
rect 132294 460294 132362 460350
rect 132418 460294 132486 460350
rect 132542 460294 162834 460350
rect 162890 460294 162958 460350
rect 163014 460294 163082 460350
rect 163138 460294 163206 460350
rect 163262 460294 163878 460350
rect 163934 460294 164002 460350
rect 164058 460294 193554 460350
rect 193610 460294 193678 460350
rect 193734 460294 193802 460350
rect 193858 460294 193926 460350
rect 193982 460294 224274 460350
rect 224330 460294 224398 460350
rect 224454 460294 224522 460350
rect 224578 460294 224646 460350
rect 224702 460294 225878 460350
rect 225934 460294 226002 460350
rect 226058 460294 254994 460350
rect 255050 460294 255118 460350
rect 255174 460294 255242 460350
rect 255298 460294 255366 460350
rect 255422 460294 287878 460350
rect 287934 460294 288002 460350
rect 288058 460294 318598 460350
rect 318654 460294 318722 460350
rect 318778 460294 347154 460350
rect 347210 460294 347278 460350
rect 347334 460294 347402 460350
rect 347458 460294 347526 460350
rect 347582 460294 371878 460350
rect 371934 460294 372002 460350
rect 372058 460294 377874 460350
rect 377930 460294 377998 460350
rect 378054 460294 378122 460350
rect 378178 460294 378246 460350
rect 378302 460294 408594 460350
rect 408650 460294 408718 460350
rect 408774 460294 408842 460350
rect 408898 460294 408966 460350
rect 409022 460294 433878 460350
rect 433934 460294 434002 460350
rect 434058 460294 439314 460350
rect 439370 460294 439438 460350
rect 439494 460294 439562 460350
rect 439618 460294 439686 460350
rect 439742 460294 470034 460350
rect 470090 460294 470158 460350
rect 470214 460294 470282 460350
rect 470338 460294 470406 460350
rect 470462 460294 495878 460350
rect 495934 460294 496002 460350
rect 496058 460294 500754 460350
rect 500810 460294 500878 460350
rect 500934 460294 501002 460350
rect 501058 460294 501126 460350
rect 501182 460294 531474 460350
rect 531530 460294 531598 460350
rect 531654 460294 531722 460350
rect 531778 460294 531846 460350
rect 531902 460294 557878 460350
rect 557934 460294 558002 460350
rect 558058 460294 562194 460350
rect 562250 460294 562318 460350
rect 562374 460294 562442 460350
rect 562498 460294 562566 460350
rect 562622 460294 592914 460350
rect 592970 460294 593038 460350
rect 593094 460294 593162 460350
rect 593218 460294 593286 460350
rect 593342 460294 597456 460350
rect 597512 460294 597580 460350
rect 597636 460294 597704 460350
rect 597760 460294 597828 460350
rect 597884 460294 597980 460350
rect -1916 460226 597980 460294
rect -1916 460170 -1820 460226
rect -1764 460170 -1696 460226
rect -1640 460170 -1572 460226
rect -1516 460170 -1448 460226
rect -1392 460170 9234 460226
rect 9290 460170 9358 460226
rect 9414 460170 9482 460226
rect 9538 460170 9606 460226
rect 9662 460170 39878 460226
rect 39934 460170 40002 460226
rect 40058 460170 70674 460226
rect 70730 460170 70798 460226
rect 70854 460170 70922 460226
rect 70978 460170 71046 460226
rect 71102 460170 101878 460226
rect 101934 460170 102002 460226
rect 102058 460170 132114 460226
rect 132170 460170 132238 460226
rect 132294 460170 132362 460226
rect 132418 460170 132486 460226
rect 132542 460170 162834 460226
rect 162890 460170 162958 460226
rect 163014 460170 163082 460226
rect 163138 460170 163206 460226
rect 163262 460170 163878 460226
rect 163934 460170 164002 460226
rect 164058 460170 193554 460226
rect 193610 460170 193678 460226
rect 193734 460170 193802 460226
rect 193858 460170 193926 460226
rect 193982 460170 224274 460226
rect 224330 460170 224398 460226
rect 224454 460170 224522 460226
rect 224578 460170 224646 460226
rect 224702 460170 225878 460226
rect 225934 460170 226002 460226
rect 226058 460170 254994 460226
rect 255050 460170 255118 460226
rect 255174 460170 255242 460226
rect 255298 460170 255366 460226
rect 255422 460170 287878 460226
rect 287934 460170 288002 460226
rect 288058 460170 318598 460226
rect 318654 460170 318722 460226
rect 318778 460170 347154 460226
rect 347210 460170 347278 460226
rect 347334 460170 347402 460226
rect 347458 460170 347526 460226
rect 347582 460170 371878 460226
rect 371934 460170 372002 460226
rect 372058 460170 377874 460226
rect 377930 460170 377998 460226
rect 378054 460170 378122 460226
rect 378178 460170 378246 460226
rect 378302 460170 408594 460226
rect 408650 460170 408718 460226
rect 408774 460170 408842 460226
rect 408898 460170 408966 460226
rect 409022 460170 433878 460226
rect 433934 460170 434002 460226
rect 434058 460170 439314 460226
rect 439370 460170 439438 460226
rect 439494 460170 439562 460226
rect 439618 460170 439686 460226
rect 439742 460170 470034 460226
rect 470090 460170 470158 460226
rect 470214 460170 470282 460226
rect 470338 460170 470406 460226
rect 470462 460170 495878 460226
rect 495934 460170 496002 460226
rect 496058 460170 500754 460226
rect 500810 460170 500878 460226
rect 500934 460170 501002 460226
rect 501058 460170 501126 460226
rect 501182 460170 531474 460226
rect 531530 460170 531598 460226
rect 531654 460170 531722 460226
rect 531778 460170 531846 460226
rect 531902 460170 557878 460226
rect 557934 460170 558002 460226
rect 558058 460170 562194 460226
rect 562250 460170 562318 460226
rect 562374 460170 562442 460226
rect 562498 460170 562566 460226
rect 562622 460170 592914 460226
rect 592970 460170 593038 460226
rect 593094 460170 593162 460226
rect 593218 460170 593286 460226
rect 593342 460170 597456 460226
rect 597512 460170 597580 460226
rect 597636 460170 597704 460226
rect 597760 460170 597828 460226
rect 597884 460170 597980 460226
rect -1916 460102 597980 460170
rect -1916 460046 -1820 460102
rect -1764 460046 -1696 460102
rect -1640 460046 -1572 460102
rect -1516 460046 -1448 460102
rect -1392 460046 9234 460102
rect 9290 460046 9358 460102
rect 9414 460046 9482 460102
rect 9538 460046 9606 460102
rect 9662 460046 39878 460102
rect 39934 460046 40002 460102
rect 40058 460046 70674 460102
rect 70730 460046 70798 460102
rect 70854 460046 70922 460102
rect 70978 460046 71046 460102
rect 71102 460046 101878 460102
rect 101934 460046 102002 460102
rect 102058 460046 132114 460102
rect 132170 460046 132238 460102
rect 132294 460046 132362 460102
rect 132418 460046 132486 460102
rect 132542 460046 162834 460102
rect 162890 460046 162958 460102
rect 163014 460046 163082 460102
rect 163138 460046 163206 460102
rect 163262 460046 163878 460102
rect 163934 460046 164002 460102
rect 164058 460046 193554 460102
rect 193610 460046 193678 460102
rect 193734 460046 193802 460102
rect 193858 460046 193926 460102
rect 193982 460046 224274 460102
rect 224330 460046 224398 460102
rect 224454 460046 224522 460102
rect 224578 460046 224646 460102
rect 224702 460046 225878 460102
rect 225934 460046 226002 460102
rect 226058 460046 254994 460102
rect 255050 460046 255118 460102
rect 255174 460046 255242 460102
rect 255298 460046 255366 460102
rect 255422 460046 287878 460102
rect 287934 460046 288002 460102
rect 288058 460046 318598 460102
rect 318654 460046 318722 460102
rect 318778 460046 347154 460102
rect 347210 460046 347278 460102
rect 347334 460046 347402 460102
rect 347458 460046 347526 460102
rect 347582 460046 371878 460102
rect 371934 460046 372002 460102
rect 372058 460046 377874 460102
rect 377930 460046 377998 460102
rect 378054 460046 378122 460102
rect 378178 460046 378246 460102
rect 378302 460046 408594 460102
rect 408650 460046 408718 460102
rect 408774 460046 408842 460102
rect 408898 460046 408966 460102
rect 409022 460046 433878 460102
rect 433934 460046 434002 460102
rect 434058 460046 439314 460102
rect 439370 460046 439438 460102
rect 439494 460046 439562 460102
rect 439618 460046 439686 460102
rect 439742 460046 470034 460102
rect 470090 460046 470158 460102
rect 470214 460046 470282 460102
rect 470338 460046 470406 460102
rect 470462 460046 495878 460102
rect 495934 460046 496002 460102
rect 496058 460046 500754 460102
rect 500810 460046 500878 460102
rect 500934 460046 501002 460102
rect 501058 460046 501126 460102
rect 501182 460046 531474 460102
rect 531530 460046 531598 460102
rect 531654 460046 531722 460102
rect 531778 460046 531846 460102
rect 531902 460046 557878 460102
rect 557934 460046 558002 460102
rect 558058 460046 562194 460102
rect 562250 460046 562318 460102
rect 562374 460046 562442 460102
rect 562498 460046 562566 460102
rect 562622 460046 592914 460102
rect 592970 460046 593038 460102
rect 593094 460046 593162 460102
rect 593218 460046 593286 460102
rect 593342 460046 597456 460102
rect 597512 460046 597580 460102
rect 597636 460046 597704 460102
rect 597760 460046 597828 460102
rect 597884 460046 597980 460102
rect -1916 459978 597980 460046
rect -1916 459922 -1820 459978
rect -1764 459922 -1696 459978
rect -1640 459922 -1572 459978
rect -1516 459922 -1448 459978
rect -1392 459922 9234 459978
rect 9290 459922 9358 459978
rect 9414 459922 9482 459978
rect 9538 459922 9606 459978
rect 9662 459922 39878 459978
rect 39934 459922 40002 459978
rect 40058 459922 70674 459978
rect 70730 459922 70798 459978
rect 70854 459922 70922 459978
rect 70978 459922 71046 459978
rect 71102 459922 101878 459978
rect 101934 459922 102002 459978
rect 102058 459922 132114 459978
rect 132170 459922 132238 459978
rect 132294 459922 132362 459978
rect 132418 459922 132486 459978
rect 132542 459922 162834 459978
rect 162890 459922 162958 459978
rect 163014 459922 163082 459978
rect 163138 459922 163206 459978
rect 163262 459922 163878 459978
rect 163934 459922 164002 459978
rect 164058 459922 193554 459978
rect 193610 459922 193678 459978
rect 193734 459922 193802 459978
rect 193858 459922 193926 459978
rect 193982 459922 224274 459978
rect 224330 459922 224398 459978
rect 224454 459922 224522 459978
rect 224578 459922 224646 459978
rect 224702 459922 225878 459978
rect 225934 459922 226002 459978
rect 226058 459922 254994 459978
rect 255050 459922 255118 459978
rect 255174 459922 255242 459978
rect 255298 459922 255366 459978
rect 255422 459922 287878 459978
rect 287934 459922 288002 459978
rect 288058 459922 318598 459978
rect 318654 459922 318722 459978
rect 318778 459922 347154 459978
rect 347210 459922 347278 459978
rect 347334 459922 347402 459978
rect 347458 459922 347526 459978
rect 347582 459922 371878 459978
rect 371934 459922 372002 459978
rect 372058 459922 377874 459978
rect 377930 459922 377998 459978
rect 378054 459922 378122 459978
rect 378178 459922 378246 459978
rect 378302 459922 408594 459978
rect 408650 459922 408718 459978
rect 408774 459922 408842 459978
rect 408898 459922 408966 459978
rect 409022 459922 433878 459978
rect 433934 459922 434002 459978
rect 434058 459922 439314 459978
rect 439370 459922 439438 459978
rect 439494 459922 439562 459978
rect 439618 459922 439686 459978
rect 439742 459922 470034 459978
rect 470090 459922 470158 459978
rect 470214 459922 470282 459978
rect 470338 459922 470406 459978
rect 470462 459922 495878 459978
rect 495934 459922 496002 459978
rect 496058 459922 500754 459978
rect 500810 459922 500878 459978
rect 500934 459922 501002 459978
rect 501058 459922 501126 459978
rect 501182 459922 531474 459978
rect 531530 459922 531598 459978
rect 531654 459922 531722 459978
rect 531778 459922 531846 459978
rect 531902 459922 557878 459978
rect 557934 459922 558002 459978
rect 558058 459922 562194 459978
rect 562250 459922 562318 459978
rect 562374 459922 562442 459978
rect 562498 459922 562566 459978
rect 562622 459922 592914 459978
rect 592970 459922 593038 459978
rect 593094 459922 593162 459978
rect 593218 459922 593286 459978
rect 593342 459922 597456 459978
rect 597512 459922 597580 459978
rect 597636 459922 597704 459978
rect 597760 459922 597828 459978
rect 597884 459922 597980 459978
rect -1916 459826 597980 459922
rect -1916 454350 597980 454446
rect -1916 454294 -860 454350
rect -804 454294 -736 454350
rect -680 454294 -612 454350
rect -556 454294 -488 454350
rect -432 454294 5514 454350
rect 5570 454294 5638 454350
rect 5694 454294 5762 454350
rect 5818 454294 5886 454350
rect 5942 454294 36234 454350
rect 36290 454294 36358 454350
rect 36414 454294 36482 454350
rect 36538 454294 36606 454350
rect 36662 454294 66954 454350
rect 67010 454294 67078 454350
rect 67134 454294 67202 454350
rect 67258 454294 67326 454350
rect 67382 454294 97674 454350
rect 97730 454294 97798 454350
rect 97854 454294 97922 454350
rect 97978 454294 98046 454350
rect 98102 454294 128394 454350
rect 128450 454294 128518 454350
rect 128574 454294 128642 454350
rect 128698 454294 128766 454350
rect 128822 454294 159114 454350
rect 159170 454294 159238 454350
rect 159294 454294 159362 454350
rect 159418 454294 159486 454350
rect 159542 454294 189834 454350
rect 189890 454294 189958 454350
rect 190014 454294 190082 454350
rect 190138 454294 190206 454350
rect 190262 454294 220554 454350
rect 220610 454294 220678 454350
rect 220734 454294 220802 454350
rect 220858 454294 220926 454350
rect 220982 454294 251274 454350
rect 251330 454294 251398 454350
rect 251454 454294 251522 454350
rect 251578 454294 251646 454350
rect 251702 454294 272518 454350
rect 272574 454294 272642 454350
rect 272698 454294 303238 454350
rect 303294 454294 303362 454350
rect 303418 454294 343434 454350
rect 343490 454294 343558 454350
rect 343614 454294 343682 454350
rect 343738 454294 343806 454350
rect 343862 454294 374154 454350
rect 374210 454294 374278 454350
rect 374334 454294 374402 454350
rect 374458 454294 374526 454350
rect 374582 454294 404874 454350
rect 404930 454294 404998 454350
rect 405054 454294 405122 454350
rect 405178 454294 405246 454350
rect 405302 454294 435594 454350
rect 435650 454294 435718 454350
rect 435774 454294 435842 454350
rect 435898 454294 435966 454350
rect 436022 454294 466314 454350
rect 466370 454294 466438 454350
rect 466494 454294 466562 454350
rect 466618 454294 466686 454350
rect 466742 454294 497034 454350
rect 497090 454294 497158 454350
rect 497214 454294 497282 454350
rect 497338 454294 497406 454350
rect 497462 454294 527754 454350
rect 527810 454294 527878 454350
rect 527934 454294 528002 454350
rect 528058 454294 528126 454350
rect 528182 454294 558474 454350
rect 558530 454294 558598 454350
rect 558654 454294 558722 454350
rect 558778 454294 558846 454350
rect 558902 454294 589194 454350
rect 589250 454294 589318 454350
rect 589374 454294 589442 454350
rect 589498 454294 589566 454350
rect 589622 454294 596496 454350
rect 596552 454294 596620 454350
rect 596676 454294 596744 454350
rect 596800 454294 596868 454350
rect 596924 454294 597980 454350
rect -1916 454226 597980 454294
rect -1916 454170 -860 454226
rect -804 454170 -736 454226
rect -680 454170 -612 454226
rect -556 454170 -488 454226
rect -432 454170 5514 454226
rect 5570 454170 5638 454226
rect 5694 454170 5762 454226
rect 5818 454170 5886 454226
rect 5942 454170 36234 454226
rect 36290 454170 36358 454226
rect 36414 454170 36482 454226
rect 36538 454170 36606 454226
rect 36662 454170 66954 454226
rect 67010 454170 67078 454226
rect 67134 454170 67202 454226
rect 67258 454170 67326 454226
rect 67382 454170 97674 454226
rect 97730 454170 97798 454226
rect 97854 454170 97922 454226
rect 97978 454170 98046 454226
rect 98102 454170 128394 454226
rect 128450 454170 128518 454226
rect 128574 454170 128642 454226
rect 128698 454170 128766 454226
rect 128822 454170 159114 454226
rect 159170 454170 159238 454226
rect 159294 454170 159362 454226
rect 159418 454170 159486 454226
rect 159542 454170 189834 454226
rect 189890 454170 189958 454226
rect 190014 454170 190082 454226
rect 190138 454170 190206 454226
rect 190262 454170 220554 454226
rect 220610 454170 220678 454226
rect 220734 454170 220802 454226
rect 220858 454170 220926 454226
rect 220982 454170 251274 454226
rect 251330 454170 251398 454226
rect 251454 454170 251522 454226
rect 251578 454170 251646 454226
rect 251702 454170 272518 454226
rect 272574 454170 272642 454226
rect 272698 454170 303238 454226
rect 303294 454170 303362 454226
rect 303418 454170 343434 454226
rect 343490 454170 343558 454226
rect 343614 454170 343682 454226
rect 343738 454170 343806 454226
rect 343862 454170 374154 454226
rect 374210 454170 374278 454226
rect 374334 454170 374402 454226
rect 374458 454170 374526 454226
rect 374582 454170 404874 454226
rect 404930 454170 404998 454226
rect 405054 454170 405122 454226
rect 405178 454170 405246 454226
rect 405302 454170 435594 454226
rect 435650 454170 435718 454226
rect 435774 454170 435842 454226
rect 435898 454170 435966 454226
rect 436022 454170 466314 454226
rect 466370 454170 466438 454226
rect 466494 454170 466562 454226
rect 466618 454170 466686 454226
rect 466742 454170 497034 454226
rect 497090 454170 497158 454226
rect 497214 454170 497282 454226
rect 497338 454170 497406 454226
rect 497462 454170 527754 454226
rect 527810 454170 527878 454226
rect 527934 454170 528002 454226
rect 528058 454170 528126 454226
rect 528182 454170 558474 454226
rect 558530 454170 558598 454226
rect 558654 454170 558722 454226
rect 558778 454170 558846 454226
rect 558902 454170 589194 454226
rect 589250 454170 589318 454226
rect 589374 454170 589442 454226
rect 589498 454170 589566 454226
rect 589622 454170 596496 454226
rect 596552 454170 596620 454226
rect 596676 454170 596744 454226
rect 596800 454170 596868 454226
rect 596924 454170 597980 454226
rect -1916 454102 597980 454170
rect -1916 454046 -860 454102
rect -804 454046 -736 454102
rect -680 454046 -612 454102
rect -556 454046 -488 454102
rect -432 454046 5514 454102
rect 5570 454046 5638 454102
rect 5694 454046 5762 454102
rect 5818 454046 5886 454102
rect 5942 454046 36234 454102
rect 36290 454046 36358 454102
rect 36414 454046 36482 454102
rect 36538 454046 36606 454102
rect 36662 454046 66954 454102
rect 67010 454046 67078 454102
rect 67134 454046 67202 454102
rect 67258 454046 67326 454102
rect 67382 454046 97674 454102
rect 97730 454046 97798 454102
rect 97854 454046 97922 454102
rect 97978 454046 98046 454102
rect 98102 454046 128394 454102
rect 128450 454046 128518 454102
rect 128574 454046 128642 454102
rect 128698 454046 128766 454102
rect 128822 454046 159114 454102
rect 159170 454046 159238 454102
rect 159294 454046 159362 454102
rect 159418 454046 159486 454102
rect 159542 454046 189834 454102
rect 189890 454046 189958 454102
rect 190014 454046 190082 454102
rect 190138 454046 190206 454102
rect 190262 454046 220554 454102
rect 220610 454046 220678 454102
rect 220734 454046 220802 454102
rect 220858 454046 220926 454102
rect 220982 454046 251274 454102
rect 251330 454046 251398 454102
rect 251454 454046 251522 454102
rect 251578 454046 251646 454102
rect 251702 454046 272518 454102
rect 272574 454046 272642 454102
rect 272698 454046 303238 454102
rect 303294 454046 303362 454102
rect 303418 454046 343434 454102
rect 343490 454046 343558 454102
rect 343614 454046 343682 454102
rect 343738 454046 343806 454102
rect 343862 454046 374154 454102
rect 374210 454046 374278 454102
rect 374334 454046 374402 454102
rect 374458 454046 374526 454102
rect 374582 454046 404874 454102
rect 404930 454046 404998 454102
rect 405054 454046 405122 454102
rect 405178 454046 405246 454102
rect 405302 454046 435594 454102
rect 435650 454046 435718 454102
rect 435774 454046 435842 454102
rect 435898 454046 435966 454102
rect 436022 454046 466314 454102
rect 466370 454046 466438 454102
rect 466494 454046 466562 454102
rect 466618 454046 466686 454102
rect 466742 454046 497034 454102
rect 497090 454046 497158 454102
rect 497214 454046 497282 454102
rect 497338 454046 497406 454102
rect 497462 454046 527754 454102
rect 527810 454046 527878 454102
rect 527934 454046 528002 454102
rect 528058 454046 528126 454102
rect 528182 454046 558474 454102
rect 558530 454046 558598 454102
rect 558654 454046 558722 454102
rect 558778 454046 558846 454102
rect 558902 454046 589194 454102
rect 589250 454046 589318 454102
rect 589374 454046 589442 454102
rect 589498 454046 589566 454102
rect 589622 454046 596496 454102
rect 596552 454046 596620 454102
rect 596676 454046 596744 454102
rect 596800 454046 596868 454102
rect 596924 454046 597980 454102
rect -1916 453978 597980 454046
rect -1916 453922 -860 453978
rect -804 453922 -736 453978
rect -680 453922 -612 453978
rect -556 453922 -488 453978
rect -432 453922 5514 453978
rect 5570 453922 5638 453978
rect 5694 453922 5762 453978
rect 5818 453922 5886 453978
rect 5942 453922 36234 453978
rect 36290 453922 36358 453978
rect 36414 453922 36482 453978
rect 36538 453922 36606 453978
rect 36662 453922 66954 453978
rect 67010 453922 67078 453978
rect 67134 453922 67202 453978
rect 67258 453922 67326 453978
rect 67382 453922 97674 453978
rect 97730 453922 97798 453978
rect 97854 453922 97922 453978
rect 97978 453922 98046 453978
rect 98102 453922 128394 453978
rect 128450 453922 128518 453978
rect 128574 453922 128642 453978
rect 128698 453922 128766 453978
rect 128822 453922 159114 453978
rect 159170 453922 159238 453978
rect 159294 453922 159362 453978
rect 159418 453922 159486 453978
rect 159542 453922 189834 453978
rect 189890 453922 189958 453978
rect 190014 453922 190082 453978
rect 190138 453922 190206 453978
rect 190262 453922 220554 453978
rect 220610 453922 220678 453978
rect 220734 453922 220802 453978
rect 220858 453922 220926 453978
rect 220982 453922 251274 453978
rect 251330 453922 251398 453978
rect 251454 453922 251522 453978
rect 251578 453922 251646 453978
rect 251702 453922 272518 453978
rect 272574 453922 272642 453978
rect 272698 453922 303238 453978
rect 303294 453922 303362 453978
rect 303418 453922 343434 453978
rect 343490 453922 343558 453978
rect 343614 453922 343682 453978
rect 343738 453922 343806 453978
rect 343862 453922 374154 453978
rect 374210 453922 374278 453978
rect 374334 453922 374402 453978
rect 374458 453922 374526 453978
rect 374582 453922 404874 453978
rect 404930 453922 404998 453978
rect 405054 453922 405122 453978
rect 405178 453922 405246 453978
rect 405302 453922 435594 453978
rect 435650 453922 435718 453978
rect 435774 453922 435842 453978
rect 435898 453922 435966 453978
rect 436022 453922 466314 453978
rect 466370 453922 466438 453978
rect 466494 453922 466562 453978
rect 466618 453922 466686 453978
rect 466742 453922 497034 453978
rect 497090 453922 497158 453978
rect 497214 453922 497282 453978
rect 497338 453922 497406 453978
rect 497462 453922 527754 453978
rect 527810 453922 527878 453978
rect 527934 453922 528002 453978
rect 528058 453922 528126 453978
rect 528182 453922 558474 453978
rect 558530 453922 558598 453978
rect 558654 453922 558722 453978
rect 558778 453922 558846 453978
rect 558902 453922 589194 453978
rect 589250 453922 589318 453978
rect 589374 453922 589442 453978
rect 589498 453922 589566 453978
rect 589622 453922 596496 453978
rect 596552 453922 596620 453978
rect 596676 453922 596744 453978
rect 596800 453922 596868 453978
rect 596924 453922 597980 453978
rect -1916 453826 597980 453922
rect -1916 442350 597980 442446
rect -1916 442294 -1820 442350
rect -1764 442294 -1696 442350
rect -1640 442294 -1572 442350
rect -1516 442294 -1448 442350
rect -1392 442294 9234 442350
rect 9290 442294 9358 442350
rect 9414 442294 9482 442350
rect 9538 442294 9606 442350
rect 9662 442294 70674 442350
rect 70730 442294 70798 442350
rect 70854 442294 70922 442350
rect 70978 442294 71046 442350
rect 71102 442294 132114 442350
rect 132170 442294 132238 442350
rect 132294 442294 132362 442350
rect 132418 442294 132486 442350
rect 132542 442294 162834 442350
rect 162890 442294 162958 442350
rect 163014 442294 163082 442350
rect 163138 442294 163206 442350
rect 163262 442294 193554 442350
rect 193610 442294 193678 442350
rect 193734 442294 193802 442350
rect 193858 442294 193926 442350
rect 193982 442294 224274 442350
rect 224330 442294 224398 442350
rect 224454 442294 224522 442350
rect 224578 442294 224646 442350
rect 224702 442294 254994 442350
rect 255050 442294 255118 442350
rect 255174 442294 255242 442350
rect 255298 442294 255366 442350
rect 255422 442294 287878 442350
rect 287934 442294 288002 442350
rect 288058 442294 318598 442350
rect 318654 442294 318722 442350
rect 318778 442294 347154 442350
rect 347210 442294 347278 442350
rect 347334 442294 347402 442350
rect 347458 442294 347526 442350
rect 347582 442294 377874 442350
rect 377930 442294 377998 442350
rect 378054 442294 378122 442350
rect 378178 442294 378246 442350
rect 378302 442294 408594 442350
rect 408650 442294 408718 442350
rect 408774 442294 408842 442350
rect 408898 442294 408966 442350
rect 409022 442294 439314 442350
rect 439370 442294 439438 442350
rect 439494 442294 439562 442350
rect 439618 442294 439686 442350
rect 439742 442294 470034 442350
rect 470090 442294 470158 442350
rect 470214 442294 470282 442350
rect 470338 442294 470406 442350
rect 470462 442294 500754 442350
rect 500810 442294 500878 442350
rect 500934 442294 501002 442350
rect 501058 442294 501126 442350
rect 501182 442294 531474 442350
rect 531530 442294 531598 442350
rect 531654 442294 531722 442350
rect 531778 442294 531846 442350
rect 531902 442294 562194 442350
rect 562250 442294 562318 442350
rect 562374 442294 562442 442350
rect 562498 442294 562566 442350
rect 562622 442294 592914 442350
rect 592970 442294 593038 442350
rect 593094 442294 593162 442350
rect 593218 442294 593286 442350
rect 593342 442294 597456 442350
rect 597512 442294 597580 442350
rect 597636 442294 597704 442350
rect 597760 442294 597828 442350
rect 597884 442294 597980 442350
rect -1916 442226 597980 442294
rect -1916 442170 -1820 442226
rect -1764 442170 -1696 442226
rect -1640 442170 -1572 442226
rect -1516 442170 -1448 442226
rect -1392 442170 9234 442226
rect 9290 442170 9358 442226
rect 9414 442170 9482 442226
rect 9538 442170 9606 442226
rect 9662 442170 70674 442226
rect 70730 442170 70798 442226
rect 70854 442170 70922 442226
rect 70978 442170 71046 442226
rect 71102 442170 132114 442226
rect 132170 442170 132238 442226
rect 132294 442170 132362 442226
rect 132418 442170 132486 442226
rect 132542 442170 162834 442226
rect 162890 442170 162958 442226
rect 163014 442170 163082 442226
rect 163138 442170 163206 442226
rect 163262 442170 193554 442226
rect 193610 442170 193678 442226
rect 193734 442170 193802 442226
rect 193858 442170 193926 442226
rect 193982 442170 224274 442226
rect 224330 442170 224398 442226
rect 224454 442170 224522 442226
rect 224578 442170 224646 442226
rect 224702 442170 254994 442226
rect 255050 442170 255118 442226
rect 255174 442170 255242 442226
rect 255298 442170 255366 442226
rect 255422 442170 287878 442226
rect 287934 442170 288002 442226
rect 288058 442170 318598 442226
rect 318654 442170 318722 442226
rect 318778 442170 347154 442226
rect 347210 442170 347278 442226
rect 347334 442170 347402 442226
rect 347458 442170 347526 442226
rect 347582 442170 377874 442226
rect 377930 442170 377998 442226
rect 378054 442170 378122 442226
rect 378178 442170 378246 442226
rect 378302 442170 408594 442226
rect 408650 442170 408718 442226
rect 408774 442170 408842 442226
rect 408898 442170 408966 442226
rect 409022 442170 439314 442226
rect 439370 442170 439438 442226
rect 439494 442170 439562 442226
rect 439618 442170 439686 442226
rect 439742 442170 470034 442226
rect 470090 442170 470158 442226
rect 470214 442170 470282 442226
rect 470338 442170 470406 442226
rect 470462 442170 500754 442226
rect 500810 442170 500878 442226
rect 500934 442170 501002 442226
rect 501058 442170 501126 442226
rect 501182 442170 531474 442226
rect 531530 442170 531598 442226
rect 531654 442170 531722 442226
rect 531778 442170 531846 442226
rect 531902 442170 562194 442226
rect 562250 442170 562318 442226
rect 562374 442170 562442 442226
rect 562498 442170 562566 442226
rect 562622 442170 592914 442226
rect 592970 442170 593038 442226
rect 593094 442170 593162 442226
rect 593218 442170 593286 442226
rect 593342 442170 597456 442226
rect 597512 442170 597580 442226
rect 597636 442170 597704 442226
rect 597760 442170 597828 442226
rect 597884 442170 597980 442226
rect -1916 442102 597980 442170
rect -1916 442046 -1820 442102
rect -1764 442046 -1696 442102
rect -1640 442046 -1572 442102
rect -1516 442046 -1448 442102
rect -1392 442046 9234 442102
rect 9290 442046 9358 442102
rect 9414 442046 9482 442102
rect 9538 442046 9606 442102
rect 9662 442046 70674 442102
rect 70730 442046 70798 442102
rect 70854 442046 70922 442102
rect 70978 442046 71046 442102
rect 71102 442046 132114 442102
rect 132170 442046 132238 442102
rect 132294 442046 132362 442102
rect 132418 442046 132486 442102
rect 132542 442046 162834 442102
rect 162890 442046 162958 442102
rect 163014 442046 163082 442102
rect 163138 442046 163206 442102
rect 163262 442046 193554 442102
rect 193610 442046 193678 442102
rect 193734 442046 193802 442102
rect 193858 442046 193926 442102
rect 193982 442046 224274 442102
rect 224330 442046 224398 442102
rect 224454 442046 224522 442102
rect 224578 442046 224646 442102
rect 224702 442046 254994 442102
rect 255050 442046 255118 442102
rect 255174 442046 255242 442102
rect 255298 442046 255366 442102
rect 255422 442046 287878 442102
rect 287934 442046 288002 442102
rect 288058 442046 318598 442102
rect 318654 442046 318722 442102
rect 318778 442046 347154 442102
rect 347210 442046 347278 442102
rect 347334 442046 347402 442102
rect 347458 442046 347526 442102
rect 347582 442046 377874 442102
rect 377930 442046 377998 442102
rect 378054 442046 378122 442102
rect 378178 442046 378246 442102
rect 378302 442046 408594 442102
rect 408650 442046 408718 442102
rect 408774 442046 408842 442102
rect 408898 442046 408966 442102
rect 409022 442046 439314 442102
rect 439370 442046 439438 442102
rect 439494 442046 439562 442102
rect 439618 442046 439686 442102
rect 439742 442046 470034 442102
rect 470090 442046 470158 442102
rect 470214 442046 470282 442102
rect 470338 442046 470406 442102
rect 470462 442046 500754 442102
rect 500810 442046 500878 442102
rect 500934 442046 501002 442102
rect 501058 442046 501126 442102
rect 501182 442046 531474 442102
rect 531530 442046 531598 442102
rect 531654 442046 531722 442102
rect 531778 442046 531846 442102
rect 531902 442046 562194 442102
rect 562250 442046 562318 442102
rect 562374 442046 562442 442102
rect 562498 442046 562566 442102
rect 562622 442046 592914 442102
rect 592970 442046 593038 442102
rect 593094 442046 593162 442102
rect 593218 442046 593286 442102
rect 593342 442046 597456 442102
rect 597512 442046 597580 442102
rect 597636 442046 597704 442102
rect 597760 442046 597828 442102
rect 597884 442046 597980 442102
rect -1916 441978 597980 442046
rect -1916 441922 -1820 441978
rect -1764 441922 -1696 441978
rect -1640 441922 -1572 441978
rect -1516 441922 -1448 441978
rect -1392 441922 9234 441978
rect 9290 441922 9358 441978
rect 9414 441922 9482 441978
rect 9538 441922 9606 441978
rect 9662 441922 70674 441978
rect 70730 441922 70798 441978
rect 70854 441922 70922 441978
rect 70978 441922 71046 441978
rect 71102 441922 132114 441978
rect 132170 441922 132238 441978
rect 132294 441922 132362 441978
rect 132418 441922 132486 441978
rect 132542 441922 162834 441978
rect 162890 441922 162958 441978
rect 163014 441922 163082 441978
rect 163138 441922 163206 441978
rect 163262 441922 193554 441978
rect 193610 441922 193678 441978
rect 193734 441922 193802 441978
rect 193858 441922 193926 441978
rect 193982 441922 224274 441978
rect 224330 441922 224398 441978
rect 224454 441922 224522 441978
rect 224578 441922 224646 441978
rect 224702 441922 254994 441978
rect 255050 441922 255118 441978
rect 255174 441922 255242 441978
rect 255298 441922 255366 441978
rect 255422 441922 287878 441978
rect 287934 441922 288002 441978
rect 288058 441922 318598 441978
rect 318654 441922 318722 441978
rect 318778 441922 347154 441978
rect 347210 441922 347278 441978
rect 347334 441922 347402 441978
rect 347458 441922 347526 441978
rect 347582 441922 377874 441978
rect 377930 441922 377998 441978
rect 378054 441922 378122 441978
rect 378178 441922 378246 441978
rect 378302 441922 408594 441978
rect 408650 441922 408718 441978
rect 408774 441922 408842 441978
rect 408898 441922 408966 441978
rect 409022 441922 439314 441978
rect 439370 441922 439438 441978
rect 439494 441922 439562 441978
rect 439618 441922 439686 441978
rect 439742 441922 470034 441978
rect 470090 441922 470158 441978
rect 470214 441922 470282 441978
rect 470338 441922 470406 441978
rect 470462 441922 500754 441978
rect 500810 441922 500878 441978
rect 500934 441922 501002 441978
rect 501058 441922 501126 441978
rect 501182 441922 531474 441978
rect 531530 441922 531598 441978
rect 531654 441922 531722 441978
rect 531778 441922 531846 441978
rect 531902 441922 562194 441978
rect 562250 441922 562318 441978
rect 562374 441922 562442 441978
rect 562498 441922 562566 441978
rect 562622 441922 592914 441978
rect 592970 441922 593038 441978
rect 593094 441922 593162 441978
rect 593218 441922 593286 441978
rect 593342 441922 597456 441978
rect 597512 441922 597580 441978
rect 597636 441922 597704 441978
rect 597760 441922 597828 441978
rect 597884 441922 597980 441978
rect -1916 441826 597980 441922
rect -1916 436350 597980 436446
rect -1916 436294 -860 436350
rect -804 436294 -736 436350
rect -680 436294 -612 436350
rect -556 436294 -488 436350
rect -432 436294 5514 436350
rect 5570 436294 5638 436350
rect 5694 436294 5762 436350
rect 5818 436294 5886 436350
rect 5942 436294 36234 436350
rect 36290 436294 36358 436350
rect 36414 436294 36482 436350
rect 36538 436294 36606 436350
rect 36662 436294 66954 436350
rect 67010 436294 67078 436350
rect 67134 436294 67202 436350
rect 67258 436294 67326 436350
rect 67382 436294 97674 436350
rect 97730 436294 97798 436350
rect 97854 436294 97922 436350
rect 97978 436294 98046 436350
rect 98102 436294 128394 436350
rect 128450 436294 128518 436350
rect 128574 436294 128642 436350
rect 128698 436294 128766 436350
rect 128822 436294 159114 436350
rect 159170 436294 159238 436350
rect 159294 436294 159362 436350
rect 159418 436294 159486 436350
rect 159542 436294 189834 436350
rect 189890 436294 189958 436350
rect 190014 436294 190082 436350
rect 190138 436294 190206 436350
rect 190262 436294 220554 436350
rect 220610 436294 220678 436350
rect 220734 436294 220802 436350
rect 220858 436294 220926 436350
rect 220982 436294 251274 436350
rect 251330 436294 251398 436350
rect 251454 436294 251522 436350
rect 251578 436294 251646 436350
rect 251702 436294 272518 436350
rect 272574 436294 272642 436350
rect 272698 436294 303238 436350
rect 303294 436294 303362 436350
rect 303418 436294 343434 436350
rect 343490 436294 343558 436350
rect 343614 436294 343682 436350
rect 343738 436294 343806 436350
rect 343862 436294 374154 436350
rect 374210 436294 374278 436350
rect 374334 436294 374402 436350
rect 374458 436294 374526 436350
rect 374582 436294 404874 436350
rect 404930 436294 404998 436350
rect 405054 436294 405122 436350
rect 405178 436294 405246 436350
rect 405302 436294 435594 436350
rect 435650 436294 435718 436350
rect 435774 436294 435842 436350
rect 435898 436294 435966 436350
rect 436022 436294 466314 436350
rect 466370 436294 466438 436350
rect 466494 436294 466562 436350
rect 466618 436294 466686 436350
rect 466742 436294 497034 436350
rect 497090 436294 497158 436350
rect 497214 436294 497282 436350
rect 497338 436294 497406 436350
rect 497462 436294 527754 436350
rect 527810 436294 527878 436350
rect 527934 436294 528002 436350
rect 528058 436294 528126 436350
rect 528182 436294 558474 436350
rect 558530 436294 558598 436350
rect 558654 436294 558722 436350
rect 558778 436294 558846 436350
rect 558902 436294 589194 436350
rect 589250 436294 589318 436350
rect 589374 436294 589442 436350
rect 589498 436294 589566 436350
rect 589622 436294 596496 436350
rect 596552 436294 596620 436350
rect 596676 436294 596744 436350
rect 596800 436294 596868 436350
rect 596924 436294 597980 436350
rect -1916 436226 597980 436294
rect -1916 436170 -860 436226
rect -804 436170 -736 436226
rect -680 436170 -612 436226
rect -556 436170 -488 436226
rect -432 436170 5514 436226
rect 5570 436170 5638 436226
rect 5694 436170 5762 436226
rect 5818 436170 5886 436226
rect 5942 436170 36234 436226
rect 36290 436170 36358 436226
rect 36414 436170 36482 436226
rect 36538 436170 36606 436226
rect 36662 436170 66954 436226
rect 67010 436170 67078 436226
rect 67134 436170 67202 436226
rect 67258 436170 67326 436226
rect 67382 436170 97674 436226
rect 97730 436170 97798 436226
rect 97854 436170 97922 436226
rect 97978 436170 98046 436226
rect 98102 436170 128394 436226
rect 128450 436170 128518 436226
rect 128574 436170 128642 436226
rect 128698 436170 128766 436226
rect 128822 436170 159114 436226
rect 159170 436170 159238 436226
rect 159294 436170 159362 436226
rect 159418 436170 159486 436226
rect 159542 436170 189834 436226
rect 189890 436170 189958 436226
rect 190014 436170 190082 436226
rect 190138 436170 190206 436226
rect 190262 436170 220554 436226
rect 220610 436170 220678 436226
rect 220734 436170 220802 436226
rect 220858 436170 220926 436226
rect 220982 436170 251274 436226
rect 251330 436170 251398 436226
rect 251454 436170 251522 436226
rect 251578 436170 251646 436226
rect 251702 436170 272518 436226
rect 272574 436170 272642 436226
rect 272698 436170 303238 436226
rect 303294 436170 303362 436226
rect 303418 436170 343434 436226
rect 343490 436170 343558 436226
rect 343614 436170 343682 436226
rect 343738 436170 343806 436226
rect 343862 436170 374154 436226
rect 374210 436170 374278 436226
rect 374334 436170 374402 436226
rect 374458 436170 374526 436226
rect 374582 436170 404874 436226
rect 404930 436170 404998 436226
rect 405054 436170 405122 436226
rect 405178 436170 405246 436226
rect 405302 436170 435594 436226
rect 435650 436170 435718 436226
rect 435774 436170 435842 436226
rect 435898 436170 435966 436226
rect 436022 436170 466314 436226
rect 466370 436170 466438 436226
rect 466494 436170 466562 436226
rect 466618 436170 466686 436226
rect 466742 436170 497034 436226
rect 497090 436170 497158 436226
rect 497214 436170 497282 436226
rect 497338 436170 497406 436226
rect 497462 436170 527754 436226
rect 527810 436170 527878 436226
rect 527934 436170 528002 436226
rect 528058 436170 528126 436226
rect 528182 436170 558474 436226
rect 558530 436170 558598 436226
rect 558654 436170 558722 436226
rect 558778 436170 558846 436226
rect 558902 436170 589194 436226
rect 589250 436170 589318 436226
rect 589374 436170 589442 436226
rect 589498 436170 589566 436226
rect 589622 436170 596496 436226
rect 596552 436170 596620 436226
rect 596676 436170 596744 436226
rect 596800 436170 596868 436226
rect 596924 436170 597980 436226
rect -1916 436102 597980 436170
rect -1916 436046 -860 436102
rect -804 436046 -736 436102
rect -680 436046 -612 436102
rect -556 436046 -488 436102
rect -432 436046 5514 436102
rect 5570 436046 5638 436102
rect 5694 436046 5762 436102
rect 5818 436046 5886 436102
rect 5942 436046 36234 436102
rect 36290 436046 36358 436102
rect 36414 436046 36482 436102
rect 36538 436046 36606 436102
rect 36662 436046 66954 436102
rect 67010 436046 67078 436102
rect 67134 436046 67202 436102
rect 67258 436046 67326 436102
rect 67382 436046 97674 436102
rect 97730 436046 97798 436102
rect 97854 436046 97922 436102
rect 97978 436046 98046 436102
rect 98102 436046 128394 436102
rect 128450 436046 128518 436102
rect 128574 436046 128642 436102
rect 128698 436046 128766 436102
rect 128822 436046 159114 436102
rect 159170 436046 159238 436102
rect 159294 436046 159362 436102
rect 159418 436046 159486 436102
rect 159542 436046 189834 436102
rect 189890 436046 189958 436102
rect 190014 436046 190082 436102
rect 190138 436046 190206 436102
rect 190262 436046 220554 436102
rect 220610 436046 220678 436102
rect 220734 436046 220802 436102
rect 220858 436046 220926 436102
rect 220982 436046 251274 436102
rect 251330 436046 251398 436102
rect 251454 436046 251522 436102
rect 251578 436046 251646 436102
rect 251702 436046 272518 436102
rect 272574 436046 272642 436102
rect 272698 436046 303238 436102
rect 303294 436046 303362 436102
rect 303418 436046 343434 436102
rect 343490 436046 343558 436102
rect 343614 436046 343682 436102
rect 343738 436046 343806 436102
rect 343862 436046 374154 436102
rect 374210 436046 374278 436102
rect 374334 436046 374402 436102
rect 374458 436046 374526 436102
rect 374582 436046 404874 436102
rect 404930 436046 404998 436102
rect 405054 436046 405122 436102
rect 405178 436046 405246 436102
rect 405302 436046 435594 436102
rect 435650 436046 435718 436102
rect 435774 436046 435842 436102
rect 435898 436046 435966 436102
rect 436022 436046 466314 436102
rect 466370 436046 466438 436102
rect 466494 436046 466562 436102
rect 466618 436046 466686 436102
rect 466742 436046 497034 436102
rect 497090 436046 497158 436102
rect 497214 436046 497282 436102
rect 497338 436046 497406 436102
rect 497462 436046 527754 436102
rect 527810 436046 527878 436102
rect 527934 436046 528002 436102
rect 528058 436046 528126 436102
rect 528182 436046 558474 436102
rect 558530 436046 558598 436102
rect 558654 436046 558722 436102
rect 558778 436046 558846 436102
rect 558902 436046 589194 436102
rect 589250 436046 589318 436102
rect 589374 436046 589442 436102
rect 589498 436046 589566 436102
rect 589622 436046 596496 436102
rect 596552 436046 596620 436102
rect 596676 436046 596744 436102
rect 596800 436046 596868 436102
rect 596924 436046 597980 436102
rect -1916 435978 597980 436046
rect -1916 435922 -860 435978
rect -804 435922 -736 435978
rect -680 435922 -612 435978
rect -556 435922 -488 435978
rect -432 435922 5514 435978
rect 5570 435922 5638 435978
rect 5694 435922 5762 435978
rect 5818 435922 5886 435978
rect 5942 435922 36234 435978
rect 36290 435922 36358 435978
rect 36414 435922 36482 435978
rect 36538 435922 36606 435978
rect 36662 435922 66954 435978
rect 67010 435922 67078 435978
rect 67134 435922 67202 435978
rect 67258 435922 67326 435978
rect 67382 435922 97674 435978
rect 97730 435922 97798 435978
rect 97854 435922 97922 435978
rect 97978 435922 98046 435978
rect 98102 435922 128394 435978
rect 128450 435922 128518 435978
rect 128574 435922 128642 435978
rect 128698 435922 128766 435978
rect 128822 435922 159114 435978
rect 159170 435922 159238 435978
rect 159294 435922 159362 435978
rect 159418 435922 159486 435978
rect 159542 435922 189834 435978
rect 189890 435922 189958 435978
rect 190014 435922 190082 435978
rect 190138 435922 190206 435978
rect 190262 435922 220554 435978
rect 220610 435922 220678 435978
rect 220734 435922 220802 435978
rect 220858 435922 220926 435978
rect 220982 435922 251274 435978
rect 251330 435922 251398 435978
rect 251454 435922 251522 435978
rect 251578 435922 251646 435978
rect 251702 435922 272518 435978
rect 272574 435922 272642 435978
rect 272698 435922 303238 435978
rect 303294 435922 303362 435978
rect 303418 435922 343434 435978
rect 343490 435922 343558 435978
rect 343614 435922 343682 435978
rect 343738 435922 343806 435978
rect 343862 435922 374154 435978
rect 374210 435922 374278 435978
rect 374334 435922 374402 435978
rect 374458 435922 374526 435978
rect 374582 435922 404874 435978
rect 404930 435922 404998 435978
rect 405054 435922 405122 435978
rect 405178 435922 405246 435978
rect 405302 435922 435594 435978
rect 435650 435922 435718 435978
rect 435774 435922 435842 435978
rect 435898 435922 435966 435978
rect 436022 435922 466314 435978
rect 466370 435922 466438 435978
rect 466494 435922 466562 435978
rect 466618 435922 466686 435978
rect 466742 435922 497034 435978
rect 497090 435922 497158 435978
rect 497214 435922 497282 435978
rect 497338 435922 497406 435978
rect 497462 435922 527754 435978
rect 527810 435922 527878 435978
rect 527934 435922 528002 435978
rect 528058 435922 528126 435978
rect 528182 435922 558474 435978
rect 558530 435922 558598 435978
rect 558654 435922 558722 435978
rect 558778 435922 558846 435978
rect 558902 435922 589194 435978
rect 589250 435922 589318 435978
rect 589374 435922 589442 435978
rect 589498 435922 589566 435978
rect 589622 435922 596496 435978
rect 596552 435922 596620 435978
rect 596676 435922 596744 435978
rect 596800 435922 596868 435978
rect 596924 435922 597980 435978
rect -1916 435826 597980 435922
rect -1916 424350 597980 424446
rect -1916 424294 -1820 424350
rect -1764 424294 -1696 424350
rect -1640 424294 -1572 424350
rect -1516 424294 -1448 424350
rect -1392 424294 9234 424350
rect 9290 424294 9358 424350
rect 9414 424294 9482 424350
rect 9538 424294 9606 424350
rect 9662 424294 70674 424350
rect 70730 424294 70798 424350
rect 70854 424294 70922 424350
rect 70978 424294 71046 424350
rect 71102 424294 132114 424350
rect 132170 424294 132238 424350
rect 132294 424294 132362 424350
rect 132418 424294 132486 424350
rect 132542 424294 162834 424350
rect 162890 424294 162958 424350
rect 163014 424294 163082 424350
rect 163138 424294 163206 424350
rect 163262 424294 193554 424350
rect 193610 424294 193678 424350
rect 193734 424294 193802 424350
rect 193858 424294 193926 424350
rect 193982 424294 224274 424350
rect 224330 424294 224398 424350
rect 224454 424294 224522 424350
rect 224578 424294 224646 424350
rect 224702 424294 254994 424350
rect 255050 424294 255118 424350
rect 255174 424294 255242 424350
rect 255298 424294 255366 424350
rect 255422 424294 287878 424350
rect 287934 424294 288002 424350
rect 288058 424294 318598 424350
rect 318654 424294 318722 424350
rect 318778 424294 347154 424350
rect 347210 424294 347278 424350
rect 347334 424294 347402 424350
rect 347458 424294 347526 424350
rect 347582 424294 377874 424350
rect 377930 424294 377998 424350
rect 378054 424294 378122 424350
rect 378178 424294 378246 424350
rect 378302 424294 408594 424350
rect 408650 424294 408718 424350
rect 408774 424294 408842 424350
rect 408898 424294 408966 424350
rect 409022 424294 439314 424350
rect 439370 424294 439438 424350
rect 439494 424294 439562 424350
rect 439618 424294 439686 424350
rect 439742 424294 470034 424350
rect 470090 424294 470158 424350
rect 470214 424294 470282 424350
rect 470338 424294 470406 424350
rect 470462 424294 500754 424350
rect 500810 424294 500878 424350
rect 500934 424294 501002 424350
rect 501058 424294 501126 424350
rect 501182 424294 531474 424350
rect 531530 424294 531598 424350
rect 531654 424294 531722 424350
rect 531778 424294 531846 424350
rect 531902 424294 562194 424350
rect 562250 424294 562318 424350
rect 562374 424294 562442 424350
rect 562498 424294 562566 424350
rect 562622 424294 592914 424350
rect 592970 424294 593038 424350
rect 593094 424294 593162 424350
rect 593218 424294 593286 424350
rect 593342 424294 597456 424350
rect 597512 424294 597580 424350
rect 597636 424294 597704 424350
rect 597760 424294 597828 424350
rect 597884 424294 597980 424350
rect -1916 424226 597980 424294
rect -1916 424170 -1820 424226
rect -1764 424170 -1696 424226
rect -1640 424170 -1572 424226
rect -1516 424170 -1448 424226
rect -1392 424170 9234 424226
rect 9290 424170 9358 424226
rect 9414 424170 9482 424226
rect 9538 424170 9606 424226
rect 9662 424170 70674 424226
rect 70730 424170 70798 424226
rect 70854 424170 70922 424226
rect 70978 424170 71046 424226
rect 71102 424170 132114 424226
rect 132170 424170 132238 424226
rect 132294 424170 132362 424226
rect 132418 424170 132486 424226
rect 132542 424170 162834 424226
rect 162890 424170 162958 424226
rect 163014 424170 163082 424226
rect 163138 424170 163206 424226
rect 163262 424170 193554 424226
rect 193610 424170 193678 424226
rect 193734 424170 193802 424226
rect 193858 424170 193926 424226
rect 193982 424170 224274 424226
rect 224330 424170 224398 424226
rect 224454 424170 224522 424226
rect 224578 424170 224646 424226
rect 224702 424170 254994 424226
rect 255050 424170 255118 424226
rect 255174 424170 255242 424226
rect 255298 424170 255366 424226
rect 255422 424170 287878 424226
rect 287934 424170 288002 424226
rect 288058 424170 318598 424226
rect 318654 424170 318722 424226
rect 318778 424170 347154 424226
rect 347210 424170 347278 424226
rect 347334 424170 347402 424226
rect 347458 424170 347526 424226
rect 347582 424170 377874 424226
rect 377930 424170 377998 424226
rect 378054 424170 378122 424226
rect 378178 424170 378246 424226
rect 378302 424170 408594 424226
rect 408650 424170 408718 424226
rect 408774 424170 408842 424226
rect 408898 424170 408966 424226
rect 409022 424170 439314 424226
rect 439370 424170 439438 424226
rect 439494 424170 439562 424226
rect 439618 424170 439686 424226
rect 439742 424170 470034 424226
rect 470090 424170 470158 424226
rect 470214 424170 470282 424226
rect 470338 424170 470406 424226
rect 470462 424170 500754 424226
rect 500810 424170 500878 424226
rect 500934 424170 501002 424226
rect 501058 424170 501126 424226
rect 501182 424170 531474 424226
rect 531530 424170 531598 424226
rect 531654 424170 531722 424226
rect 531778 424170 531846 424226
rect 531902 424170 562194 424226
rect 562250 424170 562318 424226
rect 562374 424170 562442 424226
rect 562498 424170 562566 424226
rect 562622 424170 592914 424226
rect 592970 424170 593038 424226
rect 593094 424170 593162 424226
rect 593218 424170 593286 424226
rect 593342 424170 597456 424226
rect 597512 424170 597580 424226
rect 597636 424170 597704 424226
rect 597760 424170 597828 424226
rect 597884 424170 597980 424226
rect -1916 424102 597980 424170
rect -1916 424046 -1820 424102
rect -1764 424046 -1696 424102
rect -1640 424046 -1572 424102
rect -1516 424046 -1448 424102
rect -1392 424046 9234 424102
rect 9290 424046 9358 424102
rect 9414 424046 9482 424102
rect 9538 424046 9606 424102
rect 9662 424046 70674 424102
rect 70730 424046 70798 424102
rect 70854 424046 70922 424102
rect 70978 424046 71046 424102
rect 71102 424046 132114 424102
rect 132170 424046 132238 424102
rect 132294 424046 132362 424102
rect 132418 424046 132486 424102
rect 132542 424046 162834 424102
rect 162890 424046 162958 424102
rect 163014 424046 163082 424102
rect 163138 424046 163206 424102
rect 163262 424046 193554 424102
rect 193610 424046 193678 424102
rect 193734 424046 193802 424102
rect 193858 424046 193926 424102
rect 193982 424046 224274 424102
rect 224330 424046 224398 424102
rect 224454 424046 224522 424102
rect 224578 424046 224646 424102
rect 224702 424046 254994 424102
rect 255050 424046 255118 424102
rect 255174 424046 255242 424102
rect 255298 424046 255366 424102
rect 255422 424046 287878 424102
rect 287934 424046 288002 424102
rect 288058 424046 318598 424102
rect 318654 424046 318722 424102
rect 318778 424046 347154 424102
rect 347210 424046 347278 424102
rect 347334 424046 347402 424102
rect 347458 424046 347526 424102
rect 347582 424046 377874 424102
rect 377930 424046 377998 424102
rect 378054 424046 378122 424102
rect 378178 424046 378246 424102
rect 378302 424046 408594 424102
rect 408650 424046 408718 424102
rect 408774 424046 408842 424102
rect 408898 424046 408966 424102
rect 409022 424046 439314 424102
rect 439370 424046 439438 424102
rect 439494 424046 439562 424102
rect 439618 424046 439686 424102
rect 439742 424046 470034 424102
rect 470090 424046 470158 424102
rect 470214 424046 470282 424102
rect 470338 424046 470406 424102
rect 470462 424046 500754 424102
rect 500810 424046 500878 424102
rect 500934 424046 501002 424102
rect 501058 424046 501126 424102
rect 501182 424046 531474 424102
rect 531530 424046 531598 424102
rect 531654 424046 531722 424102
rect 531778 424046 531846 424102
rect 531902 424046 562194 424102
rect 562250 424046 562318 424102
rect 562374 424046 562442 424102
rect 562498 424046 562566 424102
rect 562622 424046 592914 424102
rect 592970 424046 593038 424102
rect 593094 424046 593162 424102
rect 593218 424046 593286 424102
rect 593342 424046 597456 424102
rect 597512 424046 597580 424102
rect 597636 424046 597704 424102
rect 597760 424046 597828 424102
rect 597884 424046 597980 424102
rect -1916 423978 597980 424046
rect -1916 423922 -1820 423978
rect -1764 423922 -1696 423978
rect -1640 423922 -1572 423978
rect -1516 423922 -1448 423978
rect -1392 423922 9234 423978
rect 9290 423922 9358 423978
rect 9414 423922 9482 423978
rect 9538 423922 9606 423978
rect 9662 423922 70674 423978
rect 70730 423922 70798 423978
rect 70854 423922 70922 423978
rect 70978 423922 71046 423978
rect 71102 423922 132114 423978
rect 132170 423922 132238 423978
rect 132294 423922 132362 423978
rect 132418 423922 132486 423978
rect 132542 423922 162834 423978
rect 162890 423922 162958 423978
rect 163014 423922 163082 423978
rect 163138 423922 163206 423978
rect 163262 423922 193554 423978
rect 193610 423922 193678 423978
rect 193734 423922 193802 423978
rect 193858 423922 193926 423978
rect 193982 423922 224274 423978
rect 224330 423922 224398 423978
rect 224454 423922 224522 423978
rect 224578 423922 224646 423978
rect 224702 423922 254994 423978
rect 255050 423922 255118 423978
rect 255174 423922 255242 423978
rect 255298 423922 255366 423978
rect 255422 423922 287878 423978
rect 287934 423922 288002 423978
rect 288058 423922 318598 423978
rect 318654 423922 318722 423978
rect 318778 423922 347154 423978
rect 347210 423922 347278 423978
rect 347334 423922 347402 423978
rect 347458 423922 347526 423978
rect 347582 423922 377874 423978
rect 377930 423922 377998 423978
rect 378054 423922 378122 423978
rect 378178 423922 378246 423978
rect 378302 423922 408594 423978
rect 408650 423922 408718 423978
rect 408774 423922 408842 423978
rect 408898 423922 408966 423978
rect 409022 423922 439314 423978
rect 439370 423922 439438 423978
rect 439494 423922 439562 423978
rect 439618 423922 439686 423978
rect 439742 423922 470034 423978
rect 470090 423922 470158 423978
rect 470214 423922 470282 423978
rect 470338 423922 470406 423978
rect 470462 423922 500754 423978
rect 500810 423922 500878 423978
rect 500934 423922 501002 423978
rect 501058 423922 501126 423978
rect 501182 423922 531474 423978
rect 531530 423922 531598 423978
rect 531654 423922 531722 423978
rect 531778 423922 531846 423978
rect 531902 423922 562194 423978
rect 562250 423922 562318 423978
rect 562374 423922 562442 423978
rect 562498 423922 562566 423978
rect 562622 423922 592914 423978
rect 592970 423922 593038 423978
rect 593094 423922 593162 423978
rect 593218 423922 593286 423978
rect 593342 423922 597456 423978
rect 597512 423922 597580 423978
rect 597636 423922 597704 423978
rect 597760 423922 597828 423978
rect 597884 423922 597980 423978
rect -1916 423826 597980 423922
rect 350236 420058 472180 420074
rect 350236 420002 350252 420058
rect 350308 420002 472108 420058
rect 472164 420002 472180 420058
rect 350236 419986 472180 420002
rect -1916 418350 597980 418446
rect -1916 418294 -860 418350
rect -804 418294 -736 418350
rect -680 418294 -612 418350
rect -556 418294 -488 418350
rect -432 418294 5514 418350
rect 5570 418294 5638 418350
rect 5694 418294 5762 418350
rect 5818 418294 5886 418350
rect 5942 418294 24518 418350
rect 24574 418294 24642 418350
rect 24698 418294 36234 418350
rect 36290 418294 36358 418350
rect 36414 418294 36482 418350
rect 36538 418294 36606 418350
rect 36662 418294 55238 418350
rect 55294 418294 55362 418350
rect 55418 418294 66954 418350
rect 67010 418294 67078 418350
rect 67134 418294 67202 418350
rect 67258 418294 67326 418350
rect 67382 418294 86518 418350
rect 86574 418294 86642 418350
rect 86698 418294 97674 418350
rect 97730 418294 97798 418350
rect 97854 418294 97922 418350
rect 97978 418294 98046 418350
rect 98102 418294 117238 418350
rect 117294 418294 117362 418350
rect 117418 418294 128394 418350
rect 128450 418294 128518 418350
rect 128574 418294 128642 418350
rect 128698 418294 128766 418350
rect 128822 418294 148518 418350
rect 148574 418294 148642 418350
rect 148698 418294 159114 418350
rect 159170 418294 159238 418350
rect 159294 418294 159362 418350
rect 159418 418294 159486 418350
rect 159542 418294 179238 418350
rect 179294 418294 179362 418350
rect 179418 418294 189834 418350
rect 189890 418294 189958 418350
rect 190014 418294 190082 418350
rect 190138 418294 190206 418350
rect 190262 418294 210518 418350
rect 210574 418294 210642 418350
rect 210698 418294 220554 418350
rect 220610 418294 220678 418350
rect 220734 418294 220802 418350
rect 220858 418294 220926 418350
rect 220982 418294 241238 418350
rect 241294 418294 241362 418350
rect 241418 418294 251274 418350
rect 251330 418294 251398 418350
rect 251454 418294 251522 418350
rect 251578 418294 251646 418350
rect 251702 418294 272518 418350
rect 272574 418294 272642 418350
rect 272698 418294 303238 418350
rect 303294 418294 303362 418350
rect 303418 418294 343434 418350
rect 343490 418294 343558 418350
rect 343614 418294 343682 418350
rect 343738 418294 343806 418350
rect 343862 418294 356518 418350
rect 356574 418294 356642 418350
rect 356698 418294 374154 418350
rect 374210 418294 374278 418350
rect 374334 418294 374402 418350
rect 374458 418294 374526 418350
rect 374582 418294 387238 418350
rect 387294 418294 387362 418350
rect 387418 418294 404874 418350
rect 404930 418294 404998 418350
rect 405054 418294 405122 418350
rect 405178 418294 405246 418350
rect 405302 418294 418518 418350
rect 418574 418294 418642 418350
rect 418698 418294 435594 418350
rect 435650 418294 435718 418350
rect 435774 418294 435842 418350
rect 435898 418294 435966 418350
rect 436022 418294 449238 418350
rect 449294 418294 449362 418350
rect 449418 418294 466314 418350
rect 466370 418294 466438 418350
rect 466494 418294 466562 418350
rect 466618 418294 466686 418350
rect 466742 418294 480518 418350
rect 480574 418294 480642 418350
rect 480698 418294 497034 418350
rect 497090 418294 497158 418350
rect 497214 418294 497282 418350
rect 497338 418294 497406 418350
rect 497462 418294 511238 418350
rect 511294 418294 511362 418350
rect 511418 418294 527754 418350
rect 527810 418294 527878 418350
rect 527934 418294 528002 418350
rect 528058 418294 528126 418350
rect 528182 418294 542518 418350
rect 542574 418294 542642 418350
rect 542698 418294 558474 418350
rect 558530 418294 558598 418350
rect 558654 418294 558722 418350
rect 558778 418294 558846 418350
rect 558902 418294 573238 418350
rect 573294 418294 573362 418350
rect 573418 418294 589194 418350
rect 589250 418294 589318 418350
rect 589374 418294 589442 418350
rect 589498 418294 589566 418350
rect 589622 418294 596496 418350
rect 596552 418294 596620 418350
rect 596676 418294 596744 418350
rect 596800 418294 596868 418350
rect 596924 418294 597980 418350
rect -1916 418226 597980 418294
rect -1916 418170 -860 418226
rect -804 418170 -736 418226
rect -680 418170 -612 418226
rect -556 418170 -488 418226
rect -432 418170 5514 418226
rect 5570 418170 5638 418226
rect 5694 418170 5762 418226
rect 5818 418170 5886 418226
rect 5942 418170 24518 418226
rect 24574 418170 24642 418226
rect 24698 418170 36234 418226
rect 36290 418170 36358 418226
rect 36414 418170 36482 418226
rect 36538 418170 36606 418226
rect 36662 418170 55238 418226
rect 55294 418170 55362 418226
rect 55418 418170 66954 418226
rect 67010 418170 67078 418226
rect 67134 418170 67202 418226
rect 67258 418170 67326 418226
rect 67382 418170 86518 418226
rect 86574 418170 86642 418226
rect 86698 418170 97674 418226
rect 97730 418170 97798 418226
rect 97854 418170 97922 418226
rect 97978 418170 98046 418226
rect 98102 418170 117238 418226
rect 117294 418170 117362 418226
rect 117418 418170 128394 418226
rect 128450 418170 128518 418226
rect 128574 418170 128642 418226
rect 128698 418170 128766 418226
rect 128822 418170 148518 418226
rect 148574 418170 148642 418226
rect 148698 418170 159114 418226
rect 159170 418170 159238 418226
rect 159294 418170 159362 418226
rect 159418 418170 159486 418226
rect 159542 418170 179238 418226
rect 179294 418170 179362 418226
rect 179418 418170 189834 418226
rect 189890 418170 189958 418226
rect 190014 418170 190082 418226
rect 190138 418170 190206 418226
rect 190262 418170 210518 418226
rect 210574 418170 210642 418226
rect 210698 418170 220554 418226
rect 220610 418170 220678 418226
rect 220734 418170 220802 418226
rect 220858 418170 220926 418226
rect 220982 418170 241238 418226
rect 241294 418170 241362 418226
rect 241418 418170 251274 418226
rect 251330 418170 251398 418226
rect 251454 418170 251522 418226
rect 251578 418170 251646 418226
rect 251702 418170 272518 418226
rect 272574 418170 272642 418226
rect 272698 418170 303238 418226
rect 303294 418170 303362 418226
rect 303418 418170 343434 418226
rect 343490 418170 343558 418226
rect 343614 418170 343682 418226
rect 343738 418170 343806 418226
rect 343862 418170 356518 418226
rect 356574 418170 356642 418226
rect 356698 418170 374154 418226
rect 374210 418170 374278 418226
rect 374334 418170 374402 418226
rect 374458 418170 374526 418226
rect 374582 418170 387238 418226
rect 387294 418170 387362 418226
rect 387418 418170 404874 418226
rect 404930 418170 404998 418226
rect 405054 418170 405122 418226
rect 405178 418170 405246 418226
rect 405302 418170 418518 418226
rect 418574 418170 418642 418226
rect 418698 418170 435594 418226
rect 435650 418170 435718 418226
rect 435774 418170 435842 418226
rect 435898 418170 435966 418226
rect 436022 418170 449238 418226
rect 449294 418170 449362 418226
rect 449418 418170 466314 418226
rect 466370 418170 466438 418226
rect 466494 418170 466562 418226
rect 466618 418170 466686 418226
rect 466742 418170 480518 418226
rect 480574 418170 480642 418226
rect 480698 418170 497034 418226
rect 497090 418170 497158 418226
rect 497214 418170 497282 418226
rect 497338 418170 497406 418226
rect 497462 418170 511238 418226
rect 511294 418170 511362 418226
rect 511418 418170 527754 418226
rect 527810 418170 527878 418226
rect 527934 418170 528002 418226
rect 528058 418170 528126 418226
rect 528182 418170 542518 418226
rect 542574 418170 542642 418226
rect 542698 418170 558474 418226
rect 558530 418170 558598 418226
rect 558654 418170 558722 418226
rect 558778 418170 558846 418226
rect 558902 418170 573238 418226
rect 573294 418170 573362 418226
rect 573418 418170 589194 418226
rect 589250 418170 589318 418226
rect 589374 418170 589442 418226
rect 589498 418170 589566 418226
rect 589622 418170 596496 418226
rect 596552 418170 596620 418226
rect 596676 418170 596744 418226
rect 596800 418170 596868 418226
rect 596924 418170 597980 418226
rect -1916 418102 597980 418170
rect -1916 418046 -860 418102
rect -804 418046 -736 418102
rect -680 418046 -612 418102
rect -556 418046 -488 418102
rect -432 418046 5514 418102
rect 5570 418046 5638 418102
rect 5694 418046 5762 418102
rect 5818 418046 5886 418102
rect 5942 418046 24518 418102
rect 24574 418046 24642 418102
rect 24698 418046 36234 418102
rect 36290 418046 36358 418102
rect 36414 418046 36482 418102
rect 36538 418046 36606 418102
rect 36662 418046 55238 418102
rect 55294 418046 55362 418102
rect 55418 418046 66954 418102
rect 67010 418046 67078 418102
rect 67134 418046 67202 418102
rect 67258 418046 67326 418102
rect 67382 418046 86518 418102
rect 86574 418046 86642 418102
rect 86698 418046 97674 418102
rect 97730 418046 97798 418102
rect 97854 418046 97922 418102
rect 97978 418046 98046 418102
rect 98102 418046 117238 418102
rect 117294 418046 117362 418102
rect 117418 418046 128394 418102
rect 128450 418046 128518 418102
rect 128574 418046 128642 418102
rect 128698 418046 128766 418102
rect 128822 418046 148518 418102
rect 148574 418046 148642 418102
rect 148698 418046 159114 418102
rect 159170 418046 159238 418102
rect 159294 418046 159362 418102
rect 159418 418046 159486 418102
rect 159542 418046 179238 418102
rect 179294 418046 179362 418102
rect 179418 418046 189834 418102
rect 189890 418046 189958 418102
rect 190014 418046 190082 418102
rect 190138 418046 190206 418102
rect 190262 418046 210518 418102
rect 210574 418046 210642 418102
rect 210698 418046 220554 418102
rect 220610 418046 220678 418102
rect 220734 418046 220802 418102
rect 220858 418046 220926 418102
rect 220982 418046 241238 418102
rect 241294 418046 241362 418102
rect 241418 418046 251274 418102
rect 251330 418046 251398 418102
rect 251454 418046 251522 418102
rect 251578 418046 251646 418102
rect 251702 418046 272518 418102
rect 272574 418046 272642 418102
rect 272698 418046 303238 418102
rect 303294 418046 303362 418102
rect 303418 418046 343434 418102
rect 343490 418046 343558 418102
rect 343614 418046 343682 418102
rect 343738 418046 343806 418102
rect 343862 418046 356518 418102
rect 356574 418046 356642 418102
rect 356698 418046 374154 418102
rect 374210 418046 374278 418102
rect 374334 418046 374402 418102
rect 374458 418046 374526 418102
rect 374582 418046 387238 418102
rect 387294 418046 387362 418102
rect 387418 418046 404874 418102
rect 404930 418046 404998 418102
rect 405054 418046 405122 418102
rect 405178 418046 405246 418102
rect 405302 418046 418518 418102
rect 418574 418046 418642 418102
rect 418698 418046 435594 418102
rect 435650 418046 435718 418102
rect 435774 418046 435842 418102
rect 435898 418046 435966 418102
rect 436022 418046 449238 418102
rect 449294 418046 449362 418102
rect 449418 418046 466314 418102
rect 466370 418046 466438 418102
rect 466494 418046 466562 418102
rect 466618 418046 466686 418102
rect 466742 418046 480518 418102
rect 480574 418046 480642 418102
rect 480698 418046 497034 418102
rect 497090 418046 497158 418102
rect 497214 418046 497282 418102
rect 497338 418046 497406 418102
rect 497462 418046 511238 418102
rect 511294 418046 511362 418102
rect 511418 418046 527754 418102
rect 527810 418046 527878 418102
rect 527934 418046 528002 418102
rect 528058 418046 528126 418102
rect 528182 418046 542518 418102
rect 542574 418046 542642 418102
rect 542698 418046 558474 418102
rect 558530 418046 558598 418102
rect 558654 418046 558722 418102
rect 558778 418046 558846 418102
rect 558902 418046 573238 418102
rect 573294 418046 573362 418102
rect 573418 418046 589194 418102
rect 589250 418046 589318 418102
rect 589374 418046 589442 418102
rect 589498 418046 589566 418102
rect 589622 418046 596496 418102
rect 596552 418046 596620 418102
rect 596676 418046 596744 418102
rect 596800 418046 596868 418102
rect 596924 418046 597980 418102
rect -1916 417978 597980 418046
rect -1916 417922 -860 417978
rect -804 417922 -736 417978
rect -680 417922 -612 417978
rect -556 417922 -488 417978
rect -432 417922 5514 417978
rect 5570 417922 5638 417978
rect 5694 417922 5762 417978
rect 5818 417922 5886 417978
rect 5942 417922 24518 417978
rect 24574 417922 24642 417978
rect 24698 417922 36234 417978
rect 36290 417922 36358 417978
rect 36414 417922 36482 417978
rect 36538 417922 36606 417978
rect 36662 417922 55238 417978
rect 55294 417922 55362 417978
rect 55418 417922 66954 417978
rect 67010 417922 67078 417978
rect 67134 417922 67202 417978
rect 67258 417922 67326 417978
rect 67382 417922 86518 417978
rect 86574 417922 86642 417978
rect 86698 417922 97674 417978
rect 97730 417922 97798 417978
rect 97854 417922 97922 417978
rect 97978 417922 98046 417978
rect 98102 417922 117238 417978
rect 117294 417922 117362 417978
rect 117418 417922 128394 417978
rect 128450 417922 128518 417978
rect 128574 417922 128642 417978
rect 128698 417922 128766 417978
rect 128822 417922 148518 417978
rect 148574 417922 148642 417978
rect 148698 417922 159114 417978
rect 159170 417922 159238 417978
rect 159294 417922 159362 417978
rect 159418 417922 159486 417978
rect 159542 417922 179238 417978
rect 179294 417922 179362 417978
rect 179418 417922 189834 417978
rect 189890 417922 189958 417978
rect 190014 417922 190082 417978
rect 190138 417922 190206 417978
rect 190262 417922 210518 417978
rect 210574 417922 210642 417978
rect 210698 417922 220554 417978
rect 220610 417922 220678 417978
rect 220734 417922 220802 417978
rect 220858 417922 220926 417978
rect 220982 417922 241238 417978
rect 241294 417922 241362 417978
rect 241418 417922 251274 417978
rect 251330 417922 251398 417978
rect 251454 417922 251522 417978
rect 251578 417922 251646 417978
rect 251702 417922 272518 417978
rect 272574 417922 272642 417978
rect 272698 417922 303238 417978
rect 303294 417922 303362 417978
rect 303418 417922 343434 417978
rect 343490 417922 343558 417978
rect 343614 417922 343682 417978
rect 343738 417922 343806 417978
rect 343862 417922 356518 417978
rect 356574 417922 356642 417978
rect 356698 417922 374154 417978
rect 374210 417922 374278 417978
rect 374334 417922 374402 417978
rect 374458 417922 374526 417978
rect 374582 417922 387238 417978
rect 387294 417922 387362 417978
rect 387418 417922 404874 417978
rect 404930 417922 404998 417978
rect 405054 417922 405122 417978
rect 405178 417922 405246 417978
rect 405302 417922 418518 417978
rect 418574 417922 418642 417978
rect 418698 417922 435594 417978
rect 435650 417922 435718 417978
rect 435774 417922 435842 417978
rect 435898 417922 435966 417978
rect 436022 417922 449238 417978
rect 449294 417922 449362 417978
rect 449418 417922 466314 417978
rect 466370 417922 466438 417978
rect 466494 417922 466562 417978
rect 466618 417922 466686 417978
rect 466742 417922 480518 417978
rect 480574 417922 480642 417978
rect 480698 417922 497034 417978
rect 497090 417922 497158 417978
rect 497214 417922 497282 417978
rect 497338 417922 497406 417978
rect 497462 417922 511238 417978
rect 511294 417922 511362 417978
rect 511418 417922 527754 417978
rect 527810 417922 527878 417978
rect 527934 417922 528002 417978
rect 528058 417922 528126 417978
rect 528182 417922 542518 417978
rect 542574 417922 542642 417978
rect 542698 417922 558474 417978
rect 558530 417922 558598 417978
rect 558654 417922 558722 417978
rect 558778 417922 558846 417978
rect 558902 417922 573238 417978
rect 573294 417922 573362 417978
rect 573418 417922 589194 417978
rect 589250 417922 589318 417978
rect 589374 417922 589442 417978
rect 589498 417922 589566 417978
rect 589622 417922 596496 417978
rect 596552 417922 596620 417978
rect 596676 417922 596744 417978
rect 596800 417922 596868 417978
rect 596924 417922 597980 417978
rect -1916 417826 597980 417922
rect 206652 415018 260388 415034
rect 206652 414962 206668 415018
rect 206724 414962 260316 415018
rect 260372 414962 260388 415018
rect 206652 414946 260388 414962
rect 334444 415018 523364 415034
rect 334444 414962 334460 415018
rect 334516 414962 523292 415018
rect 523348 414962 523364 415018
rect 334444 414946 523364 414962
rect 334444 413758 414164 413774
rect 334444 413702 334460 413758
rect 334516 413702 414092 413758
rect 414148 413702 414164 413758
rect 334444 413686 414164 413702
rect 334444 413578 518324 413594
rect 334444 413522 334460 413578
rect 334516 413522 518252 413578
rect 518308 413522 518324 413578
rect 334444 413506 518324 413522
rect 414636 413398 472180 413414
rect 414636 413342 414652 413398
rect 414708 413342 472108 413398
rect 472164 413342 472180 413398
rect 414636 413326 472180 413342
rect 18380 413218 79004 413234
rect 18380 413162 18396 413218
rect 18452 413162 79004 413218
rect 18380 413146 79004 413162
rect 78916 412514 79004 413146
rect 144044 412678 149564 412694
rect 144044 412622 144060 412678
rect 144116 412622 149564 412678
rect 144044 412606 149564 412622
rect 149476 412514 149564 412606
rect 78916 412498 141108 412514
rect 78916 412442 82684 412498
rect 82740 412442 141036 412498
rect 141092 412442 141108 412498
rect 78916 412426 141108 412442
rect 149476 412498 201700 412514
rect 149476 412442 201628 412498
rect 201684 412442 201700 412498
rect 149476 412426 201700 412442
rect 428860 412138 472180 412154
rect 428860 412082 428876 412138
rect 428932 412082 472108 412138
rect 472164 412082 472180 412138
rect 428860 412066 472180 412082
rect 334444 411958 441044 411974
rect 334444 411902 334460 411958
rect 334516 411902 440972 411958
rect 441028 411902 441044 411958
rect 334444 411886 441044 411902
rect 204748 411778 263860 411794
rect 204748 411722 204764 411778
rect 204820 411722 263788 411778
rect 263844 411722 263860 411778
rect 204748 411706 263860 411722
rect 334332 411778 579700 411794
rect 334332 411722 334348 411778
rect 334404 411722 579628 411778
rect 579684 411722 579700 411778
rect 334332 411706 579700 411722
rect 352700 411598 411588 411614
rect 352700 411542 352716 411598
rect 352772 411542 411516 411598
rect 411572 411542 411588 411598
rect 352700 411526 411588 411542
rect 334444 410698 579364 410714
rect 334444 410642 334460 410698
rect 334516 410642 579292 410698
rect 579348 410642 579364 410698
rect 334444 410626 579364 410642
rect 144268 409978 252884 409994
rect 144268 409922 144284 409978
rect 144340 409922 252812 409978
rect 252868 409922 252884 409978
rect 144268 409906 252884 409922
rect 401420 409978 534452 409994
rect 401420 409922 401436 409978
rect 401492 409922 534380 409978
rect 534436 409922 534452 409978
rect 401420 409906 534452 409922
rect 351020 409798 572924 409814
rect 351020 409742 351036 409798
rect 351092 409742 572924 409798
rect 351020 409726 572924 409742
rect 334444 409618 534340 409634
rect 334444 409562 334460 409618
rect 334516 409562 534268 409618
rect 534324 409562 534340 409618
rect 334444 409546 534340 409562
rect 572836 409454 572924 409726
rect 572836 409438 579364 409454
rect 572836 409382 579292 409438
rect 579348 409382 579364 409438
rect 572836 409366 579364 409382
rect 82668 409078 249524 409094
rect 82668 409022 82684 409078
rect 82740 409022 249452 409078
rect 249508 409022 249524 409078
rect 82668 409006 249524 409022
rect 144268 408358 263524 408374
rect 144268 408302 144284 408358
rect 144340 408302 263452 408358
rect 263508 408302 263524 408358
rect 144268 408286 263524 408302
rect 334444 408178 401508 408194
rect 334444 408122 334460 408178
rect 334516 408122 401436 408178
rect 401492 408122 401508 408178
rect 334444 408106 401508 408122
rect 334444 407458 428948 407474
rect 334444 407402 334460 407458
rect 334516 407402 428876 407458
rect 428932 407402 428948 407458
rect 334444 407386 428948 407402
rect 440956 407458 579924 407474
rect 440956 407402 440972 407458
rect 441028 407402 579924 407458
rect 440956 407386 579924 407402
rect 204972 407098 263972 407114
rect 204972 407042 204988 407098
rect 205044 407042 263900 407098
rect 263956 407042 263972 407098
rect 204972 407026 263972 407042
rect 579836 407098 579924 407386
rect 579836 407042 579852 407098
rect 579908 407042 579924 407098
rect 579836 407026 579924 407042
rect 191532 406918 263860 406934
rect 191532 406862 191548 406918
rect 191604 406862 263788 406918
rect 263844 406862 263860 406918
rect 191532 406846 263860 406862
rect 20620 406738 63044 406754
rect 20620 406682 20636 406738
rect 20692 406682 62972 406738
rect 63028 406682 63044 406738
rect 20620 406666 63044 406682
rect 82332 406738 125204 406754
rect 82332 406682 82348 406738
rect 82404 406682 125132 406738
rect 125188 406682 125204 406738
rect 82332 406666 125204 406682
rect 144380 406738 262292 406754
rect 144380 406682 144396 406738
rect 144452 406682 262220 406738
rect 262276 406682 262292 406738
rect 144380 406666 262292 406682
rect 336236 406738 411252 406754
rect 336236 406682 336252 406738
rect 336308 406682 411180 406738
rect 411236 406682 411252 406738
rect 336236 406666 411252 406682
rect -1916 406350 597980 406446
rect -1916 406294 -1820 406350
rect -1764 406294 -1696 406350
rect -1640 406294 -1572 406350
rect -1516 406294 -1448 406350
rect -1392 406294 9234 406350
rect 9290 406294 9358 406350
rect 9414 406294 9482 406350
rect 9538 406294 9606 406350
rect 9662 406294 39878 406350
rect 39934 406294 40002 406350
rect 40058 406294 70674 406350
rect 70730 406294 70798 406350
rect 70854 406294 70922 406350
rect 70978 406294 71046 406350
rect 71102 406294 101878 406350
rect 101934 406294 102002 406350
rect 102058 406294 132114 406350
rect 132170 406294 132238 406350
rect 132294 406294 132362 406350
rect 132418 406294 132486 406350
rect 132542 406294 162834 406350
rect 162890 406294 162958 406350
rect 163014 406294 163082 406350
rect 163138 406294 163206 406350
rect 163262 406294 163878 406350
rect 163934 406294 164002 406350
rect 164058 406294 193554 406350
rect 193610 406294 193678 406350
rect 193734 406294 193802 406350
rect 193858 406294 193926 406350
rect 193982 406294 224274 406350
rect 224330 406294 224398 406350
rect 224454 406294 224522 406350
rect 224578 406294 224646 406350
rect 224702 406294 225878 406350
rect 225934 406294 226002 406350
rect 226058 406294 254994 406350
rect 255050 406294 255118 406350
rect 255174 406294 255242 406350
rect 255298 406294 255366 406350
rect 255422 406294 287878 406350
rect 287934 406294 288002 406350
rect 288058 406294 318598 406350
rect 318654 406294 318722 406350
rect 318778 406294 347154 406350
rect 347210 406294 347278 406350
rect 347334 406294 347402 406350
rect 347458 406294 347526 406350
rect 347582 406294 371878 406350
rect 371934 406294 372002 406350
rect 372058 406294 377874 406350
rect 377930 406294 377998 406350
rect 378054 406294 378122 406350
rect 378178 406294 378246 406350
rect 378302 406294 408594 406350
rect 408650 406294 408718 406350
rect 408774 406294 408842 406350
rect 408898 406294 408966 406350
rect 409022 406294 433878 406350
rect 433934 406294 434002 406350
rect 434058 406294 470034 406350
rect 470090 406294 470158 406350
rect 470214 406294 470282 406350
rect 470338 406294 470406 406350
rect 470462 406294 495878 406350
rect 495934 406294 496002 406350
rect 496058 406294 531474 406350
rect 531530 406294 531598 406350
rect 531654 406294 531722 406350
rect 531778 406294 531846 406350
rect 531902 406294 557878 406350
rect 557934 406294 558002 406350
rect 558058 406294 562194 406350
rect 562250 406294 562318 406350
rect 562374 406294 562442 406350
rect 562498 406294 562566 406350
rect 562622 406294 592914 406350
rect 592970 406294 593038 406350
rect 593094 406294 593162 406350
rect 593218 406294 593286 406350
rect 593342 406294 597456 406350
rect 597512 406294 597580 406350
rect 597636 406294 597704 406350
rect 597760 406294 597828 406350
rect 597884 406294 597980 406350
rect -1916 406226 597980 406294
rect -1916 406170 -1820 406226
rect -1764 406170 -1696 406226
rect -1640 406170 -1572 406226
rect -1516 406170 -1448 406226
rect -1392 406170 9234 406226
rect 9290 406170 9358 406226
rect 9414 406170 9482 406226
rect 9538 406170 9606 406226
rect 9662 406170 39878 406226
rect 39934 406170 40002 406226
rect 40058 406170 70674 406226
rect 70730 406170 70798 406226
rect 70854 406170 70922 406226
rect 70978 406170 71046 406226
rect 71102 406170 101878 406226
rect 101934 406170 102002 406226
rect 102058 406170 132114 406226
rect 132170 406170 132238 406226
rect 132294 406170 132362 406226
rect 132418 406170 132486 406226
rect 132542 406170 162834 406226
rect 162890 406170 162958 406226
rect 163014 406170 163082 406226
rect 163138 406170 163206 406226
rect 163262 406170 163878 406226
rect 163934 406170 164002 406226
rect 164058 406170 193554 406226
rect 193610 406170 193678 406226
rect 193734 406170 193802 406226
rect 193858 406170 193926 406226
rect 193982 406170 224274 406226
rect 224330 406170 224398 406226
rect 224454 406170 224522 406226
rect 224578 406170 224646 406226
rect 224702 406170 225878 406226
rect 225934 406170 226002 406226
rect 226058 406170 254994 406226
rect 255050 406170 255118 406226
rect 255174 406170 255242 406226
rect 255298 406170 255366 406226
rect 255422 406170 287878 406226
rect 287934 406170 288002 406226
rect 288058 406170 318598 406226
rect 318654 406170 318722 406226
rect 318778 406170 347154 406226
rect 347210 406170 347278 406226
rect 347334 406170 347402 406226
rect 347458 406170 347526 406226
rect 347582 406170 371878 406226
rect 371934 406170 372002 406226
rect 372058 406170 377874 406226
rect 377930 406170 377998 406226
rect 378054 406170 378122 406226
rect 378178 406170 378246 406226
rect 378302 406170 408594 406226
rect 408650 406170 408718 406226
rect 408774 406170 408842 406226
rect 408898 406170 408966 406226
rect 409022 406170 433878 406226
rect 433934 406170 434002 406226
rect 434058 406170 470034 406226
rect 470090 406170 470158 406226
rect 470214 406170 470282 406226
rect 470338 406170 470406 406226
rect 470462 406170 495878 406226
rect 495934 406170 496002 406226
rect 496058 406170 531474 406226
rect 531530 406170 531598 406226
rect 531654 406170 531722 406226
rect 531778 406170 531846 406226
rect 531902 406170 557878 406226
rect 557934 406170 558002 406226
rect 558058 406170 562194 406226
rect 562250 406170 562318 406226
rect 562374 406170 562442 406226
rect 562498 406170 562566 406226
rect 562622 406170 592914 406226
rect 592970 406170 593038 406226
rect 593094 406170 593162 406226
rect 593218 406170 593286 406226
rect 593342 406170 597456 406226
rect 597512 406170 597580 406226
rect 597636 406170 597704 406226
rect 597760 406170 597828 406226
rect 597884 406170 597980 406226
rect -1916 406102 597980 406170
rect -1916 406046 -1820 406102
rect -1764 406046 -1696 406102
rect -1640 406046 -1572 406102
rect -1516 406046 -1448 406102
rect -1392 406046 9234 406102
rect 9290 406046 9358 406102
rect 9414 406046 9482 406102
rect 9538 406046 9606 406102
rect 9662 406046 39878 406102
rect 39934 406046 40002 406102
rect 40058 406046 70674 406102
rect 70730 406046 70798 406102
rect 70854 406046 70922 406102
rect 70978 406046 71046 406102
rect 71102 406046 101878 406102
rect 101934 406046 102002 406102
rect 102058 406046 132114 406102
rect 132170 406046 132238 406102
rect 132294 406046 132362 406102
rect 132418 406046 132486 406102
rect 132542 406046 162834 406102
rect 162890 406046 162958 406102
rect 163014 406046 163082 406102
rect 163138 406046 163206 406102
rect 163262 406046 163878 406102
rect 163934 406046 164002 406102
rect 164058 406046 193554 406102
rect 193610 406046 193678 406102
rect 193734 406046 193802 406102
rect 193858 406046 193926 406102
rect 193982 406046 224274 406102
rect 224330 406046 224398 406102
rect 224454 406046 224522 406102
rect 224578 406046 224646 406102
rect 224702 406046 225878 406102
rect 225934 406046 226002 406102
rect 226058 406046 254994 406102
rect 255050 406046 255118 406102
rect 255174 406046 255242 406102
rect 255298 406046 255366 406102
rect 255422 406046 287878 406102
rect 287934 406046 288002 406102
rect 288058 406046 318598 406102
rect 318654 406046 318722 406102
rect 318778 406046 347154 406102
rect 347210 406046 347278 406102
rect 347334 406046 347402 406102
rect 347458 406046 347526 406102
rect 347582 406046 371878 406102
rect 371934 406046 372002 406102
rect 372058 406046 377874 406102
rect 377930 406046 377998 406102
rect 378054 406046 378122 406102
rect 378178 406046 378246 406102
rect 378302 406046 408594 406102
rect 408650 406046 408718 406102
rect 408774 406046 408842 406102
rect 408898 406046 408966 406102
rect 409022 406046 433878 406102
rect 433934 406046 434002 406102
rect 434058 406046 470034 406102
rect 470090 406046 470158 406102
rect 470214 406046 470282 406102
rect 470338 406046 470406 406102
rect 470462 406046 495878 406102
rect 495934 406046 496002 406102
rect 496058 406046 531474 406102
rect 531530 406046 531598 406102
rect 531654 406046 531722 406102
rect 531778 406046 531846 406102
rect 531902 406046 557878 406102
rect 557934 406046 558002 406102
rect 558058 406046 562194 406102
rect 562250 406046 562318 406102
rect 562374 406046 562442 406102
rect 562498 406046 562566 406102
rect 562622 406046 592914 406102
rect 592970 406046 593038 406102
rect 593094 406046 593162 406102
rect 593218 406046 593286 406102
rect 593342 406046 597456 406102
rect 597512 406046 597580 406102
rect 597636 406046 597704 406102
rect 597760 406046 597828 406102
rect 597884 406046 597980 406102
rect -1916 405978 597980 406046
rect -1916 405922 -1820 405978
rect -1764 405922 -1696 405978
rect -1640 405922 -1572 405978
rect -1516 405922 -1448 405978
rect -1392 405922 9234 405978
rect 9290 405922 9358 405978
rect 9414 405922 9482 405978
rect 9538 405922 9606 405978
rect 9662 405922 39878 405978
rect 39934 405922 40002 405978
rect 40058 405922 70674 405978
rect 70730 405922 70798 405978
rect 70854 405922 70922 405978
rect 70978 405922 71046 405978
rect 71102 405922 101878 405978
rect 101934 405922 102002 405978
rect 102058 405922 132114 405978
rect 132170 405922 132238 405978
rect 132294 405922 132362 405978
rect 132418 405922 132486 405978
rect 132542 405922 162834 405978
rect 162890 405922 162958 405978
rect 163014 405922 163082 405978
rect 163138 405922 163206 405978
rect 163262 405922 163878 405978
rect 163934 405922 164002 405978
rect 164058 405922 193554 405978
rect 193610 405922 193678 405978
rect 193734 405922 193802 405978
rect 193858 405922 193926 405978
rect 193982 405922 224274 405978
rect 224330 405922 224398 405978
rect 224454 405922 224522 405978
rect 224578 405922 224646 405978
rect 224702 405922 225878 405978
rect 225934 405922 226002 405978
rect 226058 405922 254994 405978
rect 255050 405922 255118 405978
rect 255174 405922 255242 405978
rect 255298 405922 255366 405978
rect 255422 405922 287878 405978
rect 287934 405922 288002 405978
rect 288058 405922 318598 405978
rect 318654 405922 318722 405978
rect 318778 405922 347154 405978
rect 347210 405922 347278 405978
rect 347334 405922 347402 405978
rect 347458 405922 347526 405978
rect 347582 405922 371878 405978
rect 371934 405922 372002 405978
rect 372058 405922 377874 405978
rect 377930 405922 377998 405978
rect 378054 405922 378122 405978
rect 378178 405922 378246 405978
rect 378302 405922 408594 405978
rect 408650 405922 408718 405978
rect 408774 405922 408842 405978
rect 408898 405922 408966 405978
rect 409022 405922 433878 405978
rect 433934 405922 434002 405978
rect 434058 405922 470034 405978
rect 470090 405922 470158 405978
rect 470214 405922 470282 405978
rect 470338 405922 470406 405978
rect 470462 405922 495878 405978
rect 495934 405922 496002 405978
rect 496058 405922 531474 405978
rect 531530 405922 531598 405978
rect 531654 405922 531722 405978
rect 531778 405922 531846 405978
rect 531902 405922 557878 405978
rect 557934 405922 558002 405978
rect 558058 405922 562194 405978
rect 562250 405922 562318 405978
rect 562374 405922 562442 405978
rect 562498 405922 562566 405978
rect 562622 405922 592914 405978
rect 592970 405922 593038 405978
rect 593094 405922 593162 405978
rect 593218 405922 593286 405978
rect 593342 405922 597456 405978
rect 597512 405922 597580 405978
rect 597636 405922 597704 405978
rect 597760 405922 597828 405978
rect 597884 405922 597980 405978
rect -1916 405826 597980 405922
rect 189292 404758 262180 404774
rect 189292 404702 189308 404758
rect 189364 404702 262108 404758
rect 262164 404702 262180 404758
rect 189292 404686 262180 404702
rect 336012 404758 472180 404774
rect 336012 404702 336028 404758
rect 336084 404702 472108 404758
rect 472164 404702 472180 404758
rect 336012 404686 472180 404702
rect 189516 404578 260388 404594
rect 189516 404522 189532 404578
rect 189588 404522 260316 404578
rect 260372 404522 260388 404578
rect 189516 404506 260388 404522
rect 144268 404218 205060 404234
rect 144268 404162 144284 404218
rect 144340 404162 204988 404218
rect 205044 404162 205060 404218
rect 144268 404146 205060 404162
rect 189404 404038 263860 404054
rect 189404 403982 189420 404038
rect 189476 403982 263788 404038
rect 263844 403982 263860 404038
rect 189404 403966 263860 403982
rect 518236 404038 579812 404054
rect 518236 403982 518252 404038
rect 518308 403982 579812 404038
rect 518236 403966 579812 403982
rect 579724 403858 579812 403966
rect 579724 403802 579740 403858
rect 579796 403802 579812 403858
rect 579724 403786 579812 403802
rect 334444 403318 517316 403334
rect 334444 403262 334460 403318
rect 334516 403262 517244 403318
rect 517300 403262 517316 403318
rect 334444 403246 517316 403262
rect 199820 403138 263860 403154
rect 199820 403082 199836 403138
rect 199892 403082 263788 403138
rect 263844 403082 263860 403138
rect 199820 403066 263860 403082
rect 334444 403138 461204 403154
rect 334444 403082 334460 403138
rect 334516 403082 461132 403138
rect 461188 403082 461204 403138
rect 334444 403066 461204 403082
rect 523276 403138 579700 403154
rect 523276 403082 523292 403138
rect 523348 403082 579700 403138
rect 523276 403066 579700 403082
rect 204972 402958 263972 402974
rect 204972 402902 204988 402958
rect 205044 402902 263900 402958
rect 263956 402902 263972 402958
rect 204972 402886 263972 402902
rect 414076 402958 534340 402974
rect 414076 402902 414092 402958
rect 414148 402902 534268 402958
rect 534324 402902 534340 402958
rect 414076 402886 534340 402902
rect 579612 402598 579700 403066
rect 579612 402542 579628 402598
rect 579684 402542 579700 402598
rect 579612 402526 579700 402542
rect 126236 402418 199124 402434
rect 126236 402362 126252 402418
rect 126308 402362 199052 402418
rect 199108 402362 199124 402418
rect 126236 402346 199124 402362
rect 351020 402418 411140 402434
rect 351020 402362 351036 402418
rect 351092 402362 411068 402418
rect 411124 402362 411140 402418
rect 351020 402346 411140 402362
rect -1916 400350 597980 400446
rect -1916 400294 -860 400350
rect -804 400294 -736 400350
rect -680 400294 -612 400350
rect -556 400294 -488 400350
rect -432 400294 5514 400350
rect 5570 400294 5638 400350
rect 5694 400294 5762 400350
rect 5818 400294 5886 400350
rect 5942 400294 24518 400350
rect 24574 400294 24642 400350
rect 24698 400294 36234 400350
rect 36290 400294 36358 400350
rect 36414 400294 36482 400350
rect 36538 400294 36606 400350
rect 36662 400294 55238 400350
rect 55294 400294 55362 400350
rect 55418 400294 66954 400350
rect 67010 400294 67078 400350
rect 67134 400294 67202 400350
rect 67258 400294 67326 400350
rect 67382 400294 86518 400350
rect 86574 400294 86642 400350
rect 86698 400294 117238 400350
rect 117294 400294 117362 400350
rect 117418 400294 128394 400350
rect 128450 400294 128518 400350
rect 128574 400294 128642 400350
rect 128698 400294 128766 400350
rect 128822 400294 148518 400350
rect 148574 400294 148642 400350
rect 148698 400294 159114 400350
rect 159170 400294 159238 400350
rect 159294 400294 159362 400350
rect 159418 400294 159486 400350
rect 159542 400294 179238 400350
rect 179294 400294 179362 400350
rect 179418 400294 189834 400350
rect 189890 400294 189958 400350
rect 190014 400294 190082 400350
rect 190138 400294 190206 400350
rect 190262 400294 210518 400350
rect 210574 400294 210642 400350
rect 210698 400294 220554 400350
rect 220610 400294 220678 400350
rect 220734 400294 220802 400350
rect 220858 400294 220926 400350
rect 220982 400294 241238 400350
rect 241294 400294 241362 400350
rect 241418 400294 251274 400350
rect 251330 400294 251398 400350
rect 251454 400294 251522 400350
rect 251578 400294 251646 400350
rect 251702 400294 272518 400350
rect 272574 400294 272642 400350
rect 272698 400294 303238 400350
rect 303294 400294 303362 400350
rect 303418 400294 343434 400350
rect 343490 400294 343558 400350
rect 343614 400294 343682 400350
rect 343738 400294 343806 400350
rect 343862 400294 356518 400350
rect 356574 400294 356642 400350
rect 356698 400294 387238 400350
rect 387294 400294 387362 400350
rect 387418 400294 404874 400350
rect 404930 400294 404998 400350
rect 405054 400294 405122 400350
rect 405178 400294 405246 400350
rect 405302 400294 418518 400350
rect 418574 400294 418642 400350
rect 418698 400294 435594 400350
rect 435650 400294 435718 400350
rect 435774 400294 435842 400350
rect 435898 400294 435966 400350
rect 436022 400294 449238 400350
rect 449294 400294 449362 400350
rect 449418 400294 466314 400350
rect 466370 400294 466438 400350
rect 466494 400294 466562 400350
rect 466618 400294 466686 400350
rect 466742 400294 480518 400350
rect 480574 400294 480642 400350
rect 480698 400294 497034 400350
rect 497090 400294 497158 400350
rect 497214 400294 497282 400350
rect 497338 400294 497406 400350
rect 497462 400294 511238 400350
rect 511294 400294 511362 400350
rect 511418 400294 527754 400350
rect 527810 400294 527878 400350
rect 527934 400294 528002 400350
rect 528058 400294 528126 400350
rect 528182 400294 542518 400350
rect 542574 400294 542642 400350
rect 542698 400294 558474 400350
rect 558530 400294 558598 400350
rect 558654 400294 558722 400350
rect 558778 400294 558846 400350
rect 558902 400294 573238 400350
rect 573294 400294 573362 400350
rect 573418 400294 589194 400350
rect 589250 400294 589318 400350
rect 589374 400294 589442 400350
rect 589498 400294 589566 400350
rect 589622 400294 596496 400350
rect 596552 400294 596620 400350
rect 596676 400294 596744 400350
rect 596800 400294 596868 400350
rect 596924 400294 597980 400350
rect -1916 400226 597980 400294
rect -1916 400170 -860 400226
rect -804 400170 -736 400226
rect -680 400170 -612 400226
rect -556 400170 -488 400226
rect -432 400170 5514 400226
rect 5570 400170 5638 400226
rect 5694 400170 5762 400226
rect 5818 400170 5886 400226
rect 5942 400170 24518 400226
rect 24574 400170 24642 400226
rect 24698 400170 36234 400226
rect 36290 400170 36358 400226
rect 36414 400170 36482 400226
rect 36538 400170 36606 400226
rect 36662 400170 55238 400226
rect 55294 400170 55362 400226
rect 55418 400170 66954 400226
rect 67010 400170 67078 400226
rect 67134 400170 67202 400226
rect 67258 400170 67326 400226
rect 67382 400170 86518 400226
rect 86574 400170 86642 400226
rect 86698 400170 117238 400226
rect 117294 400170 117362 400226
rect 117418 400170 128394 400226
rect 128450 400170 128518 400226
rect 128574 400170 128642 400226
rect 128698 400170 128766 400226
rect 128822 400170 148518 400226
rect 148574 400170 148642 400226
rect 148698 400170 159114 400226
rect 159170 400170 159238 400226
rect 159294 400170 159362 400226
rect 159418 400170 159486 400226
rect 159542 400170 179238 400226
rect 179294 400170 179362 400226
rect 179418 400170 189834 400226
rect 189890 400170 189958 400226
rect 190014 400170 190082 400226
rect 190138 400170 190206 400226
rect 190262 400170 210518 400226
rect 210574 400170 210642 400226
rect 210698 400170 220554 400226
rect 220610 400170 220678 400226
rect 220734 400170 220802 400226
rect 220858 400170 220926 400226
rect 220982 400170 241238 400226
rect 241294 400170 241362 400226
rect 241418 400170 251274 400226
rect 251330 400170 251398 400226
rect 251454 400170 251522 400226
rect 251578 400170 251646 400226
rect 251702 400170 272518 400226
rect 272574 400170 272642 400226
rect 272698 400170 303238 400226
rect 303294 400170 303362 400226
rect 303418 400170 343434 400226
rect 343490 400170 343558 400226
rect 343614 400170 343682 400226
rect 343738 400170 343806 400226
rect 343862 400170 356518 400226
rect 356574 400170 356642 400226
rect 356698 400170 387238 400226
rect 387294 400170 387362 400226
rect 387418 400170 404874 400226
rect 404930 400170 404998 400226
rect 405054 400170 405122 400226
rect 405178 400170 405246 400226
rect 405302 400170 418518 400226
rect 418574 400170 418642 400226
rect 418698 400170 435594 400226
rect 435650 400170 435718 400226
rect 435774 400170 435842 400226
rect 435898 400170 435966 400226
rect 436022 400170 449238 400226
rect 449294 400170 449362 400226
rect 449418 400170 466314 400226
rect 466370 400170 466438 400226
rect 466494 400170 466562 400226
rect 466618 400170 466686 400226
rect 466742 400170 480518 400226
rect 480574 400170 480642 400226
rect 480698 400170 497034 400226
rect 497090 400170 497158 400226
rect 497214 400170 497282 400226
rect 497338 400170 497406 400226
rect 497462 400170 511238 400226
rect 511294 400170 511362 400226
rect 511418 400170 527754 400226
rect 527810 400170 527878 400226
rect 527934 400170 528002 400226
rect 528058 400170 528126 400226
rect 528182 400170 542518 400226
rect 542574 400170 542642 400226
rect 542698 400170 558474 400226
rect 558530 400170 558598 400226
rect 558654 400170 558722 400226
rect 558778 400170 558846 400226
rect 558902 400170 573238 400226
rect 573294 400170 573362 400226
rect 573418 400170 589194 400226
rect 589250 400170 589318 400226
rect 589374 400170 589442 400226
rect 589498 400170 589566 400226
rect 589622 400170 596496 400226
rect 596552 400170 596620 400226
rect 596676 400170 596744 400226
rect 596800 400170 596868 400226
rect 596924 400170 597980 400226
rect -1916 400102 597980 400170
rect -1916 400046 -860 400102
rect -804 400046 -736 400102
rect -680 400046 -612 400102
rect -556 400046 -488 400102
rect -432 400046 5514 400102
rect 5570 400046 5638 400102
rect 5694 400046 5762 400102
rect 5818 400046 5886 400102
rect 5942 400046 24518 400102
rect 24574 400046 24642 400102
rect 24698 400046 36234 400102
rect 36290 400046 36358 400102
rect 36414 400046 36482 400102
rect 36538 400046 36606 400102
rect 36662 400046 55238 400102
rect 55294 400046 55362 400102
rect 55418 400046 66954 400102
rect 67010 400046 67078 400102
rect 67134 400046 67202 400102
rect 67258 400046 67326 400102
rect 67382 400046 86518 400102
rect 86574 400046 86642 400102
rect 86698 400046 117238 400102
rect 117294 400046 117362 400102
rect 117418 400046 128394 400102
rect 128450 400046 128518 400102
rect 128574 400046 128642 400102
rect 128698 400046 128766 400102
rect 128822 400046 148518 400102
rect 148574 400046 148642 400102
rect 148698 400046 159114 400102
rect 159170 400046 159238 400102
rect 159294 400046 159362 400102
rect 159418 400046 159486 400102
rect 159542 400046 179238 400102
rect 179294 400046 179362 400102
rect 179418 400046 189834 400102
rect 189890 400046 189958 400102
rect 190014 400046 190082 400102
rect 190138 400046 190206 400102
rect 190262 400046 210518 400102
rect 210574 400046 210642 400102
rect 210698 400046 220554 400102
rect 220610 400046 220678 400102
rect 220734 400046 220802 400102
rect 220858 400046 220926 400102
rect 220982 400046 241238 400102
rect 241294 400046 241362 400102
rect 241418 400046 251274 400102
rect 251330 400046 251398 400102
rect 251454 400046 251522 400102
rect 251578 400046 251646 400102
rect 251702 400046 272518 400102
rect 272574 400046 272642 400102
rect 272698 400046 303238 400102
rect 303294 400046 303362 400102
rect 303418 400046 343434 400102
rect 343490 400046 343558 400102
rect 343614 400046 343682 400102
rect 343738 400046 343806 400102
rect 343862 400046 356518 400102
rect 356574 400046 356642 400102
rect 356698 400046 387238 400102
rect 387294 400046 387362 400102
rect 387418 400046 404874 400102
rect 404930 400046 404998 400102
rect 405054 400046 405122 400102
rect 405178 400046 405246 400102
rect 405302 400046 418518 400102
rect 418574 400046 418642 400102
rect 418698 400046 435594 400102
rect 435650 400046 435718 400102
rect 435774 400046 435842 400102
rect 435898 400046 435966 400102
rect 436022 400046 449238 400102
rect 449294 400046 449362 400102
rect 449418 400046 466314 400102
rect 466370 400046 466438 400102
rect 466494 400046 466562 400102
rect 466618 400046 466686 400102
rect 466742 400046 480518 400102
rect 480574 400046 480642 400102
rect 480698 400046 497034 400102
rect 497090 400046 497158 400102
rect 497214 400046 497282 400102
rect 497338 400046 497406 400102
rect 497462 400046 511238 400102
rect 511294 400046 511362 400102
rect 511418 400046 527754 400102
rect 527810 400046 527878 400102
rect 527934 400046 528002 400102
rect 528058 400046 528126 400102
rect 528182 400046 542518 400102
rect 542574 400046 542642 400102
rect 542698 400046 558474 400102
rect 558530 400046 558598 400102
rect 558654 400046 558722 400102
rect 558778 400046 558846 400102
rect 558902 400046 573238 400102
rect 573294 400046 573362 400102
rect 573418 400046 589194 400102
rect 589250 400046 589318 400102
rect 589374 400046 589442 400102
rect 589498 400046 589566 400102
rect 589622 400046 596496 400102
rect 596552 400046 596620 400102
rect 596676 400046 596744 400102
rect 596800 400046 596868 400102
rect 596924 400046 597980 400102
rect -1916 399978 597980 400046
rect -1916 399922 -860 399978
rect -804 399922 -736 399978
rect -680 399922 -612 399978
rect -556 399922 -488 399978
rect -432 399922 5514 399978
rect 5570 399922 5638 399978
rect 5694 399922 5762 399978
rect 5818 399922 5886 399978
rect 5942 399922 24518 399978
rect 24574 399922 24642 399978
rect 24698 399922 36234 399978
rect 36290 399922 36358 399978
rect 36414 399922 36482 399978
rect 36538 399922 36606 399978
rect 36662 399922 55238 399978
rect 55294 399922 55362 399978
rect 55418 399922 66954 399978
rect 67010 399922 67078 399978
rect 67134 399922 67202 399978
rect 67258 399922 67326 399978
rect 67382 399922 86518 399978
rect 86574 399922 86642 399978
rect 86698 399922 117238 399978
rect 117294 399922 117362 399978
rect 117418 399922 128394 399978
rect 128450 399922 128518 399978
rect 128574 399922 128642 399978
rect 128698 399922 128766 399978
rect 128822 399922 148518 399978
rect 148574 399922 148642 399978
rect 148698 399922 159114 399978
rect 159170 399922 159238 399978
rect 159294 399922 159362 399978
rect 159418 399922 159486 399978
rect 159542 399922 179238 399978
rect 179294 399922 179362 399978
rect 179418 399922 189834 399978
rect 189890 399922 189958 399978
rect 190014 399922 190082 399978
rect 190138 399922 190206 399978
rect 190262 399922 210518 399978
rect 210574 399922 210642 399978
rect 210698 399922 220554 399978
rect 220610 399922 220678 399978
rect 220734 399922 220802 399978
rect 220858 399922 220926 399978
rect 220982 399922 241238 399978
rect 241294 399922 241362 399978
rect 241418 399922 251274 399978
rect 251330 399922 251398 399978
rect 251454 399922 251522 399978
rect 251578 399922 251646 399978
rect 251702 399922 272518 399978
rect 272574 399922 272642 399978
rect 272698 399922 303238 399978
rect 303294 399922 303362 399978
rect 303418 399922 343434 399978
rect 343490 399922 343558 399978
rect 343614 399922 343682 399978
rect 343738 399922 343806 399978
rect 343862 399922 356518 399978
rect 356574 399922 356642 399978
rect 356698 399922 387238 399978
rect 387294 399922 387362 399978
rect 387418 399922 404874 399978
rect 404930 399922 404998 399978
rect 405054 399922 405122 399978
rect 405178 399922 405246 399978
rect 405302 399922 418518 399978
rect 418574 399922 418642 399978
rect 418698 399922 435594 399978
rect 435650 399922 435718 399978
rect 435774 399922 435842 399978
rect 435898 399922 435966 399978
rect 436022 399922 449238 399978
rect 449294 399922 449362 399978
rect 449418 399922 466314 399978
rect 466370 399922 466438 399978
rect 466494 399922 466562 399978
rect 466618 399922 466686 399978
rect 466742 399922 480518 399978
rect 480574 399922 480642 399978
rect 480698 399922 497034 399978
rect 497090 399922 497158 399978
rect 497214 399922 497282 399978
rect 497338 399922 497406 399978
rect 497462 399922 511238 399978
rect 511294 399922 511362 399978
rect 511418 399922 527754 399978
rect 527810 399922 527878 399978
rect 527934 399922 528002 399978
rect 528058 399922 528126 399978
rect 528182 399922 542518 399978
rect 542574 399922 542642 399978
rect 542698 399922 558474 399978
rect 558530 399922 558598 399978
rect 558654 399922 558722 399978
rect 558778 399922 558846 399978
rect 558902 399922 573238 399978
rect 573294 399922 573362 399978
rect 573418 399922 589194 399978
rect 589250 399922 589318 399978
rect 589374 399922 589442 399978
rect 589498 399922 589566 399978
rect 589622 399922 596496 399978
rect 596552 399922 596620 399978
rect 596676 399922 596744 399978
rect 596800 399922 596868 399978
rect 596924 399922 597980 399978
rect -1916 399826 597980 399922
rect 136092 399718 263860 399734
rect 136092 399662 136108 399718
rect 136164 399662 263788 399718
rect 263844 399662 263860 399718
rect 136092 399646 263860 399662
rect 334444 399718 406660 399734
rect 334444 399662 334460 399718
rect 334516 399662 406588 399718
rect 406644 399662 406660 399718
rect 334444 399646 406660 399662
rect 189516 399538 262180 399554
rect 189516 399482 189532 399538
rect 189588 399482 262108 399538
rect 262164 399482 262180 399538
rect 189516 399466 262180 399482
rect 401420 398998 458740 399014
rect 401420 398942 401436 398998
rect 401492 398942 458668 398998
rect 458724 398942 458740 398998
rect 401420 398926 458740 398942
rect 82332 398098 263860 398114
rect 82332 398042 82348 398098
rect 82404 398042 263788 398098
rect 263844 398042 263860 398098
rect 82332 398026 263860 398042
rect 334444 398098 411252 398114
rect 334444 398042 334460 398098
rect 334516 398042 411180 398098
rect 411236 398042 411252 398098
rect 334444 398026 411252 398042
rect 334444 397918 401284 397934
rect 334444 397862 334460 397918
rect 334516 397862 401212 397918
rect 401268 397862 401284 397918
rect 334444 397846 401284 397862
rect 401308 397378 458964 397394
rect 401308 397322 401324 397378
rect 401380 397322 458892 397378
rect 458948 397322 458964 397378
rect 401308 397306 458964 397322
rect 125116 396478 263860 396494
rect 125116 396422 125132 396478
rect 125188 396422 263788 396478
rect 263844 396422 263860 396478
rect 125116 396406 263860 396422
rect 334444 396478 457060 396494
rect 334444 396422 334460 396478
rect 334516 396422 456988 396478
rect 457044 396422 457060 396478
rect 334444 396406 457060 396422
rect 199036 396298 263972 396314
rect 199036 396242 199052 396298
rect 199108 396242 263900 396298
rect 263956 396242 263972 396298
rect 199036 396226 263972 396242
rect 334332 396298 401508 396314
rect 334332 396242 334348 396298
rect 334404 396242 401436 396298
rect 401492 396242 401508 396298
rect 334332 396226 401508 396242
rect 334444 394678 455604 394694
rect 334444 394622 334460 394678
rect 334516 394622 455532 394678
rect 455588 394622 455604 394678
rect 334444 394606 455604 394622
rect 334444 394498 410804 394514
rect 334444 394442 334460 394498
rect 334516 394442 410732 394498
rect 410788 394442 410804 394498
rect 334444 394426 410804 394442
rect 135196 393058 263860 393074
rect 135196 393002 135212 393058
rect 135268 393002 263788 393058
rect 263844 393002 263860 393058
rect 135196 392986 263860 393002
rect 334444 393058 401396 393074
rect 334444 393002 334460 393058
rect 334516 393002 401324 393058
rect 401380 393002 401396 393058
rect 334444 392986 401396 393002
rect 334444 391618 455604 391634
rect 334444 391562 334460 391618
rect 334516 391562 455532 391618
rect 455588 391562 455604 391618
rect 334444 391546 455604 391562
rect 62956 391438 263860 391454
rect 62956 391382 62972 391438
rect 63028 391382 263788 391438
rect 263844 391382 263860 391438
rect 62956 391366 263860 391382
rect 350348 391438 579700 391454
rect 350348 391382 350364 391438
rect 350420 391382 579700 391438
rect 350348 391366 579700 391382
rect 579612 391078 579700 391366
rect 579612 391022 579628 391078
rect 579684 391022 579700 391078
rect 579612 391006 579700 391022
rect -1916 388389 597980 388446
rect -1916 388350 39836 388389
rect -1916 388294 -1820 388350
rect -1764 388294 -1696 388350
rect -1640 388294 -1572 388350
rect -1516 388294 -1448 388350
rect -1392 388294 9234 388350
rect 9290 388294 9358 388350
rect 9414 388294 9482 388350
rect 9538 388294 9606 388350
rect 9662 388333 39836 388350
rect 39892 388333 39940 388389
rect 39996 388333 40044 388389
rect 40100 388350 101836 388389
rect 40100 388333 70674 388350
rect 9662 388294 70674 388333
rect 70730 388294 70798 388350
rect 70854 388294 70922 388350
rect 70978 388294 71046 388350
rect 71102 388333 101836 388350
rect 101892 388333 101940 388389
rect 101996 388333 102044 388389
rect 102100 388350 163836 388389
rect 102100 388333 132114 388350
rect 71102 388294 132114 388333
rect 132170 388294 132238 388350
rect 132294 388294 132362 388350
rect 132418 388294 132486 388350
rect 132542 388294 162834 388350
rect 162890 388294 162958 388350
rect 163014 388294 163082 388350
rect 163138 388294 163206 388350
rect 163262 388333 163836 388350
rect 163892 388333 163940 388389
rect 163996 388333 164044 388389
rect 164100 388350 225836 388389
rect 164100 388333 193554 388350
rect 163262 388294 193554 388333
rect 193610 388294 193678 388350
rect 193734 388294 193802 388350
rect 193858 388294 193926 388350
rect 193982 388294 224274 388350
rect 224330 388294 224398 388350
rect 224454 388294 224522 388350
rect 224578 388294 224646 388350
rect 224702 388333 225836 388350
rect 225892 388333 225940 388389
rect 225996 388333 226044 388389
rect 226100 388350 371836 388389
rect 226100 388333 254994 388350
rect 224702 388294 254994 388333
rect 255050 388294 255118 388350
rect 255174 388294 255242 388350
rect 255298 388294 255366 388350
rect 255422 388294 287878 388350
rect 287934 388294 288002 388350
rect 288058 388294 318598 388350
rect 318654 388294 318722 388350
rect 318778 388294 347154 388350
rect 347210 388294 347278 388350
rect 347334 388294 347402 388350
rect 347458 388294 347526 388350
rect 347582 388333 371836 388350
rect 371892 388333 371940 388389
rect 371996 388333 372044 388389
rect 372100 388350 433836 388389
rect 372100 388333 377874 388350
rect 347582 388294 377874 388333
rect 377930 388294 377998 388350
rect 378054 388294 378122 388350
rect 378178 388294 378246 388350
rect 378302 388294 408594 388350
rect 408650 388294 408718 388350
rect 408774 388294 408842 388350
rect 408898 388294 408966 388350
rect 409022 388333 433836 388350
rect 433892 388333 433940 388389
rect 433996 388333 434044 388389
rect 434100 388350 495836 388389
rect 434100 388333 439314 388350
rect 409022 388294 439314 388333
rect 439370 388294 439438 388350
rect 439494 388294 439562 388350
rect 439618 388294 439686 388350
rect 439742 388294 470034 388350
rect 470090 388294 470158 388350
rect 470214 388294 470282 388350
rect 470338 388294 470406 388350
rect 470462 388333 495836 388350
rect 495892 388333 495940 388389
rect 495996 388333 496044 388389
rect 496100 388350 557836 388389
rect 496100 388333 500754 388350
rect 470462 388294 500754 388333
rect 500810 388294 500878 388350
rect 500934 388294 501002 388350
rect 501058 388294 501126 388350
rect 501182 388294 531474 388350
rect 531530 388294 531598 388350
rect 531654 388294 531722 388350
rect 531778 388294 531846 388350
rect 531902 388333 557836 388350
rect 557892 388333 557940 388389
rect 557996 388333 558044 388389
rect 558100 388350 597980 388389
rect 558100 388333 562194 388350
rect 531902 388294 562194 388333
rect 562250 388294 562318 388350
rect 562374 388294 562442 388350
rect 562498 388294 562566 388350
rect 562622 388294 592914 388350
rect 592970 388294 593038 388350
rect 593094 388294 593162 388350
rect 593218 388294 593286 388350
rect 593342 388294 597456 388350
rect 597512 388294 597580 388350
rect 597636 388294 597704 388350
rect 597760 388294 597828 388350
rect 597884 388294 597980 388350
rect -1916 388226 597980 388294
rect -1916 388170 -1820 388226
rect -1764 388170 -1696 388226
rect -1640 388170 -1572 388226
rect -1516 388170 -1448 388226
rect -1392 388170 9234 388226
rect 9290 388170 9358 388226
rect 9414 388170 9482 388226
rect 9538 388170 9606 388226
rect 9662 388170 70674 388226
rect 70730 388170 70798 388226
rect 70854 388170 70922 388226
rect 70978 388170 71046 388226
rect 71102 388170 132114 388226
rect 132170 388170 132238 388226
rect 132294 388170 132362 388226
rect 132418 388170 132486 388226
rect 132542 388170 162834 388226
rect 162890 388170 162958 388226
rect 163014 388170 163082 388226
rect 163138 388170 163206 388226
rect 163262 388170 193554 388226
rect 193610 388170 193678 388226
rect 193734 388170 193802 388226
rect 193858 388170 193926 388226
rect 193982 388170 224274 388226
rect 224330 388170 224398 388226
rect 224454 388170 224522 388226
rect 224578 388170 224646 388226
rect 224702 388170 254994 388226
rect 255050 388170 255118 388226
rect 255174 388170 255242 388226
rect 255298 388170 255366 388226
rect 255422 388170 287878 388226
rect 287934 388170 288002 388226
rect 288058 388170 318598 388226
rect 318654 388170 318722 388226
rect 318778 388170 347154 388226
rect 347210 388170 347278 388226
rect 347334 388170 347402 388226
rect 347458 388170 347526 388226
rect 347582 388170 377874 388226
rect 377930 388170 377998 388226
rect 378054 388170 378122 388226
rect 378178 388170 378246 388226
rect 378302 388170 408594 388226
rect 408650 388170 408718 388226
rect 408774 388170 408842 388226
rect 408898 388170 408966 388226
rect 409022 388170 439314 388226
rect 439370 388170 439438 388226
rect 439494 388170 439562 388226
rect 439618 388170 439686 388226
rect 439742 388170 470034 388226
rect 470090 388170 470158 388226
rect 470214 388170 470282 388226
rect 470338 388170 470406 388226
rect 470462 388170 500754 388226
rect 500810 388170 500878 388226
rect 500934 388170 501002 388226
rect 501058 388170 501126 388226
rect 501182 388170 531474 388226
rect 531530 388170 531598 388226
rect 531654 388170 531722 388226
rect 531778 388170 531846 388226
rect 531902 388170 562194 388226
rect 562250 388170 562318 388226
rect 562374 388170 562442 388226
rect 562498 388170 562566 388226
rect 562622 388170 592914 388226
rect 592970 388170 593038 388226
rect 593094 388170 593162 388226
rect 593218 388170 593286 388226
rect 593342 388170 597456 388226
rect 597512 388170 597580 388226
rect 597636 388170 597704 388226
rect 597760 388170 597828 388226
rect 597884 388170 597980 388226
rect -1916 388102 597980 388170
rect -1916 388046 -1820 388102
rect -1764 388046 -1696 388102
rect -1640 388046 -1572 388102
rect -1516 388046 -1448 388102
rect -1392 388046 9234 388102
rect 9290 388046 9358 388102
rect 9414 388046 9482 388102
rect 9538 388046 9606 388102
rect 9662 388046 70674 388102
rect 70730 388046 70798 388102
rect 70854 388046 70922 388102
rect 70978 388046 71046 388102
rect 71102 388046 132114 388102
rect 132170 388046 132238 388102
rect 132294 388046 132362 388102
rect 132418 388046 132486 388102
rect 132542 388046 162834 388102
rect 162890 388046 162958 388102
rect 163014 388046 163082 388102
rect 163138 388046 163206 388102
rect 163262 388046 193554 388102
rect 193610 388046 193678 388102
rect 193734 388046 193802 388102
rect 193858 388046 193926 388102
rect 193982 388046 224274 388102
rect 224330 388046 224398 388102
rect 224454 388046 224522 388102
rect 224578 388046 224646 388102
rect 224702 388046 254994 388102
rect 255050 388046 255118 388102
rect 255174 388046 255242 388102
rect 255298 388046 255366 388102
rect 255422 388046 287878 388102
rect 287934 388046 288002 388102
rect 288058 388046 318598 388102
rect 318654 388046 318722 388102
rect 318778 388046 347154 388102
rect 347210 388046 347278 388102
rect 347334 388046 347402 388102
rect 347458 388046 347526 388102
rect 347582 388046 377874 388102
rect 377930 388046 377998 388102
rect 378054 388046 378122 388102
rect 378178 388046 378246 388102
rect 378302 388046 408594 388102
rect 408650 388046 408718 388102
rect 408774 388046 408842 388102
rect 408898 388046 408966 388102
rect 409022 388046 439314 388102
rect 439370 388046 439438 388102
rect 439494 388046 439562 388102
rect 439618 388046 439686 388102
rect 439742 388046 470034 388102
rect 470090 388046 470158 388102
rect 470214 388046 470282 388102
rect 470338 388046 470406 388102
rect 470462 388046 500754 388102
rect 500810 388046 500878 388102
rect 500934 388046 501002 388102
rect 501058 388046 501126 388102
rect 501182 388046 531474 388102
rect 531530 388046 531598 388102
rect 531654 388046 531722 388102
rect 531778 388046 531846 388102
rect 531902 388046 562194 388102
rect 562250 388046 562318 388102
rect 562374 388046 562442 388102
rect 562498 388046 562566 388102
rect 562622 388046 592914 388102
rect 592970 388046 593038 388102
rect 593094 388046 593162 388102
rect 593218 388046 593286 388102
rect 593342 388046 597456 388102
rect 597512 388046 597580 388102
rect 597636 388046 597704 388102
rect 597760 388046 597828 388102
rect 597884 388046 597980 388102
rect -1916 387978 597980 388046
rect -1916 387922 -1820 387978
rect -1764 387922 -1696 387978
rect -1640 387922 -1572 387978
rect -1516 387922 -1448 387978
rect -1392 387922 9234 387978
rect 9290 387922 9358 387978
rect 9414 387922 9482 387978
rect 9538 387922 9606 387978
rect 9662 387922 70674 387978
rect 70730 387922 70798 387978
rect 70854 387922 70922 387978
rect 70978 387922 71046 387978
rect 71102 387922 132114 387978
rect 132170 387922 132238 387978
rect 132294 387922 132362 387978
rect 132418 387922 132486 387978
rect 132542 387922 162834 387978
rect 162890 387922 162958 387978
rect 163014 387922 163082 387978
rect 163138 387922 163206 387978
rect 163262 387922 193554 387978
rect 193610 387922 193678 387978
rect 193734 387922 193802 387978
rect 193858 387922 193926 387978
rect 193982 387922 224274 387978
rect 224330 387922 224398 387978
rect 224454 387922 224522 387978
rect 224578 387922 224646 387978
rect 224702 387922 254994 387978
rect 255050 387922 255118 387978
rect 255174 387922 255242 387978
rect 255298 387922 255366 387978
rect 255422 387922 287878 387978
rect 287934 387922 288002 387978
rect 288058 387922 318598 387978
rect 318654 387922 318722 387978
rect 318778 387922 347154 387978
rect 347210 387922 347278 387978
rect 347334 387922 347402 387978
rect 347458 387922 347526 387978
rect 347582 387922 377874 387978
rect 377930 387922 377998 387978
rect 378054 387922 378122 387978
rect 378178 387922 378246 387978
rect 378302 387922 408594 387978
rect 408650 387922 408718 387978
rect 408774 387922 408842 387978
rect 408898 387922 408966 387978
rect 409022 387922 439314 387978
rect 439370 387922 439438 387978
rect 439494 387922 439562 387978
rect 439618 387922 439686 387978
rect 439742 387922 470034 387978
rect 470090 387922 470158 387978
rect 470214 387922 470282 387978
rect 470338 387922 470406 387978
rect 470462 387922 500754 387978
rect 500810 387922 500878 387978
rect 500934 387922 501002 387978
rect 501058 387922 501126 387978
rect 501182 387922 531474 387978
rect 531530 387922 531598 387978
rect 531654 387922 531722 387978
rect 531778 387922 531846 387978
rect 531902 387922 562194 387978
rect 562250 387922 562318 387978
rect 562374 387922 562442 387978
rect 562498 387922 562566 387978
rect 562622 387922 592914 387978
rect 592970 387922 593038 387978
rect 593094 387922 593162 387978
rect 593218 387922 593286 387978
rect 593342 387922 597456 387978
rect 597512 387922 597580 387978
rect 597636 387922 597704 387978
rect 597760 387922 597828 387978
rect 597884 387922 597980 387978
rect -1916 387826 597980 387922
rect -1916 382350 597980 382446
rect -1916 382294 -860 382350
rect -804 382294 -736 382350
rect -680 382294 -612 382350
rect -556 382294 -488 382350
rect -432 382294 5514 382350
rect 5570 382294 5638 382350
rect 5694 382294 5762 382350
rect 5818 382294 5886 382350
rect 5942 382294 36234 382350
rect 36290 382294 36358 382350
rect 36414 382294 36482 382350
rect 36538 382294 36606 382350
rect 36662 382294 66954 382350
rect 67010 382294 67078 382350
rect 67134 382294 67202 382350
rect 67258 382294 67326 382350
rect 67382 382294 97674 382350
rect 97730 382294 97798 382350
rect 97854 382294 97922 382350
rect 97978 382294 98046 382350
rect 98102 382294 128394 382350
rect 128450 382294 128518 382350
rect 128574 382294 128642 382350
rect 128698 382294 128766 382350
rect 128822 382294 159114 382350
rect 159170 382294 159238 382350
rect 159294 382294 159362 382350
rect 159418 382294 159486 382350
rect 159542 382294 189834 382350
rect 189890 382294 189958 382350
rect 190014 382294 190082 382350
rect 190138 382294 190206 382350
rect 190262 382294 220554 382350
rect 220610 382294 220678 382350
rect 220734 382294 220802 382350
rect 220858 382294 220926 382350
rect 220982 382294 251274 382350
rect 251330 382294 251398 382350
rect 251454 382294 251522 382350
rect 251578 382294 251646 382350
rect 251702 382294 272518 382350
rect 272574 382294 272642 382350
rect 272698 382294 303238 382350
rect 303294 382294 303362 382350
rect 303418 382294 343434 382350
rect 343490 382294 343558 382350
rect 343614 382294 343682 382350
rect 343738 382294 343806 382350
rect 343862 382294 374154 382350
rect 374210 382294 374278 382350
rect 374334 382294 374402 382350
rect 374458 382294 374526 382350
rect 374582 382294 404874 382350
rect 404930 382294 404998 382350
rect 405054 382294 405122 382350
rect 405178 382294 405246 382350
rect 405302 382294 435594 382350
rect 435650 382294 435718 382350
rect 435774 382294 435842 382350
rect 435898 382294 435966 382350
rect 436022 382294 466314 382350
rect 466370 382294 466438 382350
rect 466494 382294 466562 382350
rect 466618 382294 466686 382350
rect 466742 382294 497034 382350
rect 497090 382294 497158 382350
rect 497214 382294 497282 382350
rect 497338 382294 497406 382350
rect 497462 382294 527754 382350
rect 527810 382294 527878 382350
rect 527934 382294 528002 382350
rect 528058 382294 528126 382350
rect 528182 382294 558474 382350
rect 558530 382294 558598 382350
rect 558654 382294 558722 382350
rect 558778 382294 558846 382350
rect 558902 382294 589194 382350
rect 589250 382294 589318 382350
rect 589374 382294 589442 382350
rect 589498 382294 589566 382350
rect 589622 382294 596496 382350
rect 596552 382294 596620 382350
rect 596676 382294 596744 382350
rect 596800 382294 596868 382350
rect 596924 382294 597980 382350
rect -1916 382226 597980 382294
rect -1916 382170 -860 382226
rect -804 382170 -736 382226
rect -680 382170 -612 382226
rect -556 382170 -488 382226
rect -432 382170 5514 382226
rect 5570 382170 5638 382226
rect 5694 382170 5762 382226
rect 5818 382170 5886 382226
rect 5942 382170 36234 382226
rect 36290 382170 36358 382226
rect 36414 382170 36482 382226
rect 36538 382170 36606 382226
rect 36662 382170 66954 382226
rect 67010 382170 67078 382226
rect 67134 382170 67202 382226
rect 67258 382170 67326 382226
rect 67382 382170 97674 382226
rect 97730 382170 97798 382226
rect 97854 382170 97922 382226
rect 97978 382170 98046 382226
rect 98102 382170 128394 382226
rect 128450 382170 128518 382226
rect 128574 382170 128642 382226
rect 128698 382170 128766 382226
rect 128822 382170 159114 382226
rect 159170 382170 159238 382226
rect 159294 382170 159362 382226
rect 159418 382170 159486 382226
rect 159542 382170 189834 382226
rect 189890 382170 189958 382226
rect 190014 382170 190082 382226
rect 190138 382170 190206 382226
rect 190262 382170 220554 382226
rect 220610 382170 220678 382226
rect 220734 382170 220802 382226
rect 220858 382170 220926 382226
rect 220982 382170 251274 382226
rect 251330 382170 251398 382226
rect 251454 382170 251522 382226
rect 251578 382170 251646 382226
rect 251702 382170 272518 382226
rect 272574 382170 272642 382226
rect 272698 382170 303238 382226
rect 303294 382170 303362 382226
rect 303418 382170 343434 382226
rect 343490 382170 343558 382226
rect 343614 382170 343682 382226
rect 343738 382170 343806 382226
rect 343862 382170 374154 382226
rect 374210 382170 374278 382226
rect 374334 382170 374402 382226
rect 374458 382170 374526 382226
rect 374582 382170 404874 382226
rect 404930 382170 404998 382226
rect 405054 382170 405122 382226
rect 405178 382170 405246 382226
rect 405302 382170 435594 382226
rect 435650 382170 435718 382226
rect 435774 382170 435842 382226
rect 435898 382170 435966 382226
rect 436022 382170 466314 382226
rect 466370 382170 466438 382226
rect 466494 382170 466562 382226
rect 466618 382170 466686 382226
rect 466742 382170 497034 382226
rect 497090 382170 497158 382226
rect 497214 382170 497282 382226
rect 497338 382170 497406 382226
rect 497462 382170 527754 382226
rect 527810 382170 527878 382226
rect 527934 382170 528002 382226
rect 528058 382170 528126 382226
rect 528182 382170 558474 382226
rect 558530 382170 558598 382226
rect 558654 382170 558722 382226
rect 558778 382170 558846 382226
rect 558902 382170 589194 382226
rect 589250 382170 589318 382226
rect 589374 382170 589442 382226
rect 589498 382170 589566 382226
rect 589622 382170 596496 382226
rect 596552 382170 596620 382226
rect 596676 382170 596744 382226
rect 596800 382170 596868 382226
rect 596924 382170 597980 382226
rect -1916 382102 597980 382170
rect -1916 382046 -860 382102
rect -804 382046 -736 382102
rect -680 382046 -612 382102
rect -556 382046 -488 382102
rect -432 382046 5514 382102
rect 5570 382046 5638 382102
rect 5694 382046 5762 382102
rect 5818 382046 5886 382102
rect 5942 382046 36234 382102
rect 36290 382046 36358 382102
rect 36414 382046 36482 382102
rect 36538 382046 36606 382102
rect 36662 382046 66954 382102
rect 67010 382046 67078 382102
rect 67134 382046 67202 382102
rect 67258 382046 67326 382102
rect 67382 382046 97674 382102
rect 97730 382046 97798 382102
rect 97854 382046 97922 382102
rect 97978 382046 98046 382102
rect 98102 382046 128394 382102
rect 128450 382046 128518 382102
rect 128574 382046 128642 382102
rect 128698 382046 128766 382102
rect 128822 382046 159114 382102
rect 159170 382046 159238 382102
rect 159294 382046 159362 382102
rect 159418 382046 159486 382102
rect 159542 382046 189834 382102
rect 189890 382046 189958 382102
rect 190014 382046 190082 382102
rect 190138 382046 190206 382102
rect 190262 382046 220554 382102
rect 220610 382046 220678 382102
rect 220734 382046 220802 382102
rect 220858 382046 220926 382102
rect 220982 382046 251274 382102
rect 251330 382046 251398 382102
rect 251454 382046 251522 382102
rect 251578 382046 251646 382102
rect 251702 382046 272518 382102
rect 272574 382046 272642 382102
rect 272698 382046 303238 382102
rect 303294 382046 303362 382102
rect 303418 382046 343434 382102
rect 343490 382046 343558 382102
rect 343614 382046 343682 382102
rect 343738 382046 343806 382102
rect 343862 382046 374154 382102
rect 374210 382046 374278 382102
rect 374334 382046 374402 382102
rect 374458 382046 374526 382102
rect 374582 382046 404874 382102
rect 404930 382046 404998 382102
rect 405054 382046 405122 382102
rect 405178 382046 405246 382102
rect 405302 382046 435594 382102
rect 435650 382046 435718 382102
rect 435774 382046 435842 382102
rect 435898 382046 435966 382102
rect 436022 382046 466314 382102
rect 466370 382046 466438 382102
rect 466494 382046 466562 382102
rect 466618 382046 466686 382102
rect 466742 382046 497034 382102
rect 497090 382046 497158 382102
rect 497214 382046 497282 382102
rect 497338 382046 497406 382102
rect 497462 382046 527754 382102
rect 527810 382046 527878 382102
rect 527934 382046 528002 382102
rect 528058 382046 528126 382102
rect 528182 382046 558474 382102
rect 558530 382046 558598 382102
rect 558654 382046 558722 382102
rect 558778 382046 558846 382102
rect 558902 382046 589194 382102
rect 589250 382046 589318 382102
rect 589374 382046 589442 382102
rect 589498 382046 589566 382102
rect 589622 382046 596496 382102
rect 596552 382046 596620 382102
rect 596676 382046 596744 382102
rect 596800 382046 596868 382102
rect 596924 382046 597980 382102
rect -1916 381978 597980 382046
rect -1916 381922 -860 381978
rect -804 381922 -736 381978
rect -680 381922 -612 381978
rect -556 381922 -488 381978
rect -432 381922 5514 381978
rect 5570 381922 5638 381978
rect 5694 381922 5762 381978
rect 5818 381922 5886 381978
rect 5942 381922 36234 381978
rect 36290 381922 36358 381978
rect 36414 381922 36482 381978
rect 36538 381922 36606 381978
rect 36662 381922 66954 381978
rect 67010 381922 67078 381978
rect 67134 381922 67202 381978
rect 67258 381922 67326 381978
rect 67382 381922 97674 381978
rect 97730 381922 97798 381978
rect 97854 381922 97922 381978
rect 97978 381922 98046 381978
rect 98102 381922 128394 381978
rect 128450 381922 128518 381978
rect 128574 381922 128642 381978
rect 128698 381922 128766 381978
rect 128822 381922 159114 381978
rect 159170 381922 159238 381978
rect 159294 381922 159362 381978
rect 159418 381922 159486 381978
rect 159542 381922 189834 381978
rect 189890 381922 189958 381978
rect 190014 381922 190082 381978
rect 190138 381922 190206 381978
rect 190262 381922 220554 381978
rect 220610 381922 220678 381978
rect 220734 381922 220802 381978
rect 220858 381922 220926 381978
rect 220982 381922 251274 381978
rect 251330 381922 251398 381978
rect 251454 381922 251522 381978
rect 251578 381922 251646 381978
rect 251702 381922 272518 381978
rect 272574 381922 272642 381978
rect 272698 381922 303238 381978
rect 303294 381922 303362 381978
rect 303418 381922 343434 381978
rect 343490 381922 343558 381978
rect 343614 381922 343682 381978
rect 343738 381922 343806 381978
rect 343862 381922 374154 381978
rect 374210 381922 374278 381978
rect 374334 381922 374402 381978
rect 374458 381922 374526 381978
rect 374582 381922 404874 381978
rect 404930 381922 404998 381978
rect 405054 381922 405122 381978
rect 405178 381922 405246 381978
rect 405302 381922 435594 381978
rect 435650 381922 435718 381978
rect 435774 381922 435842 381978
rect 435898 381922 435966 381978
rect 436022 381922 466314 381978
rect 466370 381922 466438 381978
rect 466494 381922 466562 381978
rect 466618 381922 466686 381978
rect 466742 381922 497034 381978
rect 497090 381922 497158 381978
rect 497214 381922 497282 381978
rect 497338 381922 497406 381978
rect 497462 381922 527754 381978
rect 527810 381922 527878 381978
rect 527934 381922 528002 381978
rect 528058 381922 528126 381978
rect 528182 381922 558474 381978
rect 558530 381922 558598 381978
rect 558654 381922 558722 381978
rect 558778 381922 558846 381978
rect 558902 381922 589194 381978
rect 589250 381922 589318 381978
rect 589374 381922 589442 381978
rect 589498 381922 589566 381978
rect 589622 381922 596496 381978
rect 596552 381922 596620 381978
rect 596676 381922 596744 381978
rect 596800 381922 596868 381978
rect 596924 381922 597980 381978
rect -1916 381826 597980 381922
rect -1916 370350 597980 370446
rect -1916 370294 -1820 370350
rect -1764 370294 -1696 370350
rect -1640 370294 -1572 370350
rect -1516 370294 -1448 370350
rect -1392 370294 9234 370350
rect 9290 370294 9358 370350
rect 9414 370294 9482 370350
rect 9538 370294 9606 370350
rect 9662 370294 70674 370350
rect 70730 370294 70798 370350
rect 70854 370294 70922 370350
rect 70978 370294 71046 370350
rect 71102 370294 132114 370350
rect 132170 370294 132238 370350
rect 132294 370294 132362 370350
rect 132418 370294 132486 370350
rect 132542 370294 162834 370350
rect 162890 370294 162958 370350
rect 163014 370294 163082 370350
rect 163138 370294 163206 370350
rect 163262 370294 193554 370350
rect 193610 370294 193678 370350
rect 193734 370294 193802 370350
rect 193858 370294 193926 370350
rect 193982 370294 224274 370350
rect 224330 370294 224398 370350
rect 224454 370294 224522 370350
rect 224578 370294 224646 370350
rect 224702 370294 254994 370350
rect 255050 370294 255118 370350
rect 255174 370294 255242 370350
rect 255298 370294 255366 370350
rect 255422 370294 287878 370350
rect 287934 370294 288002 370350
rect 288058 370294 318598 370350
rect 318654 370294 318722 370350
rect 318778 370294 347154 370350
rect 347210 370294 347278 370350
rect 347334 370294 347402 370350
rect 347458 370294 347526 370350
rect 347582 370294 377874 370350
rect 377930 370294 377998 370350
rect 378054 370294 378122 370350
rect 378178 370294 378246 370350
rect 378302 370294 408594 370350
rect 408650 370294 408718 370350
rect 408774 370294 408842 370350
rect 408898 370294 408966 370350
rect 409022 370294 439314 370350
rect 439370 370294 439438 370350
rect 439494 370294 439562 370350
rect 439618 370294 439686 370350
rect 439742 370294 470034 370350
rect 470090 370294 470158 370350
rect 470214 370294 470282 370350
rect 470338 370294 470406 370350
rect 470462 370294 500754 370350
rect 500810 370294 500878 370350
rect 500934 370294 501002 370350
rect 501058 370294 501126 370350
rect 501182 370294 531474 370350
rect 531530 370294 531598 370350
rect 531654 370294 531722 370350
rect 531778 370294 531846 370350
rect 531902 370294 562194 370350
rect 562250 370294 562318 370350
rect 562374 370294 562442 370350
rect 562498 370294 562566 370350
rect 562622 370294 592914 370350
rect 592970 370294 593038 370350
rect 593094 370294 593162 370350
rect 593218 370294 593286 370350
rect 593342 370294 597456 370350
rect 597512 370294 597580 370350
rect 597636 370294 597704 370350
rect 597760 370294 597828 370350
rect 597884 370294 597980 370350
rect -1916 370226 597980 370294
rect -1916 370170 -1820 370226
rect -1764 370170 -1696 370226
rect -1640 370170 -1572 370226
rect -1516 370170 -1448 370226
rect -1392 370170 9234 370226
rect 9290 370170 9358 370226
rect 9414 370170 9482 370226
rect 9538 370170 9606 370226
rect 9662 370170 70674 370226
rect 70730 370170 70798 370226
rect 70854 370170 70922 370226
rect 70978 370170 71046 370226
rect 71102 370170 132114 370226
rect 132170 370170 132238 370226
rect 132294 370170 132362 370226
rect 132418 370170 132486 370226
rect 132542 370170 162834 370226
rect 162890 370170 162958 370226
rect 163014 370170 163082 370226
rect 163138 370170 163206 370226
rect 163262 370170 193554 370226
rect 193610 370170 193678 370226
rect 193734 370170 193802 370226
rect 193858 370170 193926 370226
rect 193982 370170 224274 370226
rect 224330 370170 224398 370226
rect 224454 370170 224522 370226
rect 224578 370170 224646 370226
rect 224702 370170 254994 370226
rect 255050 370170 255118 370226
rect 255174 370170 255242 370226
rect 255298 370170 255366 370226
rect 255422 370170 287878 370226
rect 287934 370170 288002 370226
rect 288058 370170 318598 370226
rect 318654 370170 318722 370226
rect 318778 370170 347154 370226
rect 347210 370170 347278 370226
rect 347334 370170 347402 370226
rect 347458 370170 347526 370226
rect 347582 370170 377874 370226
rect 377930 370170 377998 370226
rect 378054 370170 378122 370226
rect 378178 370170 378246 370226
rect 378302 370170 408594 370226
rect 408650 370170 408718 370226
rect 408774 370170 408842 370226
rect 408898 370170 408966 370226
rect 409022 370170 439314 370226
rect 439370 370170 439438 370226
rect 439494 370170 439562 370226
rect 439618 370170 439686 370226
rect 439742 370170 470034 370226
rect 470090 370170 470158 370226
rect 470214 370170 470282 370226
rect 470338 370170 470406 370226
rect 470462 370170 500754 370226
rect 500810 370170 500878 370226
rect 500934 370170 501002 370226
rect 501058 370170 501126 370226
rect 501182 370170 531474 370226
rect 531530 370170 531598 370226
rect 531654 370170 531722 370226
rect 531778 370170 531846 370226
rect 531902 370170 562194 370226
rect 562250 370170 562318 370226
rect 562374 370170 562442 370226
rect 562498 370170 562566 370226
rect 562622 370170 592914 370226
rect 592970 370170 593038 370226
rect 593094 370170 593162 370226
rect 593218 370170 593286 370226
rect 593342 370170 597456 370226
rect 597512 370170 597580 370226
rect 597636 370170 597704 370226
rect 597760 370170 597828 370226
rect 597884 370170 597980 370226
rect -1916 370102 597980 370170
rect -1916 370046 -1820 370102
rect -1764 370046 -1696 370102
rect -1640 370046 -1572 370102
rect -1516 370046 -1448 370102
rect -1392 370046 9234 370102
rect 9290 370046 9358 370102
rect 9414 370046 9482 370102
rect 9538 370046 9606 370102
rect 9662 370046 70674 370102
rect 70730 370046 70798 370102
rect 70854 370046 70922 370102
rect 70978 370046 71046 370102
rect 71102 370046 132114 370102
rect 132170 370046 132238 370102
rect 132294 370046 132362 370102
rect 132418 370046 132486 370102
rect 132542 370046 162834 370102
rect 162890 370046 162958 370102
rect 163014 370046 163082 370102
rect 163138 370046 163206 370102
rect 163262 370046 193554 370102
rect 193610 370046 193678 370102
rect 193734 370046 193802 370102
rect 193858 370046 193926 370102
rect 193982 370046 224274 370102
rect 224330 370046 224398 370102
rect 224454 370046 224522 370102
rect 224578 370046 224646 370102
rect 224702 370046 254994 370102
rect 255050 370046 255118 370102
rect 255174 370046 255242 370102
rect 255298 370046 255366 370102
rect 255422 370046 287878 370102
rect 287934 370046 288002 370102
rect 288058 370046 318598 370102
rect 318654 370046 318722 370102
rect 318778 370046 347154 370102
rect 347210 370046 347278 370102
rect 347334 370046 347402 370102
rect 347458 370046 347526 370102
rect 347582 370046 377874 370102
rect 377930 370046 377998 370102
rect 378054 370046 378122 370102
rect 378178 370046 378246 370102
rect 378302 370046 408594 370102
rect 408650 370046 408718 370102
rect 408774 370046 408842 370102
rect 408898 370046 408966 370102
rect 409022 370046 439314 370102
rect 439370 370046 439438 370102
rect 439494 370046 439562 370102
rect 439618 370046 439686 370102
rect 439742 370046 470034 370102
rect 470090 370046 470158 370102
rect 470214 370046 470282 370102
rect 470338 370046 470406 370102
rect 470462 370046 500754 370102
rect 500810 370046 500878 370102
rect 500934 370046 501002 370102
rect 501058 370046 501126 370102
rect 501182 370046 531474 370102
rect 531530 370046 531598 370102
rect 531654 370046 531722 370102
rect 531778 370046 531846 370102
rect 531902 370046 562194 370102
rect 562250 370046 562318 370102
rect 562374 370046 562442 370102
rect 562498 370046 562566 370102
rect 562622 370046 592914 370102
rect 592970 370046 593038 370102
rect 593094 370046 593162 370102
rect 593218 370046 593286 370102
rect 593342 370046 597456 370102
rect 597512 370046 597580 370102
rect 597636 370046 597704 370102
rect 597760 370046 597828 370102
rect 597884 370046 597980 370102
rect -1916 369978 597980 370046
rect -1916 369922 -1820 369978
rect -1764 369922 -1696 369978
rect -1640 369922 -1572 369978
rect -1516 369922 -1448 369978
rect -1392 369922 9234 369978
rect 9290 369922 9358 369978
rect 9414 369922 9482 369978
rect 9538 369922 9606 369978
rect 9662 369922 70674 369978
rect 70730 369922 70798 369978
rect 70854 369922 70922 369978
rect 70978 369922 71046 369978
rect 71102 369922 132114 369978
rect 132170 369922 132238 369978
rect 132294 369922 132362 369978
rect 132418 369922 132486 369978
rect 132542 369922 162834 369978
rect 162890 369922 162958 369978
rect 163014 369922 163082 369978
rect 163138 369922 163206 369978
rect 163262 369922 193554 369978
rect 193610 369922 193678 369978
rect 193734 369922 193802 369978
rect 193858 369922 193926 369978
rect 193982 369922 224274 369978
rect 224330 369922 224398 369978
rect 224454 369922 224522 369978
rect 224578 369922 224646 369978
rect 224702 369922 254994 369978
rect 255050 369922 255118 369978
rect 255174 369922 255242 369978
rect 255298 369922 255366 369978
rect 255422 369922 287878 369978
rect 287934 369922 288002 369978
rect 288058 369922 318598 369978
rect 318654 369922 318722 369978
rect 318778 369922 347154 369978
rect 347210 369922 347278 369978
rect 347334 369922 347402 369978
rect 347458 369922 347526 369978
rect 347582 369922 377874 369978
rect 377930 369922 377998 369978
rect 378054 369922 378122 369978
rect 378178 369922 378246 369978
rect 378302 369922 408594 369978
rect 408650 369922 408718 369978
rect 408774 369922 408842 369978
rect 408898 369922 408966 369978
rect 409022 369922 439314 369978
rect 439370 369922 439438 369978
rect 439494 369922 439562 369978
rect 439618 369922 439686 369978
rect 439742 369922 470034 369978
rect 470090 369922 470158 369978
rect 470214 369922 470282 369978
rect 470338 369922 470406 369978
rect 470462 369922 500754 369978
rect 500810 369922 500878 369978
rect 500934 369922 501002 369978
rect 501058 369922 501126 369978
rect 501182 369922 531474 369978
rect 531530 369922 531598 369978
rect 531654 369922 531722 369978
rect 531778 369922 531846 369978
rect 531902 369922 562194 369978
rect 562250 369922 562318 369978
rect 562374 369922 562442 369978
rect 562498 369922 562566 369978
rect 562622 369922 592914 369978
rect 592970 369922 593038 369978
rect 593094 369922 593162 369978
rect 593218 369922 593286 369978
rect 593342 369922 597456 369978
rect 597512 369922 597580 369978
rect 597636 369922 597704 369978
rect 597760 369922 597828 369978
rect 597884 369922 597980 369978
rect -1916 369826 597980 369922
rect -1916 364350 597980 364446
rect -1916 364294 -860 364350
rect -804 364294 -736 364350
rect -680 364294 -612 364350
rect -556 364294 -488 364350
rect -432 364294 5514 364350
rect 5570 364294 5638 364350
rect 5694 364294 5762 364350
rect 5818 364294 5886 364350
rect 5942 364294 36234 364350
rect 36290 364294 36358 364350
rect 36414 364294 36482 364350
rect 36538 364294 36606 364350
rect 36662 364294 66954 364350
rect 67010 364294 67078 364350
rect 67134 364294 67202 364350
rect 67258 364294 67326 364350
rect 67382 364294 97674 364350
rect 97730 364294 97798 364350
rect 97854 364294 97922 364350
rect 97978 364294 98046 364350
rect 98102 364294 128394 364350
rect 128450 364294 128518 364350
rect 128574 364294 128642 364350
rect 128698 364294 128766 364350
rect 128822 364294 159114 364350
rect 159170 364294 159238 364350
rect 159294 364294 159362 364350
rect 159418 364294 159486 364350
rect 159542 364294 189834 364350
rect 189890 364294 189958 364350
rect 190014 364294 190082 364350
rect 190138 364294 190206 364350
rect 190262 364294 220554 364350
rect 220610 364294 220678 364350
rect 220734 364294 220802 364350
rect 220858 364294 220926 364350
rect 220982 364294 251274 364350
rect 251330 364294 251398 364350
rect 251454 364294 251522 364350
rect 251578 364294 251646 364350
rect 251702 364294 272518 364350
rect 272574 364294 272642 364350
rect 272698 364294 303238 364350
rect 303294 364294 303362 364350
rect 303418 364294 343434 364350
rect 343490 364294 343558 364350
rect 343614 364294 343682 364350
rect 343738 364294 343806 364350
rect 343862 364294 374154 364350
rect 374210 364294 374278 364350
rect 374334 364294 374402 364350
rect 374458 364294 374526 364350
rect 374582 364294 404874 364350
rect 404930 364294 404998 364350
rect 405054 364294 405122 364350
rect 405178 364294 405246 364350
rect 405302 364294 435594 364350
rect 435650 364294 435718 364350
rect 435774 364294 435842 364350
rect 435898 364294 435966 364350
rect 436022 364294 466314 364350
rect 466370 364294 466438 364350
rect 466494 364294 466562 364350
rect 466618 364294 466686 364350
rect 466742 364294 497034 364350
rect 497090 364294 497158 364350
rect 497214 364294 497282 364350
rect 497338 364294 497406 364350
rect 497462 364294 527754 364350
rect 527810 364294 527878 364350
rect 527934 364294 528002 364350
rect 528058 364294 528126 364350
rect 528182 364294 558474 364350
rect 558530 364294 558598 364350
rect 558654 364294 558722 364350
rect 558778 364294 558846 364350
rect 558902 364294 589194 364350
rect 589250 364294 589318 364350
rect 589374 364294 589442 364350
rect 589498 364294 589566 364350
rect 589622 364294 596496 364350
rect 596552 364294 596620 364350
rect 596676 364294 596744 364350
rect 596800 364294 596868 364350
rect 596924 364294 597980 364350
rect -1916 364226 597980 364294
rect -1916 364170 -860 364226
rect -804 364170 -736 364226
rect -680 364170 -612 364226
rect -556 364170 -488 364226
rect -432 364170 5514 364226
rect 5570 364170 5638 364226
rect 5694 364170 5762 364226
rect 5818 364170 5886 364226
rect 5942 364170 36234 364226
rect 36290 364170 36358 364226
rect 36414 364170 36482 364226
rect 36538 364170 36606 364226
rect 36662 364170 66954 364226
rect 67010 364170 67078 364226
rect 67134 364170 67202 364226
rect 67258 364170 67326 364226
rect 67382 364170 97674 364226
rect 97730 364170 97798 364226
rect 97854 364170 97922 364226
rect 97978 364170 98046 364226
rect 98102 364170 128394 364226
rect 128450 364170 128518 364226
rect 128574 364170 128642 364226
rect 128698 364170 128766 364226
rect 128822 364170 159114 364226
rect 159170 364170 159238 364226
rect 159294 364170 159362 364226
rect 159418 364170 159486 364226
rect 159542 364170 189834 364226
rect 189890 364170 189958 364226
rect 190014 364170 190082 364226
rect 190138 364170 190206 364226
rect 190262 364170 220554 364226
rect 220610 364170 220678 364226
rect 220734 364170 220802 364226
rect 220858 364170 220926 364226
rect 220982 364170 251274 364226
rect 251330 364170 251398 364226
rect 251454 364170 251522 364226
rect 251578 364170 251646 364226
rect 251702 364170 272518 364226
rect 272574 364170 272642 364226
rect 272698 364170 303238 364226
rect 303294 364170 303362 364226
rect 303418 364170 343434 364226
rect 343490 364170 343558 364226
rect 343614 364170 343682 364226
rect 343738 364170 343806 364226
rect 343862 364170 374154 364226
rect 374210 364170 374278 364226
rect 374334 364170 374402 364226
rect 374458 364170 374526 364226
rect 374582 364170 404874 364226
rect 404930 364170 404998 364226
rect 405054 364170 405122 364226
rect 405178 364170 405246 364226
rect 405302 364170 435594 364226
rect 435650 364170 435718 364226
rect 435774 364170 435842 364226
rect 435898 364170 435966 364226
rect 436022 364170 466314 364226
rect 466370 364170 466438 364226
rect 466494 364170 466562 364226
rect 466618 364170 466686 364226
rect 466742 364170 497034 364226
rect 497090 364170 497158 364226
rect 497214 364170 497282 364226
rect 497338 364170 497406 364226
rect 497462 364170 527754 364226
rect 527810 364170 527878 364226
rect 527934 364170 528002 364226
rect 528058 364170 528126 364226
rect 528182 364170 558474 364226
rect 558530 364170 558598 364226
rect 558654 364170 558722 364226
rect 558778 364170 558846 364226
rect 558902 364170 589194 364226
rect 589250 364170 589318 364226
rect 589374 364170 589442 364226
rect 589498 364170 589566 364226
rect 589622 364170 596496 364226
rect 596552 364170 596620 364226
rect 596676 364170 596744 364226
rect 596800 364170 596868 364226
rect 596924 364170 597980 364226
rect -1916 364102 597980 364170
rect -1916 364046 -860 364102
rect -804 364046 -736 364102
rect -680 364046 -612 364102
rect -556 364046 -488 364102
rect -432 364046 5514 364102
rect 5570 364046 5638 364102
rect 5694 364046 5762 364102
rect 5818 364046 5886 364102
rect 5942 364046 36234 364102
rect 36290 364046 36358 364102
rect 36414 364046 36482 364102
rect 36538 364046 36606 364102
rect 36662 364046 66954 364102
rect 67010 364046 67078 364102
rect 67134 364046 67202 364102
rect 67258 364046 67326 364102
rect 67382 364046 97674 364102
rect 97730 364046 97798 364102
rect 97854 364046 97922 364102
rect 97978 364046 98046 364102
rect 98102 364046 128394 364102
rect 128450 364046 128518 364102
rect 128574 364046 128642 364102
rect 128698 364046 128766 364102
rect 128822 364046 159114 364102
rect 159170 364046 159238 364102
rect 159294 364046 159362 364102
rect 159418 364046 159486 364102
rect 159542 364046 189834 364102
rect 189890 364046 189958 364102
rect 190014 364046 190082 364102
rect 190138 364046 190206 364102
rect 190262 364046 220554 364102
rect 220610 364046 220678 364102
rect 220734 364046 220802 364102
rect 220858 364046 220926 364102
rect 220982 364046 251274 364102
rect 251330 364046 251398 364102
rect 251454 364046 251522 364102
rect 251578 364046 251646 364102
rect 251702 364046 272518 364102
rect 272574 364046 272642 364102
rect 272698 364046 303238 364102
rect 303294 364046 303362 364102
rect 303418 364046 343434 364102
rect 343490 364046 343558 364102
rect 343614 364046 343682 364102
rect 343738 364046 343806 364102
rect 343862 364046 374154 364102
rect 374210 364046 374278 364102
rect 374334 364046 374402 364102
rect 374458 364046 374526 364102
rect 374582 364046 404874 364102
rect 404930 364046 404998 364102
rect 405054 364046 405122 364102
rect 405178 364046 405246 364102
rect 405302 364046 435594 364102
rect 435650 364046 435718 364102
rect 435774 364046 435842 364102
rect 435898 364046 435966 364102
rect 436022 364046 466314 364102
rect 466370 364046 466438 364102
rect 466494 364046 466562 364102
rect 466618 364046 466686 364102
rect 466742 364046 497034 364102
rect 497090 364046 497158 364102
rect 497214 364046 497282 364102
rect 497338 364046 497406 364102
rect 497462 364046 527754 364102
rect 527810 364046 527878 364102
rect 527934 364046 528002 364102
rect 528058 364046 528126 364102
rect 528182 364046 558474 364102
rect 558530 364046 558598 364102
rect 558654 364046 558722 364102
rect 558778 364046 558846 364102
rect 558902 364046 589194 364102
rect 589250 364046 589318 364102
rect 589374 364046 589442 364102
rect 589498 364046 589566 364102
rect 589622 364046 596496 364102
rect 596552 364046 596620 364102
rect 596676 364046 596744 364102
rect 596800 364046 596868 364102
rect 596924 364046 597980 364102
rect -1916 363978 597980 364046
rect -1916 363922 -860 363978
rect -804 363922 -736 363978
rect -680 363922 -612 363978
rect -556 363922 -488 363978
rect -432 363922 5514 363978
rect 5570 363922 5638 363978
rect 5694 363922 5762 363978
rect 5818 363922 5886 363978
rect 5942 363922 36234 363978
rect 36290 363922 36358 363978
rect 36414 363922 36482 363978
rect 36538 363922 36606 363978
rect 36662 363922 66954 363978
rect 67010 363922 67078 363978
rect 67134 363922 67202 363978
rect 67258 363922 67326 363978
rect 67382 363922 97674 363978
rect 97730 363922 97798 363978
rect 97854 363922 97922 363978
rect 97978 363922 98046 363978
rect 98102 363922 128394 363978
rect 128450 363922 128518 363978
rect 128574 363922 128642 363978
rect 128698 363922 128766 363978
rect 128822 363922 159114 363978
rect 159170 363922 159238 363978
rect 159294 363922 159362 363978
rect 159418 363922 159486 363978
rect 159542 363922 189834 363978
rect 189890 363922 189958 363978
rect 190014 363922 190082 363978
rect 190138 363922 190206 363978
rect 190262 363922 220554 363978
rect 220610 363922 220678 363978
rect 220734 363922 220802 363978
rect 220858 363922 220926 363978
rect 220982 363922 251274 363978
rect 251330 363922 251398 363978
rect 251454 363922 251522 363978
rect 251578 363922 251646 363978
rect 251702 363922 272518 363978
rect 272574 363922 272642 363978
rect 272698 363922 303238 363978
rect 303294 363922 303362 363978
rect 303418 363922 343434 363978
rect 343490 363922 343558 363978
rect 343614 363922 343682 363978
rect 343738 363922 343806 363978
rect 343862 363922 374154 363978
rect 374210 363922 374278 363978
rect 374334 363922 374402 363978
rect 374458 363922 374526 363978
rect 374582 363922 404874 363978
rect 404930 363922 404998 363978
rect 405054 363922 405122 363978
rect 405178 363922 405246 363978
rect 405302 363922 435594 363978
rect 435650 363922 435718 363978
rect 435774 363922 435842 363978
rect 435898 363922 435966 363978
rect 436022 363922 466314 363978
rect 466370 363922 466438 363978
rect 466494 363922 466562 363978
rect 466618 363922 466686 363978
rect 466742 363922 497034 363978
rect 497090 363922 497158 363978
rect 497214 363922 497282 363978
rect 497338 363922 497406 363978
rect 497462 363922 527754 363978
rect 527810 363922 527878 363978
rect 527934 363922 528002 363978
rect 528058 363922 528126 363978
rect 528182 363922 558474 363978
rect 558530 363922 558598 363978
rect 558654 363922 558722 363978
rect 558778 363922 558846 363978
rect 558902 363922 589194 363978
rect 589250 363922 589318 363978
rect 589374 363922 589442 363978
rect 589498 363922 589566 363978
rect 589622 363922 596496 363978
rect 596552 363922 596620 363978
rect 596676 363922 596744 363978
rect 596800 363922 596868 363978
rect 596924 363922 597980 363978
rect -1916 363826 597980 363922
rect -1916 352350 597980 352446
rect -1916 352294 -1820 352350
rect -1764 352294 -1696 352350
rect -1640 352294 -1572 352350
rect -1516 352294 -1448 352350
rect -1392 352294 9234 352350
rect 9290 352294 9358 352350
rect 9414 352294 9482 352350
rect 9538 352294 9606 352350
rect 9662 352294 39878 352350
rect 39934 352294 40002 352350
rect 40058 352294 70674 352350
rect 70730 352294 70798 352350
rect 70854 352294 70922 352350
rect 70978 352294 71046 352350
rect 71102 352294 101878 352350
rect 101934 352294 102002 352350
rect 102058 352294 132114 352350
rect 132170 352294 132238 352350
rect 132294 352294 132362 352350
rect 132418 352294 132486 352350
rect 132542 352294 162834 352350
rect 162890 352294 162958 352350
rect 163014 352294 163082 352350
rect 163138 352294 163206 352350
rect 163262 352294 163878 352350
rect 163934 352294 164002 352350
rect 164058 352294 193554 352350
rect 193610 352294 193678 352350
rect 193734 352294 193802 352350
rect 193858 352294 193926 352350
rect 193982 352294 224274 352350
rect 224330 352294 224398 352350
rect 224454 352294 224522 352350
rect 224578 352294 224646 352350
rect 224702 352294 225878 352350
rect 225934 352294 226002 352350
rect 226058 352294 254994 352350
rect 255050 352294 255118 352350
rect 255174 352294 255242 352350
rect 255298 352294 255366 352350
rect 255422 352294 287878 352350
rect 287934 352294 288002 352350
rect 288058 352294 318598 352350
rect 318654 352294 318722 352350
rect 318778 352294 347154 352350
rect 347210 352294 347278 352350
rect 347334 352294 347402 352350
rect 347458 352294 347526 352350
rect 347582 352294 371878 352350
rect 371934 352294 372002 352350
rect 372058 352294 377874 352350
rect 377930 352294 377998 352350
rect 378054 352294 378122 352350
rect 378178 352294 378246 352350
rect 378302 352294 408594 352350
rect 408650 352294 408718 352350
rect 408774 352294 408842 352350
rect 408898 352294 408966 352350
rect 409022 352294 433878 352350
rect 433934 352294 434002 352350
rect 434058 352294 439314 352350
rect 439370 352294 439438 352350
rect 439494 352294 439562 352350
rect 439618 352294 439686 352350
rect 439742 352294 470034 352350
rect 470090 352294 470158 352350
rect 470214 352294 470282 352350
rect 470338 352294 470406 352350
rect 470462 352294 495878 352350
rect 495934 352294 496002 352350
rect 496058 352294 500754 352350
rect 500810 352294 500878 352350
rect 500934 352294 501002 352350
rect 501058 352294 501126 352350
rect 501182 352294 531474 352350
rect 531530 352294 531598 352350
rect 531654 352294 531722 352350
rect 531778 352294 531846 352350
rect 531902 352294 557878 352350
rect 557934 352294 558002 352350
rect 558058 352294 562194 352350
rect 562250 352294 562318 352350
rect 562374 352294 562442 352350
rect 562498 352294 562566 352350
rect 562622 352294 592914 352350
rect 592970 352294 593038 352350
rect 593094 352294 593162 352350
rect 593218 352294 593286 352350
rect 593342 352294 597456 352350
rect 597512 352294 597580 352350
rect 597636 352294 597704 352350
rect 597760 352294 597828 352350
rect 597884 352294 597980 352350
rect -1916 352226 597980 352294
rect -1916 352170 -1820 352226
rect -1764 352170 -1696 352226
rect -1640 352170 -1572 352226
rect -1516 352170 -1448 352226
rect -1392 352170 9234 352226
rect 9290 352170 9358 352226
rect 9414 352170 9482 352226
rect 9538 352170 9606 352226
rect 9662 352170 39878 352226
rect 39934 352170 40002 352226
rect 40058 352170 70674 352226
rect 70730 352170 70798 352226
rect 70854 352170 70922 352226
rect 70978 352170 71046 352226
rect 71102 352170 101878 352226
rect 101934 352170 102002 352226
rect 102058 352170 132114 352226
rect 132170 352170 132238 352226
rect 132294 352170 132362 352226
rect 132418 352170 132486 352226
rect 132542 352170 162834 352226
rect 162890 352170 162958 352226
rect 163014 352170 163082 352226
rect 163138 352170 163206 352226
rect 163262 352170 163878 352226
rect 163934 352170 164002 352226
rect 164058 352170 193554 352226
rect 193610 352170 193678 352226
rect 193734 352170 193802 352226
rect 193858 352170 193926 352226
rect 193982 352170 224274 352226
rect 224330 352170 224398 352226
rect 224454 352170 224522 352226
rect 224578 352170 224646 352226
rect 224702 352170 225878 352226
rect 225934 352170 226002 352226
rect 226058 352170 254994 352226
rect 255050 352170 255118 352226
rect 255174 352170 255242 352226
rect 255298 352170 255366 352226
rect 255422 352170 287878 352226
rect 287934 352170 288002 352226
rect 288058 352170 318598 352226
rect 318654 352170 318722 352226
rect 318778 352170 347154 352226
rect 347210 352170 347278 352226
rect 347334 352170 347402 352226
rect 347458 352170 347526 352226
rect 347582 352170 371878 352226
rect 371934 352170 372002 352226
rect 372058 352170 377874 352226
rect 377930 352170 377998 352226
rect 378054 352170 378122 352226
rect 378178 352170 378246 352226
rect 378302 352170 408594 352226
rect 408650 352170 408718 352226
rect 408774 352170 408842 352226
rect 408898 352170 408966 352226
rect 409022 352170 433878 352226
rect 433934 352170 434002 352226
rect 434058 352170 439314 352226
rect 439370 352170 439438 352226
rect 439494 352170 439562 352226
rect 439618 352170 439686 352226
rect 439742 352170 470034 352226
rect 470090 352170 470158 352226
rect 470214 352170 470282 352226
rect 470338 352170 470406 352226
rect 470462 352170 495878 352226
rect 495934 352170 496002 352226
rect 496058 352170 500754 352226
rect 500810 352170 500878 352226
rect 500934 352170 501002 352226
rect 501058 352170 501126 352226
rect 501182 352170 531474 352226
rect 531530 352170 531598 352226
rect 531654 352170 531722 352226
rect 531778 352170 531846 352226
rect 531902 352170 557878 352226
rect 557934 352170 558002 352226
rect 558058 352170 562194 352226
rect 562250 352170 562318 352226
rect 562374 352170 562442 352226
rect 562498 352170 562566 352226
rect 562622 352170 592914 352226
rect 592970 352170 593038 352226
rect 593094 352170 593162 352226
rect 593218 352170 593286 352226
rect 593342 352170 597456 352226
rect 597512 352170 597580 352226
rect 597636 352170 597704 352226
rect 597760 352170 597828 352226
rect 597884 352170 597980 352226
rect -1916 352102 597980 352170
rect -1916 352046 -1820 352102
rect -1764 352046 -1696 352102
rect -1640 352046 -1572 352102
rect -1516 352046 -1448 352102
rect -1392 352046 9234 352102
rect 9290 352046 9358 352102
rect 9414 352046 9482 352102
rect 9538 352046 9606 352102
rect 9662 352046 39878 352102
rect 39934 352046 40002 352102
rect 40058 352046 70674 352102
rect 70730 352046 70798 352102
rect 70854 352046 70922 352102
rect 70978 352046 71046 352102
rect 71102 352046 101878 352102
rect 101934 352046 102002 352102
rect 102058 352046 132114 352102
rect 132170 352046 132238 352102
rect 132294 352046 132362 352102
rect 132418 352046 132486 352102
rect 132542 352046 162834 352102
rect 162890 352046 162958 352102
rect 163014 352046 163082 352102
rect 163138 352046 163206 352102
rect 163262 352046 163878 352102
rect 163934 352046 164002 352102
rect 164058 352046 193554 352102
rect 193610 352046 193678 352102
rect 193734 352046 193802 352102
rect 193858 352046 193926 352102
rect 193982 352046 224274 352102
rect 224330 352046 224398 352102
rect 224454 352046 224522 352102
rect 224578 352046 224646 352102
rect 224702 352046 225878 352102
rect 225934 352046 226002 352102
rect 226058 352046 254994 352102
rect 255050 352046 255118 352102
rect 255174 352046 255242 352102
rect 255298 352046 255366 352102
rect 255422 352046 287878 352102
rect 287934 352046 288002 352102
rect 288058 352046 318598 352102
rect 318654 352046 318722 352102
rect 318778 352046 347154 352102
rect 347210 352046 347278 352102
rect 347334 352046 347402 352102
rect 347458 352046 347526 352102
rect 347582 352046 371878 352102
rect 371934 352046 372002 352102
rect 372058 352046 377874 352102
rect 377930 352046 377998 352102
rect 378054 352046 378122 352102
rect 378178 352046 378246 352102
rect 378302 352046 408594 352102
rect 408650 352046 408718 352102
rect 408774 352046 408842 352102
rect 408898 352046 408966 352102
rect 409022 352046 433878 352102
rect 433934 352046 434002 352102
rect 434058 352046 439314 352102
rect 439370 352046 439438 352102
rect 439494 352046 439562 352102
rect 439618 352046 439686 352102
rect 439742 352046 470034 352102
rect 470090 352046 470158 352102
rect 470214 352046 470282 352102
rect 470338 352046 470406 352102
rect 470462 352046 495878 352102
rect 495934 352046 496002 352102
rect 496058 352046 500754 352102
rect 500810 352046 500878 352102
rect 500934 352046 501002 352102
rect 501058 352046 501126 352102
rect 501182 352046 531474 352102
rect 531530 352046 531598 352102
rect 531654 352046 531722 352102
rect 531778 352046 531846 352102
rect 531902 352046 557878 352102
rect 557934 352046 558002 352102
rect 558058 352046 562194 352102
rect 562250 352046 562318 352102
rect 562374 352046 562442 352102
rect 562498 352046 562566 352102
rect 562622 352046 592914 352102
rect 592970 352046 593038 352102
rect 593094 352046 593162 352102
rect 593218 352046 593286 352102
rect 593342 352046 597456 352102
rect 597512 352046 597580 352102
rect 597636 352046 597704 352102
rect 597760 352046 597828 352102
rect 597884 352046 597980 352102
rect -1916 351978 597980 352046
rect -1916 351922 -1820 351978
rect -1764 351922 -1696 351978
rect -1640 351922 -1572 351978
rect -1516 351922 -1448 351978
rect -1392 351922 9234 351978
rect 9290 351922 9358 351978
rect 9414 351922 9482 351978
rect 9538 351922 9606 351978
rect 9662 351922 39878 351978
rect 39934 351922 40002 351978
rect 40058 351922 70674 351978
rect 70730 351922 70798 351978
rect 70854 351922 70922 351978
rect 70978 351922 71046 351978
rect 71102 351922 101878 351978
rect 101934 351922 102002 351978
rect 102058 351922 132114 351978
rect 132170 351922 132238 351978
rect 132294 351922 132362 351978
rect 132418 351922 132486 351978
rect 132542 351922 162834 351978
rect 162890 351922 162958 351978
rect 163014 351922 163082 351978
rect 163138 351922 163206 351978
rect 163262 351922 163878 351978
rect 163934 351922 164002 351978
rect 164058 351922 193554 351978
rect 193610 351922 193678 351978
rect 193734 351922 193802 351978
rect 193858 351922 193926 351978
rect 193982 351922 224274 351978
rect 224330 351922 224398 351978
rect 224454 351922 224522 351978
rect 224578 351922 224646 351978
rect 224702 351922 225878 351978
rect 225934 351922 226002 351978
rect 226058 351922 254994 351978
rect 255050 351922 255118 351978
rect 255174 351922 255242 351978
rect 255298 351922 255366 351978
rect 255422 351922 287878 351978
rect 287934 351922 288002 351978
rect 288058 351922 318598 351978
rect 318654 351922 318722 351978
rect 318778 351922 347154 351978
rect 347210 351922 347278 351978
rect 347334 351922 347402 351978
rect 347458 351922 347526 351978
rect 347582 351922 371878 351978
rect 371934 351922 372002 351978
rect 372058 351922 377874 351978
rect 377930 351922 377998 351978
rect 378054 351922 378122 351978
rect 378178 351922 378246 351978
rect 378302 351922 408594 351978
rect 408650 351922 408718 351978
rect 408774 351922 408842 351978
rect 408898 351922 408966 351978
rect 409022 351922 433878 351978
rect 433934 351922 434002 351978
rect 434058 351922 439314 351978
rect 439370 351922 439438 351978
rect 439494 351922 439562 351978
rect 439618 351922 439686 351978
rect 439742 351922 470034 351978
rect 470090 351922 470158 351978
rect 470214 351922 470282 351978
rect 470338 351922 470406 351978
rect 470462 351922 495878 351978
rect 495934 351922 496002 351978
rect 496058 351922 500754 351978
rect 500810 351922 500878 351978
rect 500934 351922 501002 351978
rect 501058 351922 501126 351978
rect 501182 351922 531474 351978
rect 531530 351922 531598 351978
rect 531654 351922 531722 351978
rect 531778 351922 531846 351978
rect 531902 351922 557878 351978
rect 557934 351922 558002 351978
rect 558058 351922 562194 351978
rect 562250 351922 562318 351978
rect 562374 351922 562442 351978
rect 562498 351922 562566 351978
rect 562622 351922 592914 351978
rect 592970 351922 593038 351978
rect 593094 351922 593162 351978
rect 593218 351922 593286 351978
rect 593342 351922 597456 351978
rect 597512 351922 597580 351978
rect 597636 351922 597704 351978
rect 597760 351922 597828 351978
rect 597884 351922 597980 351978
rect -1916 351826 597980 351922
rect 205980 349498 263860 349514
rect 205980 349442 205996 349498
rect 206052 349442 263788 349498
rect 263844 349442 263860 349498
rect 205980 349426 263860 349442
rect 334444 349498 523364 349514
rect 334444 349442 334460 349498
rect 334516 349442 523292 349498
rect 523348 349442 523364 349498
rect 334444 349426 523364 349442
rect 384676 349318 393444 349334
rect 384676 349262 393372 349318
rect 393428 349262 393444 349318
rect 384676 349246 393444 349262
rect 384676 348794 384764 349246
rect 350236 348778 384764 348794
rect 350236 348722 350252 348778
rect 350308 348722 384764 348778
rect 350236 348706 384764 348722
rect 203068 348598 263412 348614
rect 203068 348542 203084 348598
rect 203140 348542 263340 348598
rect 263396 348542 263412 348598
rect 203068 348526 263412 348542
rect 394812 348598 473300 348614
rect 394812 348542 394828 348598
rect 394884 348542 473228 348598
rect 473284 348542 473300 348598
rect 394812 348526 473300 348542
rect 197356 347878 263860 347894
rect 197356 347822 197372 347878
rect 197428 347822 263788 347878
rect 263844 347822 263860 347878
rect 197356 347806 263860 347822
rect -1916 346350 597980 346446
rect -1916 346294 -860 346350
rect -804 346294 -736 346350
rect -680 346294 -612 346350
rect -556 346294 -488 346350
rect -432 346294 5514 346350
rect 5570 346294 5638 346350
rect 5694 346294 5762 346350
rect 5818 346294 5886 346350
rect 5942 346294 24518 346350
rect 24574 346294 24642 346350
rect 24698 346294 36234 346350
rect 36290 346294 36358 346350
rect 36414 346294 36482 346350
rect 36538 346294 36606 346350
rect 36662 346294 55238 346350
rect 55294 346294 55362 346350
rect 55418 346294 66954 346350
rect 67010 346294 67078 346350
rect 67134 346294 67202 346350
rect 67258 346294 67326 346350
rect 67382 346294 86518 346350
rect 86574 346294 86642 346350
rect 86698 346294 97674 346350
rect 97730 346294 97798 346350
rect 97854 346294 97922 346350
rect 97978 346294 98046 346350
rect 98102 346294 117238 346350
rect 117294 346294 117362 346350
rect 117418 346294 128394 346350
rect 128450 346294 128518 346350
rect 128574 346294 128642 346350
rect 128698 346294 128766 346350
rect 128822 346294 148518 346350
rect 148574 346294 148642 346350
rect 148698 346294 159114 346350
rect 159170 346294 159238 346350
rect 159294 346294 159362 346350
rect 159418 346294 159486 346350
rect 159542 346294 179238 346350
rect 179294 346294 179362 346350
rect 179418 346294 189834 346350
rect 189890 346294 189958 346350
rect 190014 346294 190082 346350
rect 190138 346294 190206 346350
rect 190262 346294 210518 346350
rect 210574 346294 210642 346350
rect 210698 346294 220554 346350
rect 220610 346294 220678 346350
rect 220734 346294 220802 346350
rect 220858 346294 220926 346350
rect 220982 346294 241238 346350
rect 241294 346294 241362 346350
rect 241418 346294 251274 346350
rect 251330 346294 251398 346350
rect 251454 346294 251522 346350
rect 251578 346294 251646 346350
rect 251702 346294 272518 346350
rect 272574 346294 272642 346350
rect 272698 346294 303238 346350
rect 303294 346294 303362 346350
rect 303418 346294 343434 346350
rect 343490 346294 343558 346350
rect 343614 346294 343682 346350
rect 343738 346294 343806 346350
rect 343862 346294 356518 346350
rect 356574 346294 356642 346350
rect 356698 346294 374154 346350
rect 374210 346294 374278 346350
rect 374334 346294 374402 346350
rect 374458 346294 374526 346350
rect 374582 346294 387238 346350
rect 387294 346294 387362 346350
rect 387418 346294 404874 346350
rect 404930 346294 404998 346350
rect 405054 346294 405122 346350
rect 405178 346294 405246 346350
rect 405302 346294 418518 346350
rect 418574 346294 418642 346350
rect 418698 346294 435594 346350
rect 435650 346294 435718 346350
rect 435774 346294 435842 346350
rect 435898 346294 435966 346350
rect 436022 346294 449238 346350
rect 449294 346294 449362 346350
rect 449418 346294 466314 346350
rect 466370 346294 466438 346350
rect 466494 346294 466562 346350
rect 466618 346294 466686 346350
rect 466742 346294 480518 346350
rect 480574 346294 480642 346350
rect 480698 346294 497034 346350
rect 497090 346294 497158 346350
rect 497214 346294 497282 346350
rect 497338 346294 497406 346350
rect 497462 346294 511238 346350
rect 511294 346294 511362 346350
rect 511418 346294 527754 346350
rect 527810 346294 527878 346350
rect 527934 346294 528002 346350
rect 528058 346294 528126 346350
rect 528182 346294 542518 346350
rect 542574 346294 542642 346350
rect 542698 346294 558474 346350
rect 558530 346294 558598 346350
rect 558654 346294 558722 346350
rect 558778 346294 558846 346350
rect 558902 346294 573238 346350
rect 573294 346294 573362 346350
rect 573418 346294 589194 346350
rect 589250 346294 589318 346350
rect 589374 346294 589442 346350
rect 589498 346294 589566 346350
rect 589622 346294 596496 346350
rect 596552 346294 596620 346350
rect 596676 346294 596744 346350
rect 596800 346294 596868 346350
rect 596924 346294 597980 346350
rect -1916 346226 597980 346294
rect -1916 346170 -860 346226
rect -804 346170 -736 346226
rect -680 346170 -612 346226
rect -556 346170 -488 346226
rect -432 346170 5514 346226
rect 5570 346170 5638 346226
rect 5694 346170 5762 346226
rect 5818 346170 5886 346226
rect 5942 346170 24518 346226
rect 24574 346170 24642 346226
rect 24698 346170 36234 346226
rect 36290 346170 36358 346226
rect 36414 346170 36482 346226
rect 36538 346170 36606 346226
rect 36662 346170 55238 346226
rect 55294 346170 55362 346226
rect 55418 346170 66954 346226
rect 67010 346170 67078 346226
rect 67134 346170 67202 346226
rect 67258 346170 67326 346226
rect 67382 346170 86518 346226
rect 86574 346170 86642 346226
rect 86698 346170 97674 346226
rect 97730 346170 97798 346226
rect 97854 346170 97922 346226
rect 97978 346170 98046 346226
rect 98102 346170 117238 346226
rect 117294 346170 117362 346226
rect 117418 346170 128394 346226
rect 128450 346170 128518 346226
rect 128574 346170 128642 346226
rect 128698 346170 128766 346226
rect 128822 346170 148518 346226
rect 148574 346170 148642 346226
rect 148698 346170 159114 346226
rect 159170 346170 159238 346226
rect 159294 346170 159362 346226
rect 159418 346170 159486 346226
rect 159542 346170 179238 346226
rect 179294 346170 179362 346226
rect 179418 346170 189834 346226
rect 189890 346170 189958 346226
rect 190014 346170 190082 346226
rect 190138 346170 190206 346226
rect 190262 346170 210518 346226
rect 210574 346170 210642 346226
rect 210698 346170 220554 346226
rect 220610 346170 220678 346226
rect 220734 346170 220802 346226
rect 220858 346170 220926 346226
rect 220982 346170 241238 346226
rect 241294 346170 241362 346226
rect 241418 346170 251274 346226
rect 251330 346170 251398 346226
rect 251454 346170 251522 346226
rect 251578 346170 251646 346226
rect 251702 346170 272518 346226
rect 272574 346170 272642 346226
rect 272698 346170 303238 346226
rect 303294 346170 303362 346226
rect 303418 346170 343434 346226
rect 343490 346170 343558 346226
rect 343614 346170 343682 346226
rect 343738 346170 343806 346226
rect 343862 346170 356518 346226
rect 356574 346170 356642 346226
rect 356698 346170 374154 346226
rect 374210 346170 374278 346226
rect 374334 346170 374402 346226
rect 374458 346170 374526 346226
rect 374582 346170 387238 346226
rect 387294 346170 387362 346226
rect 387418 346170 404874 346226
rect 404930 346170 404998 346226
rect 405054 346170 405122 346226
rect 405178 346170 405246 346226
rect 405302 346170 418518 346226
rect 418574 346170 418642 346226
rect 418698 346170 435594 346226
rect 435650 346170 435718 346226
rect 435774 346170 435842 346226
rect 435898 346170 435966 346226
rect 436022 346170 449238 346226
rect 449294 346170 449362 346226
rect 449418 346170 466314 346226
rect 466370 346170 466438 346226
rect 466494 346170 466562 346226
rect 466618 346170 466686 346226
rect 466742 346170 480518 346226
rect 480574 346170 480642 346226
rect 480698 346170 497034 346226
rect 497090 346170 497158 346226
rect 497214 346170 497282 346226
rect 497338 346170 497406 346226
rect 497462 346170 511238 346226
rect 511294 346170 511362 346226
rect 511418 346170 527754 346226
rect 527810 346170 527878 346226
rect 527934 346170 528002 346226
rect 528058 346170 528126 346226
rect 528182 346170 542518 346226
rect 542574 346170 542642 346226
rect 542698 346170 558474 346226
rect 558530 346170 558598 346226
rect 558654 346170 558722 346226
rect 558778 346170 558846 346226
rect 558902 346170 573238 346226
rect 573294 346170 573362 346226
rect 573418 346170 589194 346226
rect 589250 346170 589318 346226
rect 589374 346170 589442 346226
rect 589498 346170 589566 346226
rect 589622 346170 596496 346226
rect 596552 346170 596620 346226
rect 596676 346170 596744 346226
rect 596800 346170 596868 346226
rect 596924 346170 597980 346226
rect -1916 346102 597980 346170
rect -1916 346046 -860 346102
rect -804 346046 -736 346102
rect -680 346046 -612 346102
rect -556 346046 -488 346102
rect -432 346046 5514 346102
rect 5570 346046 5638 346102
rect 5694 346046 5762 346102
rect 5818 346046 5886 346102
rect 5942 346046 24518 346102
rect 24574 346046 24642 346102
rect 24698 346046 36234 346102
rect 36290 346046 36358 346102
rect 36414 346046 36482 346102
rect 36538 346046 36606 346102
rect 36662 346046 55238 346102
rect 55294 346046 55362 346102
rect 55418 346046 66954 346102
rect 67010 346046 67078 346102
rect 67134 346046 67202 346102
rect 67258 346046 67326 346102
rect 67382 346046 86518 346102
rect 86574 346046 86642 346102
rect 86698 346046 97674 346102
rect 97730 346046 97798 346102
rect 97854 346046 97922 346102
rect 97978 346046 98046 346102
rect 98102 346046 117238 346102
rect 117294 346046 117362 346102
rect 117418 346046 128394 346102
rect 128450 346046 128518 346102
rect 128574 346046 128642 346102
rect 128698 346046 128766 346102
rect 128822 346046 148518 346102
rect 148574 346046 148642 346102
rect 148698 346046 159114 346102
rect 159170 346046 159238 346102
rect 159294 346046 159362 346102
rect 159418 346046 159486 346102
rect 159542 346046 179238 346102
rect 179294 346046 179362 346102
rect 179418 346046 189834 346102
rect 189890 346046 189958 346102
rect 190014 346046 190082 346102
rect 190138 346046 190206 346102
rect 190262 346046 210518 346102
rect 210574 346046 210642 346102
rect 210698 346046 220554 346102
rect 220610 346046 220678 346102
rect 220734 346046 220802 346102
rect 220858 346046 220926 346102
rect 220982 346046 241238 346102
rect 241294 346046 241362 346102
rect 241418 346046 251274 346102
rect 251330 346046 251398 346102
rect 251454 346046 251522 346102
rect 251578 346046 251646 346102
rect 251702 346046 272518 346102
rect 272574 346046 272642 346102
rect 272698 346046 303238 346102
rect 303294 346046 303362 346102
rect 303418 346046 343434 346102
rect 343490 346046 343558 346102
rect 343614 346046 343682 346102
rect 343738 346046 343806 346102
rect 343862 346046 356518 346102
rect 356574 346046 356642 346102
rect 356698 346046 374154 346102
rect 374210 346046 374278 346102
rect 374334 346046 374402 346102
rect 374458 346046 374526 346102
rect 374582 346046 387238 346102
rect 387294 346046 387362 346102
rect 387418 346046 404874 346102
rect 404930 346046 404998 346102
rect 405054 346046 405122 346102
rect 405178 346046 405246 346102
rect 405302 346046 418518 346102
rect 418574 346046 418642 346102
rect 418698 346046 435594 346102
rect 435650 346046 435718 346102
rect 435774 346046 435842 346102
rect 435898 346046 435966 346102
rect 436022 346046 449238 346102
rect 449294 346046 449362 346102
rect 449418 346046 466314 346102
rect 466370 346046 466438 346102
rect 466494 346046 466562 346102
rect 466618 346046 466686 346102
rect 466742 346046 480518 346102
rect 480574 346046 480642 346102
rect 480698 346046 497034 346102
rect 497090 346046 497158 346102
rect 497214 346046 497282 346102
rect 497338 346046 497406 346102
rect 497462 346046 511238 346102
rect 511294 346046 511362 346102
rect 511418 346046 527754 346102
rect 527810 346046 527878 346102
rect 527934 346046 528002 346102
rect 528058 346046 528126 346102
rect 528182 346046 542518 346102
rect 542574 346046 542642 346102
rect 542698 346046 558474 346102
rect 558530 346046 558598 346102
rect 558654 346046 558722 346102
rect 558778 346046 558846 346102
rect 558902 346046 573238 346102
rect 573294 346046 573362 346102
rect 573418 346046 589194 346102
rect 589250 346046 589318 346102
rect 589374 346046 589442 346102
rect 589498 346046 589566 346102
rect 589622 346046 596496 346102
rect 596552 346046 596620 346102
rect 596676 346046 596744 346102
rect 596800 346046 596868 346102
rect 596924 346046 597980 346102
rect -1916 345978 597980 346046
rect -1916 345922 -860 345978
rect -804 345922 -736 345978
rect -680 345922 -612 345978
rect -556 345922 -488 345978
rect -432 345922 5514 345978
rect 5570 345922 5638 345978
rect 5694 345922 5762 345978
rect 5818 345922 5886 345978
rect 5942 345922 24518 345978
rect 24574 345922 24642 345978
rect 24698 345922 36234 345978
rect 36290 345922 36358 345978
rect 36414 345922 36482 345978
rect 36538 345922 36606 345978
rect 36662 345922 55238 345978
rect 55294 345922 55362 345978
rect 55418 345922 66954 345978
rect 67010 345922 67078 345978
rect 67134 345922 67202 345978
rect 67258 345922 67326 345978
rect 67382 345922 86518 345978
rect 86574 345922 86642 345978
rect 86698 345922 97674 345978
rect 97730 345922 97798 345978
rect 97854 345922 97922 345978
rect 97978 345922 98046 345978
rect 98102 345922 117238 345978
rect 117294 345922 117362 345978
rect 117418 345922 128394 345978
rect 128450 345922 128518 345978
rect 128574 345922 128642 345978
rect 128698 345922 128766 345978
rect 128822 345922 148518 345978
rect 148574 345922 148642 345978
rect 148698 345922 159114 345978
rect 159170 345922 159238 345978
rect 159294 345922 159362 345978
rect 159418 345922 159486 345978
rect 159542 345922 179238 345978
rect 179294 345922 179362 345978
rect 179418 345922 189834 345978
rect 189890 345922 189958 345978
rect 190014 345922 190082 345978
rect 190138 345922 190206 345978
rect 190262 345922 210518 345978
rect 210574 345922 210642 345978
rect 210698 345922 220554 345978
rect 220610 345922 220678 345978
rect 220734 345922 220802 345978
rect 220858 345922 220926 345978
rect 220982 345922 241238 345978
rect 241294 345922 241362 345978
rect 241418 345922 251274 345978
rect 251330 345922 251398 345978
rect 251454 345922 251522 345978
rect 251578 345922 251646 345978
rect 251702 345922 272518 345978
rect 272574 345922 272642 345978
rect 272698 345922 303238 345978
rect 303294 345922 303362 345978
rect 303418 345922 343434 345978
rect 343490 345922 343558 345978
rect 343614 345922 343682 345978
rect 343738 345922 343806 345978
rect 343862 345922 356518 345978
rect 356574 345922 356642 345978
rect 356698 345922 374154 345978
rect 374210 345922 374278 345978
rect 374334 345922 374402 345978
rect 374458 345922 374526 345978
rect 374582 345922 387238 345978
rect 387294 345922 387362 345978
rect 387418 345922 404874 345978
rect 404930 345922 404998 345978
rect 405054 345922 405122 345978
rect 405178 345922 405246 345978
rect 405302 345922 418518 345978
rect 418574 345922 418642 345978
rect 418698 345922 435594 345978
rect 435650 345922 435718 345978
rect 435774 345922 435842 345978
rect 435898 345922 435966 345978
rect 436022 345922 449238 345978
rect 449294 345922 449362 345978
rect 449418 345922 466314 345978
rect 466370 345922 466438 345978
rect 466494 345922 466562 345978
rect 466618 345922 466686 345978
rect 466742 345922 480518 345978
rect 480574 345922 480642 345978
rect 480698 345922 497034 345978
rect 497090 345922 497158 345978
rect 497214 345922 497282 345978
rect 497338 345922 497406 345978
rect 497462 345922 511238 345978
rect 511294 345922 511362 345978
rect 511418 345922 527754 345978
rect 527810 345922 527878 345978
rect 527934 345922 528002 345978
rect 528058 345922 528126 345978
rect 528182 345922 542518 345978
rect 542574 345922 542642 345978
rect 542698 345922 558474 345978
rect 558530 345922 558598 345978
rect 558654 345922 558722 345978
rect 558778 345922 558846 345978
rect 558902 345922 573238 345978
rect 573294 345922 573362 345978
rect 573418 345922 589194 345978
rect 589250 345922 589318 345978
rect 589374 345922 589442 345978
rect 589498 345922 589566 345978
rect 589622 345922 596496 345978
rect 596552 345922 596620 345978
rect 596676 345922 596744 345978
rect 596800 345922 596868 345978
rect 596924 345922 597980 345978
rect -1916 345826 597980 345922
rect 195676 344638 263860 344654
rect 195676 344582 195692 344638
rect 195748 344582 263788 344638
rect 263844 344582 263860 344638
rect 195676 344566 263860 344582
rect 192428 344458 263972 344474
rect 192428 344402 192444 344458
rect 192500 344402 263900 344458
rect 263956 344402 263972 344458
rect 192428 344386 263972 344402
rect 334444 344458 460308 344474
rect 334444 344402 334460 344458
rect 334516 344402 460236 344458
rect 460292 344402 460308 344458
rect 334444 344386 460308 344402
rect 334444 344278 394900 344294
rect 334444 344222 334460 344278
rect 334516 344222 394828 344278
rect 394884 344222 394900 344278
rect 334444 344206 394900 344222
rect 189068 343558 262180 343574
rect 189068 343502 189084 343558
rect 189140 343502 262108 343558
rect 262164 343502 262180 343558
rect 189068 343486 262180 343502
rect 334332 343558 521124 343574
rect 334332 343502 334348 343558
rect 334404 343502 521052 343558
rect 521108 343502 521124 343558
rect 334332 343486 521124 343502
rect 195788 343018 263860 343034
rect 195788 342962 195804 343018
rect 195860 342962 263788 343018
rect 263844 342962 263860 343018
rect 195788 342946 263860 342962
rect 160508 342838 264756 342854
rect 160508 342782 160524 342838
rect 160580 342782 264684 342838
rect 264740 342782 264756 342838
rect 160508 342766 264756 342782
rect 20116 341938 126044 341954
rect 20116 341882 82684 341938
rect 82740 341882 126044 341938
rect 20116 341866 126044 341882
rect 20116 341774 20204 341866
rect 20060 341758 20204 341774
rect 20060 341702 20076 341758
rect 20132 341702 20204 341758
rect 20060 341686 20204 341702
rect 125956 341234 126044 341866
rect 478756 341938 534340 341954
rect 478756 341882 534268 341938
rect 534324 341882 534340 341938
rect 478756 341866 534340 341882
rect 478756 341774 478844 341866
rect 130044 341758 149564 341774
rect 130044 341702 130060 341758
rect 130116 341702 149564 341758
rect 130044 341686 149564 341702
rect 192316 341758 263860 341774
rect 192316 341702 192332 341758
rect 192388 341702 263788 341758
rect 263844 341702 263860 341758
rect 192316 341686 263860 341702
rect 476012 341758 478844 341774
rect 476012 341702 476028 341758
rect 476084 341702 478844 341758
rect 476012 341686 478844 341702
rect 144044 341578 144132 341594
rect 144044 341522 144060 341578
rect 144116 341522 144132 341578
rect 144044 341234 144132 341522
rect 149476 341414 149564 341686
rect 159724 341578 263972 341594
rect 159724 341522 159740 341578
rect 159796 341522 263900 341578
rect 263956 341522 263972 341578
rect 159724 341506 263972 341522
rect 334444 341578 407444 341594
rect 334444 341522 334460 341578
rect 334516 341522 407372 341578
rect 407428 341522 407444 341578
rect 334444 341506 407444 341522
rect 149476 341398 263860 341414
rect 149476 341342 263788 341398
rect 263844 341342 263860 341398
rect 149476 341326 263860 341342
rect 334332 341398 461204 341414
rect 334332 341342 334348 341398
rect 334404 341342 461132 341398
rect 461188 341342 461204 341398
rect 334332 341326 461204 341342
rect 125956 341218 141108 341234
rect 125956 341162 141036 341218
rect 141092 341162 141108 341218
rect 125956 341146 141108 341162
rect 144044 341218 201364 341234
rect 144044 341162 201292 341218
rect 201348 341162 201364 341218
rect 144044 341146 201364 341162
rect 352700 341218 473748 341234
rect 352700 341162 352716 341218
rect 352772 341162 414652 341218
rect 414708 341162 473676 341218
rect 473732 341162 473748 341218
rect 352700 341146 473748 341162
rect 122652 340498 263860 340514
rect 122652 340442 122668 340498
rect 122724 340442 263788 340498
rect 263844 340442 263860 340498
rect 122652 340426 263860 340442
rect 82444 340318 260388 340334
rect 82444 340262 82460 340318
rect 82516 340262 260316 340318
rect 260372 340262 260388 340318
rect 82444 340246 260388 340262
rect 460220 340138 521012 340154
rect 460220 340082 460236 340138
rect 460292 340082 520940 340138
rect 520996 340082 521012 340138
rect 460220 340066 521012 340082
rect 334444 339778 404532 339794
rect 334444 339722 334460 339778
rect 334516 339722 404460 339778
rect 404516 339722 404532 339778
rect 334444 339706 404532 339722
rect 455404 339778 455492 339794
rect 455404 339722 455420 339778
rect 455476 339722 455492 339778
rect 455404 339614 455492 339722
rect 351132 339598 455492 339614
rect 351132 339542 351148 339598
rect 351204 339542 455492 339598
rect 351132 339526 455492 339542
rect 334444 339418 455492 339434
rect 334444 339362 334460 339418
rect 334516 339362 455420 339418
rect 455476 339362 455492 339418
rect 334444 339346 455492 339362
rect 127580 339238 159812 339254
rect 127580 339182 127596 339238
rect 127652 339182 159740 339238
rect 159796 339182 159812 339238
rect 127580 339166 159812 339182
rect 384676 339238 393444 339254
rect 384676 339182 393372 339238
rect 393428 339182 393444 339238
rect 384676 339166 393444 339182
rect 461116 339238 502364 339254
rect 461116 339182 461132 339238
rect 461188 339182 502364 339238
rect 461116 339166 502364 339182
rect 384676 338714 384764 339166
rect 502276 338894 502364 339166
rect 338588 338698 384764 338714
rect 338588 338642 338604 338698
rect 338660 338642 384764 338698
rect 338588 338626 384764 338642
rect 455516 338878 455604 338894
rect 455516 338822 455532 338878
rect 455588 338822 455604 338878
rect 455516 338534 455604 338822
rect 502276 338878 517540 338894
rect 502276 338822 517468 338878
rect 517524 338822 517540 338878
rect 502276 338806 517540 338822
rect 82220 338518 122740 338534
rect 82220 338462 82236 338518
rect 82292 338462 122668 338518
rect 122724 338462 122740 338518
rect 82220 338446 122740 338462
rect 189404 338518 260164 338534
rect 189404 338462 189420 338518
rect 189476 338462 260092 338518
rect 260148 338462 260164 338518
rect 189404 338446 260164 338462
rect 394812 338518 455604 338534
rect 394812 338462 394828 338518
rect 394884 338462 455604 338518
rect 394812 338446 455604 338462
rect 334332 337978 396580 337994
rect 334332 337922 334348 337978
rect 334404 337922 396508 337978
rect 396564 337922 396580 337978
rect 334332 337906 396580 337922
rect 334444 337798 396580 337814
rect 334444 337742 334460 337798
rect 334516 337742 396580 337798
rect 334444 337726 396580 337742
rect 404556 337798 455380 337814
rect 404556 337742 404572 337798
rect 404628 337742 455308 337798
rect 455364 337742 455380 337798
rect 404556 337726 455380 337742
rect 396492 337634 396580 337726
rect 64188 337618 160596 337634
rect 64188 337562 64204 337618
rect 64260 337562 160524 337618
rect 160580 337562 160596 337618
rect 64188 337546 160596 337562
rect 334444 337618 394900 337634
rect 334444 337562 334460 337618
rect 334516 337562 394828 337618
rect 394884 337562 394900 337618
rect 334444 337546 394900 337562
rect 396492 337546 455324 337634
rect 455236 337094 455324 337546
rect 455236 337078 455380 337094
rect 455236 337022 455308 337078
rect 455364 337022 455380 337078
rect 455236 337006 455380 337022
rect 396492 336898 455716 336914
rect 396492 336842 396508 336898
rect 396564 336842 455716 336898
rect 396492 336826 455716 336842
rect 455628 336538 455716 336826
rect 455628 336482 455644 336538
rect 455700 336482 455716 336538
rect 455628 336466 455716 336482
rect 334444 336358 393220 336374
rect 334444 336302 334460 336358
rect 334516 336302 393148 336358
rect 393204 336302 393220 336358
rect 334444 336286 393220 336302
rect 20620 336178 124420 336194
rect 20620 336122 20636 336178
rect 20692 336122 124348 336178
rect 124404 336122 124420 336178
rect 20620 336106 124420 336122
rect 127580 336178 160484 336194
rect 127580 336122 127596 336178
rect 127652 336122 160412 336178
rect 160468 336122 160484 336178
rect 127580 336106 160484 336122
rect 334332 336178 399828 336194
rect 334332 336122 334348 336178
rect 334404 336122 399756 336178
rect 399812 336122 399828 336178
rect 334332 336106 399828 336122
rect 334444 335998 404644 336014
rect 334444 335942 334460 335998
rect 334516 335942 404572 335998
rect 404628 335942 404644 335998
rect 334444 335926 404644 335942
rect 404444 335098 455324 335114
rect 404444 335042 404460 335098
rect 404516 335042 455324 335098
rect 404444 335026 455324 335042
rect 455236 334754 455324 335026
rect 334444 334738 403300 334754
rect 334444 334682 334460 334738
rect 334516 334682 403228 334738
rect 403284 334682 403300 334738
rect 334444 334666 403300 334682
rect 455236 334738 455380 334754
rect 455236 334682 455308 334738
rect 455364 334682 455380 334738
rect 455236 334666 455380 334682
rect -1916 334350 597980 334446
rect -1916 334294 -1820 334350
rect -1764 334294 -1696 334350
rect -1640 334294 -1572 334350
rect -1516 334294 -1448 334350
rect -1392 334294 9234 334350
rect 9290 334294 9358 334350
rect 9414 334294 9482 334350
rect 9538 334294 9606 334350
rect 9662 334294 39878 334350
rect 39934 334294 40002 334350
rect 40058 334294 70674 334350
rect 70730 334294 70798 334350
rect 70854 334294 70922 334350
rect 70978 334294 71046 334350
rect 71102 334294 101878 334350
rect 101934 334294 102002 334350
rect 102058 334294 132114 334350
rect 132170 334294 132238 334350
rect 132294 334294 132362 334350
rect 132418 334294 132486 334350
rect 132542 334294 163878 334350
rect 163934 334294 164002 334350
rect 164058 334294 193554 334350
rect 193610 334294 193678 334350
rect 193734 334294 193802 334350
rect 193858 334294 193926 334350
rect 193982 334294 224274 334350
rect 224330 334294 224398 334350
rect 224454 334294 224522 334350
rect 224578 334294 224646 334350
rect 224702 334294 225878 334350
rect 225934 334294 226002 334350
rect 226058 334294 254994 334350
rect 255050 334294 255118 334350
rect 255174 334294 255242 334350
rect 255298 334294 255366 334350
rect 255422 334294 287878 334350
rect 287934 334294 288002 334350
rect 288058 334294 318598 334350
rect 318654 334294 318722 334350
rect 318778 334294 347154 334350
rect 347210 334294 347278 334350
rect 347334 334294 347402 334350
rect 347458 334294 347526 334350
rect 347582 334294 371878 334350
rect 371934 334294 372002 334350
rect 372058 334294 377874 334350
rect 377930 334294 377998 334350
rect 378054 334294 378122 334350
rect 378178 334294 378246 334350
rect 378302 334294 408594 334350
rect 408650 334294 408718 334350
rect 408774 334294 408842 334350
rect 408898 334294 408966 334350
rect 409022 334294 433878 334350
rect 433934 334294 434002 334350
rect 434058 334294 439314 334350
rect 439370 334294 439438 334350
rect 439494 334294 439562 334350
rect 439618 334294 439686 334350
rect 439742 334294 470034 334350
rect 470090 334294 470158 334350
rect 470214 334294 470282 334350
rect 470338 334294 470406 334350
rect 470462 334294 495878 334350
rect 495934 334294 496002 334350
rect 496058 334294 500754 334350
rect 500810 334294 500878 334350
rect 500934 334294 501002 334350
rect 501058 334294 501126 334350
rect 501182 334294 531474 334350
rect 531530 334294 531598 334350
rect 531654 334294 531722 334350
rect 531778 334294 531846 334350
rect 531902 334294 557878 334350
rect 557934 334294 558002 334350
rect 558058 334294 592914 334350
rect 592970 334294 593038 334350
rect 593094 334294 593162 334350
rect 593218 334294 593286 334350
rect 593342 334294 597456 334350
rect 597512 334294 597580 334350
rect 597636 334294 597704 334350
rect 597760 334294 597828 334350
rect 597884 334294 597980 334350
rect -1916 334226 597980 334294
rect -1916 334170 -1820 334226
rect -1764 334170 -1696 334226
rect -1640 334170 -1572 334226
rect -1516 334170 -1448 334226
rect -1392 334170 9234 334226
rect 9290 334170 9358 334226
rect 9414 334170 9482 334226
rect 9538 334170 9606 334226
rect 9662 334170 39878 334226
rect 39934 334170 40002 334226
rect 40058 334170 70674 334226
rect 70730 334170 70798 334226
rect 70854 334170 70922 334226
rect 70978 334170 71046 334226
rect 71102 334170 101878 334226
rect 101934 334170 102002 334226
rect 102058 334170 132114 334226
rect 132170 334170 132238 334226
rect 132294 334170 132362 334226
rect 132418 334170 132486 334226
rect 132542 334170 163878 334226
rect 163934 334170 164002 334226
rect 164058 334170 193554 334226
rect 193610 334170 193678 334226
rect 193734 334170 193802 334226
rect 193858 334170 193926 334226
rect 193982 334170 224274 334226
rect 224330 334170 224398 334226
rect 224454 334170 224522 334226
rect 224578 334170 224646 334226
rect 224702 334170 225878 334226
rect 225934 334170 226002 334226
rect 226058 334170 254994 334226
rect 255050 334170 255118 334226
rect 255174 334170 255242 334226
rect 255298 334170 255366 334226
rect 255422 334170 287878 334226
rect 287934 334170 288002 334226
rect 288058 334170 318598 334226
rect 318654 334170 318722 334226
rect 318778 334170 347154 334226
rect 347210 334170 347278 334226
rect 347334 334170 347402 334226
rect 347458 334170 347526 334226
rect 347582 334170 371878 334226
rect 371934 334170 372002 334226
rect 372058 334170 377874 334226
rect 377930 334170 377998 334226
rect 378054 334170 378122 334226
rect 378178 334170 378246 334226
rect 378302 334170 408594 334226
rect 408650 334170 408718 334226
rect 408774 334170 408842 334226
rect 408898 334170 408966 334226
rect 409022 334170 433878 334226
rect 433934 334170 434002 334226
rect 434058 334170 439314 334226
rect 439370 334170 439438 334226
rect 439494 334170 439562 334226
rect 439618 334170 439686 334226
rect 439742 334170 470034 334226
rect 470090 334170 470158 334226
rect 470214 334170 470282 334226
rect 470338 334170 470406 334226
rect 470462 334170 495878 334226
rect 495934 334170 496002 334226
rect 496058 334170 500754 334226
rect 500810 334170 500878 334226
rect 500934 334170 501002 334226
rect 501058 334170 501126 334226
rect 501182 334170 531474 334226
rect 531530 334170 531598 334226
rect 531654 334170 531722 334226
rect 531778 334170 531846 334226
rect 531902 334170 557878 334226
rect 557934 334170 558002 334226
rect 558058 334170 592914 334226
rect 592970 334170 593038 334226
rect 593094 334170 593162 334226
rect 593218 334170 593286 334226
rect 593342 334170 597456 334226
rect 597512 334170 597580 334226
rect 597636 334170 597704 334226
rect 597760 334170 597828 334226
rect 597884 334170 597980 334226
rect -1916 334102 597980 334170
rect -1916 334046 -1820 334102
rect -1764 334046 -1696 334102
rect -1640 334046 -1572 334102
rect -1516 334046 -1448 334102
rect -1392 334046 9234 334102
rect 9290 334046 9358 334102
rect 9414 334046 9482 334102
rect 9538 334046 9606 334102
rect 9662 334046 39878 334102
rect 39934 334046 40002 334102
rect 40058 334046 70674 334102
rect 70730 334046 70798 334102
rect 70854 334046 70922 334102
rect 70978 334046 71046 334102
rect 71102 334046 101878 334102
rect 101934 334046 102002 334102
rect 102058 334046 132114 334102
rect 132170 334046 132238 334102
rect 132294 334046 132362 334102
rect 132418 334046 132486 334102
rect 132542 334046 163878 334102
rect 163934 334046 164002 334102
rect 164058 334046 193554 334102
rect 193610 334046 193678 334102
rect 193734 334046 193802 334102
rect 193858 334046 193926 334102
rect 193982 334046 224274 334102
rect 224330 334046 224398 334102
rect 224454 334046 224522 334102
rect 224578 334046 224646 334102
rect 224702 334046 225878 334102
rect 225934 334046 226002 334102
rect 226058 334046 254994 334102
rect 255050 334046 255118 334102
rect 255174 334046 255242 334102
rect 255298 334046 255366 334102
rect 255422 334046 287878 334102
rect 287934 334046 288002 334102
rect 288058 334046 318598 334102
rect 318654 334046 318722 334102
rect 318778 334046 347154 334102
rect 347210 334046 347278 334102
rect 347334 334046 347402 334102
rect 347458 334046 347526 334102
rect 347582 334046 371878 334102
rect 371934 334046 372002 334102
rect 372058 334046 377874 334102
rect 377930 334046 377998 334102
rect 378054 334046 378122 334102
rect 378178 334046 378246 334102
rect 378302 334046 408594 334102
rect 408650 334046 408718 334102
rect 408774 334046 408842 334102
rect 408898 334046 408966 334102
rect 409022 334046 433878 334102
rect 433934 334046 434002 334102
rect 434058 334046 439314 334102
rect 439370 334046 439438 334102
rect 439494 334046 439562 334102
rect 439618 334046 439686 334102
rect 439742 334046 470034 334102
rect 470090 334046 470158 334102
rect 470214 334046 470282 334102
rect 470338 334046 470406 334102
rect 470462 334046 495878 334102
rect 495934 334046 496002 334102
rect 496058 334046 500754 334102
rect 500810 334046 500878 334102
rect 500934 334046 501002 334102
rect 501058 334046 501126 334102
rect 501182 334046 531474 334102
rect 531530 334046 531598 334102
rect 531654 334046 531722 334102
rect 531778 334046 531846 334102
rect 531902 334046 557878 334102
rect 557934 334046 558002 334102
rect 558058 334046 592914 334102
rect 592970 334046 593038 334102
rect 593094 334046 593162 334102
rect 593218 334046 593286 334102
rect 593342 334046 597456 334102
rect 597512 334046 597580 334102
rect 597636 334046 597704 334102
rect 597760 334046 597828 334102
rect 597884 334046 597980 334102
rect -1916 333978 597980 334046
rect -1916 333922 -1820 333978
rect -1764 333922 -1696 333978
rect -1640 333922 -1572 333978
rect -1516 333922 -1448 333978
rect -1392 333922 9234 333978
rect 9290 333922 9358 333978
rect 9414 333922 9482 333978
rect 9538 333922 9606 333978
rect 9662 333922 39878 333978
rect 39934 333922 40002 333978
rect 40058 333922 70674 333978
rect 70730 333922 70798 333978
rect 70854 333922 70922 333978
rect 70978 333922 71046 333978
rect 71102 333922 101878 333978
rect 101934 333922 102002 333978
rect 102058 333922 132114 333978
rect 132170 333922 132238 333978
rect 132294 333922 132362 333978
rect 132418 333922 132486 333978
rect 132542 333922 163878 333978
rect 163934 333922 164002 333978
rect 164058 333922 193554 333978
rect 193610 333922 193678 333978
rect 193734 333922 193802 333978
rect 193858 333922 193926 333978
rect 193982 333922 224274 333978
rect 224330 333922 224398 333978
rect 224454 333922 224522 333978
rect 224578 333922 224646 333978
rect 224702 333922 225878 333978
rect 225934 333922 226002 333978
rect 226058 333922 254994 333978
rect 255050 333922 255118 333978
rect 255174 333922 255242 333978
rect 255298 333922 255366 333978
rect 255422 333922 287878 333978
rect 287934 333922 288002 333978
rect 288058 333922 318598 333978
rect 318654 333922 318722 333978
rect 318778 333922 347154 333978
rect 347210 333922 347278 333978
rect 347334 333922 347402 333978
rect 347458 333922 347526 333978
rect 347582 333922 371878 333978
rect 371934 333922 372002 333978
rect 372058 333922 377874 333978
rect 377930 333922 377998 333978
rect 378054 333922 378122 333978
rect 378178 333922 378246 333978
rect 378302 333922 408594 333978
rect 408650 333922 408718 333978
rect 408774 333922 408842 333978
rect 408898 333922 408966 333978
rect 409022 333922 433878 333978
rect 433934 333922 434002 333978
rect 434058 333922 439314 333978
rect 439370 333922 439438 333978
rect 439494 333922 439562 333978
rect 439618 333922 439686 333978
rect 439742 333922 470034 333978
rect 470090 333922 470158 333978
rect 470214 333922 470282 333978
rect 470338 333922 470406 333978
rect 470462 333922 495878 333978
rect 495934 333922 496002 333978
rect 496058 333922 500754 333978
rect 500810 333922 500878 333978
rect 500934 333922 501002 333978
rect 501058 333922 501126 333978
rect 501182 333922 531474 333978
rect 531530 333922 531598 333978
rect 531654 333922 531722 333978
rect 531778 333922 531846 333978
rect 531902 333922 557878 333978
rect 557934 333922 558002 333978
rect 558058 333922 592914 333978
rect 592970 333922 593038 333978
rect 593094 333922 593162 333978
rect 593218 333922 593286 333978
rect 593342 333922 597456 333978
rect 597512 333922 597580 333978
rect 597636 333922 597704 333978
rect 597760 333922 597828 333978
rect 597884 333922 597980 333978
rect -1916 333826 597980 333922
rect 334444 333658 393556 333674
rect 334444 333602 334460 333658
rect 334516 333602 393484 333658
rect 393540 333602 393556 333658
rect 334444 333586 393556 333602
rect 127580 332758 160596 332774
rect 127580 332702 127596 332758
rect 127652 332702 160524 332758
rect 160580 332702 160596 332758
rect 127580 332686 160596 332702
rect 393132 332686 393668 332774
rect 393132 332594 393220 332686
rect 393580 332594 393668 332686
rect 334444 332578 393220 332594
rect 334444 332522 334460 332578
rect 334516 332522 393220 332578
rect 334444 332506 393220 332522
rect 393356 332578 393444 332594
rect 393356 332522 393372 332578
rect 393428 332522 393444 332578
rect 393356 332054 393444 332522
rect 393580 332578 394900 332594
rect 393580 332522 394828 332578
rect 394884 332522 394900 332578
rect 393580 332506 394900 332522
rect 344412 332038 393444 332054
rect 344412 331982 344428 332038
rect 344484 331982 393444 332038
rect 344412 331966 393444 331982
rect 18044 331858 162612 331874
rect 18044 331802 18060 331858
rect 18116 331802 162540 331858
rect 162596 331802 162612 331858
rect 18044 331786 162612 331802
rect 393132 331858 455604 331874
rect 393132 331802 393148 331858
rect 393204 331802 455532 331858
rect 455588 331802 455604 331858
rect 393132 331786 455604 331802
rect 572836 331678 579700 331694
rect 572836 331622 579628 331678
rect 579684 331622 579700 331678
rect 572836 331606 579700 331622
rect 64188 331498 263860 331514
rect 64188 331442 64204 331498
rect 64260 331442 263788 331498
rect 263844 331442 263860 331498
rect 64188 331426 263860 331442
rect 572836 331154 572924 331606
rect 166220 331138 263972 331154
rect 166220 331082 166236 331138
rect 166292 331082 263900 331138
rect 263956 331082 263972 331138
rect 166220 331066 263972 331082
rect 464476 331138 572924 331154
rect 464476 331082 464492 331138
rect 464548 331082 572924 331138
rect 464476 331066 572924 331082
rect 65196 330958 263860 330974
rect 65196 330902 65212 330958
rect 65268 330902 263788 330958
rect 263844 330902 263860 330958
rect 65196 330886 263860 330902
rect 337692 330958 455380 330974
rect 337692 330902 337708 330958
rect 337764 330902 455308 330958
rect 455364 330902 455380 330958
rect 337692 330886 455380 330902
rect 127580 330778 264084 330794
rect 127580 330722 127596 330778
rect 127652 330722 264012 330778
rect 264068 330722 264084 330778
rect 127580 330706 264084 330722
rect 334444 330778 395012 330794
rect 334444 330722 334460 330778
rect 334516 330722 394940 330778
rect 394996 330722 395012 330778
rect 334444 330706 395012 330722
rect 162524 330598 263860 330614
rect 162524 330542 162540 330598
rect 162596 330542 263788 330598
rect 263844 330542 263860 330598
rect 162524 330526 263860 330542
rect 64188 330418 166308 330434
rect 64188 330362 64204 330418
rect 64260 330362 166236 330418
rect 166292 330362 166308 330418
rect 64188 330346 166308 330362
rect 403212 330058 455492 330074
rect 403212 330002 403228 330058
rect 403284 330002 455492 330058
rect 403212 329986 455492 330002
rect 462796 330058 534340 330074
rect 462796 330002 462812 330058
rect 462868 330002 534268 330058
rect 534324 330002 534340 330058
rect 462796 329986 534340 330002
rect 455404 329878 455492 329986
rect 455404 329822 455420 329878
rect 455476 329822 455492 329878
rect 455404 329806 455492 329822
rect 384676 329518 393332 329534
rect 384676 329462 393260 329518
rect 393316 329462 393332 329518
rect 384676 329446 393332 329462
rect 384676 329354 384764 329446
rect 334444 329338 384764 329354
rect 334444 329282 334460 329338
rect 334516 329282 384764 329338
rect 334444 329266 384764 329282
rect -1916 328350 597980 328446
rect -1916 328294 -860 328350
rect -804 328294 -736 328350
rect -680 328294 -612 328350
rect -556 328294 -488 328350
rect -432 328294 5514 328350
rect 5570 328294 5638 328350
rect 5694 328294 5762 328350
rect 5818 328294 5886 328350
rect 5942 328294 24518 328350
rect 24574 328294 24642 328350
rect 24698 328294 36234 328350
rect 36290 328294 36358 328350
rect 36414 328294 36482 328350
rect 36538 328294 36606 328350
rect 36662 328294 55238 328350
rect 55294 328294 55362 328350
rect 55418 328294 66954 328350
rect 67010 328294 67078 328350
rect 67134 328294 67202 328350
rect 67258 328294 67326 328350
rect 67382 328294 86518 328350
rect 86574 328294 86642 328350
rect 86698 328294 97674 328350
rect 97730 328294 97798 328350
rect 97854 328294 97922 328350
rect 97978 328294 98046 328350
rect 98102 328294 117238 328350
rect 117294 328294 117362 328350
rect 117418 328294 128394 328350
rect 128450 328294 128518 328350
rect 128574 328294 128642 328350
rect 128698 328294 128766 328350
rect 128822 328294 148518 328350
rect 148574 328294 148642 328350
rect 148698 328294 159114 328350
rect 159170 328294 159238 328350
rect 159294 328294 159362 328350
rect 159418 328294 159486 328350
rect 159542 328294 179238 328350
rect 179294 328294 179362 328350
rect 179418 328294 189834 328350
rect 189890 328294 189958 328350
rect 190014 328294 190082 328350
rect 190138 328294 190206 328350
rect 190262 328294 210518 328350
rect 210574 328294 210642 328350
rect 210698 328294 220554 328350
rect 220610 328294 220678 328350
rect 220734 328294 220802 328350
rect 220858 328294 220926 328350
rect 220982 328294 241238 328350
rect 241294 328294 241362 328350
rect 241418 328294 251274 328350
rect 251330 328294 251398 328350
rect 251454 328294 251522 328350
rect 251578 328294 251646 328350
rect 251702 328294 272518 328350
rect 272574 328294 272642 328350
rect 272698 328294 303238 328350
rect 303294 328294 303362 328350
rect 303418 328294 343434 328350
rect 343490 328294 343558 328350
rect 343614 328294 343682 328350
rect 343738 328294 343806 328350
rect 343862 328294 356518 328350
rect 356574 328294 356642 328350
rect 356698 328294 374154 328350
rect 374210 328294 374278 328350
rect 374334 328294 374402 328350
rect 374458 328294 374526 328350
rect 374582 328294 387238 328350
rect 387294 328294 387362 328350
rect 387418 328294 404874 328350
rect 404930 328294 404998 328350
rect 405054 328294 405122 328350
rect 405178 328294 405246 328350
rect 405302 328294 418518 328350
rect 418574 328294 418642 328350
rect 418698 328294 435594 328350
rect 435650 328294 435718 328350
rect 435774 328294 435842 328350
rect 435898 328294 435966 328350
rect 436022 328294 449238 328350
rect 449294 328294 449362 328350
rect 449418 328294 466314 328350
rect 466370 328294 466438 328350
rect 466494 328294 466562 328350
rect 466618 328294 466686 328350
rect 466742 328294 480518 328350
rect 480574 328294 480642 328350
rect 480698 328294 497034 328350
rect 497090 328294 497158 328350
rect 497214 328294 497282 328350
rect 497338 328294 497406 328350
rect 497462 328294 511238 328350
rect 511294 328294 511362 328350
rect 511418 328294 527754 328350
rect 527810 328294 527878 328350
rect 527934 328294 528002 328350
rect 528058 328294 528126 328350
rect 528182 328294 542518 328350
rect 542574 328294 542642 328350
rect 542698 328294 558474 328350
rect 558530 328294 558598 328350
rect 558654 328294 558722 328350
rect 558778 328294 558846 328350
rect 558902 328294 573238 328350
rect 573294 328294 573362 328350
rect 573418 328294 589194 328350
rect 589250 328294 589318 328350
rect 589374 328294 589442 328350
rect 589498 328294 589566 328350
rect 589622 328294 596496 328350
rect 596552 328294 596620 328350
rect 596676 328294 596744 328350
rect 596800 328294 596868 328350
rect 596924 328294 597980 328350
rect -1916 328226 597980 328294
rect -1916 328170 -860 328226
rect -804 328170 -736 328226
rect -680 328170 -612 328226
rect -556 328170 -488 328226
rect -432 328170 5514 328226
rect 5570 328170 5638 328226
rect 5694 328170 5762 328226
rect 5818 328170 5886 328226
rect 5942 328170 24518 328226
rect 24574 328170 24642 328226
rect 24698 328170 36234 328226
rect 36290 328170 36358 328226
rect 36414 328170 36482 328226
rect 36538 328170 36606 328226
rect 36662 328170 55238 328226
rect 55294 328170 55362 328226
rect 55418 328170 66954 328226
rect 67010 328170 67078 328226
rect 67134 328170 67202 328226
rect 67258 328170 67326 328226
rect 67382 328170 86518 328226
rect 86574 328170 86642 328226
rect 86698 328170 97674 328226
rect 97730 328170 97798 328226
rect 97854 328170 97922 328226
rect 97978 328170 98046 328226
rect 98102 328170 117238 328226
rect 117294 328170 117362 328226
rect 117418 328170 128394 328226
rect 128450 328170 128518 328226
rect 128574 328170 128642 328226
rect 128698 328170 128766 328226
rect 128822 328170 148518 328226
rect 148574 328170 148642 328226
rect 148698 328170 159114 328226
rect 159170 328170 159238 328226
rect 159294 328170 159362 328226
rect 159418 328170 159486 328226
rect 159542 328170 179238 328226
rect 179294 328170 179362 328226
rect 179418 328170 189834 328226
rect 189890 328170 189958 328226
rect 190014 328170 190082 328226
rect 190138 328170 190206 328226
rect 190262 328170 210518 328226
rect 210574 328170 210642 328226
rect 210698 328170 220554 328226
rect 220610 328170 220678 328226
rect 220734 328170 220802 328226
rect 220858 328170 220926 328226
rect 220982 328170 241238 328226
rect 241294 328170 241362 328226
rect 241418 328170 251274 328226
rect 251330 328170 251398 328226
rect 251454 328170 251522 328226
rect 251578 328170 251646 328226
rect 251702 328170 272518 328226
rect 272574 328170 272642 328226
rect 272698 328170 303238 328226
rect 303294 328170 303362 328226
rect 303418 328170 343434 328226
rect 343490 328170 343558 328226
rect 343614 328170 343682 328226
rect 343738 328170 343806 328226
rect 343862 328170 356518 328226
rect 356574 328170 356642 328226
rect 356698 328170 374154 328226
rect 374210 328170 374278 328226
rect 374334 328170 374402 328226
rect 374458 328170 374526 328226
rect 374582 328170 387238 328226
rect 387294 328170 387362 328226
rect 387418 328170 404874 328226
rect 404930 328170 404998 328226
rect 405054 328170 405122 328226
rect 405178 328170 405246 328226
rect 405302 328170 418518 328226
rect 418574 328170 418642 328226
rect 418698 328170 435594 328226
rect 435650 328170 435718 328226
rect 435774 328170 435842 328226
rect 435898 328170 435966 328226
rect 436022 328170 449238 328226
rect 449294 328170 449362 328226
rect 449418 328170 466314 328226
rect 466370 328170 466438 328226
rect 466494 328170 466562 328226
rect 466618 328170 466686 328226
rect 466742 328170 480518 328226
rect 480574 328170 480642 328226
rect 480698 328170 497034 328226
rect 497090 328170 497158 328226
rect 497214 328170 497282 328226
rect 497338 328170 497406 328226
rect 497462 328170 511238 328226
rect 511294 328170 511362 328226
rect 511418 328170 527754 328226
rect 527810 328170 527878 328226
rect 527934 328170 528002 328226
rect 528058 328170 528126 328226
rect 528182 328170 542518 328226
rect 542574 328170 542642 328226
rect 542698 328170 558474 328226
rect 558530 328170 558598 328226
rect 558654 328170 558722 328226
rect 558778 328170 558846 328226
rect 558902 328170 573238 328226
rect 573294 328170 573362 328226
rect 573418 328170 589194 328226
rect 589250 328170 589318 328226
rect 589374 328170 589442 328226
rect 589498 328170 589566 328226
rect 589622 328170 596496 328226
rect 596552 328170 596620 328226
rect 596676 328170 596744 328226
rect 596800 328170 596868 328226
rect 596924 328170 597980 328226
rect -1916 328102 597980 328170
rect -1916 328046 -860 328102
rect -804 328046 -736 328102
rect -680 328046 -612 328102
rect -556 328046 -488 328102
rect -432 328046 5514 328102
rect 5570 328046 5638 328102
rect 5694 328046 5762 328102
rect 5818 328046 5886 328102
rect 5942 328046 24518 328102
rect 24574 328046 24642 328102
rect 24698 328046 36234 328102
rect 36290 328046 36358 328102
rect 36414 328046 36482 328102
rect 36538 328046 36606 328102
rect 36662 328046 55238 328102
rect 55294 328046 55362 328102
rect 55418 328046 66954 328102
rect 67010 328046 67078 328102
rect 67134 328046 67202 328102
rect 67258 328046 67326 328102
rect 67382 328046 86518 328102
rect 86574 328046 86642 328102
rect 86698 328046 97674 328102
rect 97730 328046 97798 328102
rect 97854 328046 97922 328102
rect 97978 328046 98046 328102
rect 98102 328046 117238 328102
rect 117294 328046 117362 328102
rect 117418 328046 128394 328102
rect 128450 328046 128518 328102
rect 128574 328046 128642 328102
rect 128698 328046 128766 328102
rect 128822 328046 148518 328102
rect 148574 328046 148642 328102
rect 148698 328046 159114 328102
rect 159170 328046 159238 328102
rect 159294 328046 159362 328102
rect 159418 328046 159486 328102
rect 159542 328046 179238 328102
rect 179294 328046 179362 328102
rect 179418 328046 189834 328102
rect 189890 328046 189958 328102
rect 190014 328046 190082 328102
rect 190138 328046 190206 328102
rect 190262 328046 210518 328102
rect 210574 328046 210642 328102
rect 210698 328046 220554 328102
rect 220610 328046 220678 328102
rect 220734 328046 220802 328102
rect 220858 328046 220926 328102
rect 220982 328046 241238 328102
rect 241294 328046 241362 328102
rect 241418 328046 251274 328102
rect 251330 328046 251398 328102
rect 251454 328046 251522 328102
rect 251578 328046 251646 328102
rect 251702 328046 272518 328102
rect 272574 328046 272642 328102
rect 272698 328046 303238 328102
rect 303294 328046 303362 328102
rect 303418 328046 343434 328102
rect 343490 328046 343558 328102
rect 343614 328046 343682 328102
rect 343738 328046 343806 328102
rect 343862 328046 356518 328102
rect 356574 328046 356642 328102
rect 356698 328046 374154 328102
rect 374210 328046 374278 328102
rect 374334 328046 374402 328102
rect 374458 328046 374526 328102
rect 374582 328046 387238 328102
rect 387294 328046 387362 328102
rect 387418 328046 404874 328102
rect 404930 328046 404998 328102
rect 405054 328046 405122 328102
rect 405178 328046 405246 328102
rect 405302 328046 418518 328102
rect 418574 328046 418642 328102
rect 418698 328046 435594 328102
rect 435650 328046 435718 328102
rect 435774 328046 435842 328102
rect 435898 328046 435966 328102
rect 436022 328046 449238 328102
rect 449294 328046 449362 328102
rect 449418 328046 466314 328102
rect 466370 328046 466438 328102
rect 466494 328046 466562 328102
rect 466618 328046 466686 328102
rect 466742 328046 480518 328102
rect 480574 328046 480642 328102
rect 480698 328046 497034 328102
rect 497090 328046 497158 328102
rect 497214 328046 497282 328102
rect 497338 328046 497406 328102
rect 497462 328046 511238 328102
rect 511294 328046 511362 328102
rect 511418 328046 527754 328102
rect 527810 328046 527878 328102
rect 527934 328046 528002 328102
rect 528058 328046 528126 328102
rect 528182 328046 542518 328102
rect 542574 328046 542642 328102
rect 542698 328046 558474 328102
rect 558530 328046 558598 328102
rect 558654 328046 558722 328102
rect 558778 328046 558846 328102
rect 558902 328046 573238 328102
rect 573294 328046 573362 328102
rect 573418 328046 589194 328102
rect 589250 328046 589318 328102
rect 589374 328046 589442 328102
rect 589498 328046 589566 328102
rect 589622 328046 596496 328102
rect 596552 328046 596620 328102
rect 596676 328046 596744 328102
rect 596800 328046 596868 328102
rect 596924 328046 597980 328102
rect -1916 327978 597980 328046
rect -1916 327922 -860 327978
rect -804 327922 -736 327978
rect -680 327922 -612 327978
rect -556 327922 -488 327978
rect -432 327922 5514 327978
rect 5570 327922 5638 327978
rect 5694 327922 5762 327978
rect 5818 327922 5886 327978
rect 5942 327922 24518 327978
rect 24574 327922 24642 327978
rect 24698 327922 36234 327978
rect 36290 327922 36358 327978
rect 36414 327922 36482 327978
rect 36538 327922 36606 327978
rect 36662 327922 55238 327978
rect 55294 327922 55362 327978
rect 55418 327922 66954 327978
rect 67010 327922 67078 327978
rect 67134 327922 67202 327978
rect 67258 327922 67326 327978
rect 67382 327922 86518 327978
rect 86574 327922 86642 327978
rect 86698 327922 97674 327978
rect 97730 327922 97798 327978
rect 97854 327922 97922 327978
rect 97978 327922 98046 327978
rect 98102 327922 117238 327978
rect 117294 327922 117362 327978
rect 117418 327922 128394 327978
rect 128450 327922 128518 327978
rect 128574 327922 128642 327978
rect 128698 327922 128766 327978
rect 128822 327922 148518 327978
rect 148574 327922 148642 327978
rect 148698 327922 159114 327978
rect 159170 327922 159238 327978
rect 159294 327922 159362 327978
rect 159418 327922 159486 327978
rect 159542 327922 179238 327978
rect 179294 327922 179362 327978
rect 179418 327922 189834 327978
rect 189890 327922 189958 327978
rect 190014 327922 190082 327978
rect 190138 327922 190206 327978
rect 190262 327922 210518 327978
rect 210574 327922 210642 327978
rect 210698 327922 220554 327978
rect 220610 327922 220678 327978
rect 220734 327922 220802 327978
rect 220858 327922 220926 327978
rect 220982 327922 241238 327978
rect 241294 327922 241362 327978
rect 241418 327922 251274 327978
rect 251330 327922 251398 327978
rect 251454 327922 251522 327978
rect 251578 327922 251646 327978
rect 251702 327922 272518 327978
rect 272574 327922 272642 327978
rect 272698 327922 303238 327978
rect 303294 327922 303362 327978
rect 303418 327922 343434 327978
rect 343490 327922 343558 327978
rect 343614 327922 343682 327978
rect 343738 327922 343806 327978
rect 343862 327922 356518 327978
rect 356574 327922 356642 327978
rect 356698 327922 374154 327978
rect 374210 327922 374278 327978
rect 374334 327922 374402 327978
rect 374458 327922 374526 327978
rect 374582 327922 387238 327978
rect 387294 327922 387362 327978
rect 387418 327922 404874 327978
rect 404930 327922 404998 327978
rect 405054 327922 405122 327978
rect 405178 327922 405246 327978
rect 405302 327922 418518 327978
rect 418574 327922 418642 327978
rect 418698 327922 435594 327978
rect 435650 327922 435718 327978
rect 435774 327922 435842 327978
rect 435898 327922 435966 327978
rect 436022 327922 449238 327978
rect 449294 327922 449362 327978
rect 449418 327922 466314 327978
rect 466370 327922 466438 327978
rect 466494 327922 466562 327978
rect 466618 327922 466686 327978
rect 466742 327922 480518 327978
rect 480574 327922 480642 327978
rect 480698 327922 497034 327978
rect 497090 327922 497158 327978
rect 497214 327922 497282 327978
rect 497338 327922 497406 327978
rect 497462 327922 511238 327978
rect 511294 327922 511362 327978
rect 511418 327922 527754 327978
rect 527810 327922 527878 327978
rect 527934 327922 528002 327978
rect 528058 327922 528126 327978
rect 528182 327922 542518 327978
rect 542574 327922 542642 327978
rect 542698 327922 558474 327978
rect 558530 327922 558598 327978
rect 558654 327922 558722 327978
rect 558778 327922 558846 327978
rect 558902 327922 573238 327978
rect 573294 327922 573362 327978
rect 573418 327922 589194 327978
rect 589250 327922 589318 327978
rect 589374 327922 589442 327978
rect 589498 327922 589566 327978
rect 589622 327922 596496 327978
rect 596552 327922 596620 327978
rect 596676 327922 596744 327978
rect 596800 327922 596868 327978
rect 596924 327922 597980 327978
rect -1916 327826 597980 327922
rect 20060 327538 263860 327554
rect 20060 327482 20076 327538
rect 20132 327482 263788 327538
rect 263844 327482 263860 327538
rect 20060 327466 263860 327482
rect 334444 327538 394900 327554
rect 334444 327482 334460 327538
rect 334516 327482 394828 327538
rect 394884 327482 394900 327538
rect 334444 327466 394900 327482
rect 124332 327358 263972 327374
rect 124332 327302 124348 327358
rect 124404 327302 263900 327358
rect 263956 327302 263972 327358
rect 124332 327286 263972 327302
rect 334444 327358 394116 327374
rect 334444 327302 334460 327358
rect 334516 327302 394044 327358
rect 394100 327302 394116 327358
rect 334444 327286 394116 327302
rect 404556 326818 583060 326834
rect 404556 326762 404572 326818
rect 404628 326762 582988 326818
rect 583044 326762 583060 326818
rect 404556 326746 583060 326762
rect 160396 325918 264980 325934
rect 160396 325862 160412 325918
rect 160468 325862 264908 325918
rect 264964 325862 264980 325918
rect 160396 325846 264980 325862
rect 334444 325918 462884 325934
rect 334444 325862 334460 325918
rect 334516 325862 462812 325918
rect 462868 325862 462884 325918
rect 334444 325846 462884 325862
rect 160508 325738 264644 325754
rect 160508 325682 160524 325738
rect 160580 325682 264572 325738
rect 264628 325682 264644 325738
rect 160508 325666 264644 325682
rect 206092 325558 263860 325574
rect 206092 325502 206108 325558
rect 206164 325502 263788 325558
rect 263844 325502 263860 325558
rect 206092 325486 263860 325502
rect 460220 325018 535124 325034
rect 460220 324962 460236 325018
rect 460292 324962 535052 325018
rect 535108 324962 535124 325018
rect 460220 324946 535124 324962
rect 204860 324118 263860 324134
rect 204860 324062 204876 324118
rect 204932 324062 263788 324118
rect 263844 324062 263860 324118
rect 204860 324046 263860 324062
rect 334444 324118 523364 324134
rect 334444 324062 334460 324118
rect 334516 324062 523292 324118
rect 523348 324062 523364 324118
rect 334444 324046 523364 324062
rect 334332 323938 464564 323954
rect 334332 323882 334348 323938
rect 334404 323882 464492 323938
rect 464548 323882 464564 323938
rect 334332 323866 464564 323882
rect 334444 322498 460308 322514
rect 334444 322442 334460 322498
rect 334516 322442 460236 322498
rect 460292 322442 460308 322498
rect 334444 322426 460308 322442
rect 334444 320878 404644 320894
rect 334444 320822 334460 320878
rect 334516 320822 404572 320878
rect 404628 320822 404644 320878
rect 334444 320806 404644 320822
rect 334444 319078 461204 319094
rect 334444 319022 334460 319078
rect 334516 319022 461132 319078
rect 461188 319022 461204 319078
rect 334444 319006 461204 319022
rect -1916 316350 597980 316446
rect -1916 316294 -1820 316350
rect -1764 316294 -1696 316350
rect -1640 316294 -1572 316350
rect -1516 316294 -1448 316350
rect -1392 316294 9234 316350
rect 9290 316294 9358 316350
rect 9414 316294 9482 316350
rect 9538 316294 9606 316350
rect 9662 316294 70674 316350
rect 70730 316294 70798 316350
rect 70854 316294 70922 316350
rect 70978 316294 71046 316350
rect 71102 316294 132114 316350
rect 132170 316294 132238 316350
rect 132294 316294 132362 316350
rect 132418 316294 132486 316350
rect 132542 316294 162834 316350
rect 162890 316294 162958 316350
rect 163014 316294 163082 316350
rect 163138 316294 163206 316350
rect 163262 316294 193554 316350
rect 193610 316294 193678 316350
rect 193734 316294 193802 316350
rect 193858 316294 193926 316350
rect 193982 316294 224274 316350
rect 224330 316294 224398 316350
rect 224454 316294 224522 316350
rect 224578 316294 224646 316350
rect 224702 316294 254994 316350
rect 255050 316294 255118 316350
rect 255174 316294 255242 316350
rect 255298 316294 255366 316350
rect 255422 316294 287878 316350
rect 287934 316294 288002 316350
rect 288058 316294 318598 316350
rect 318654 316294 318722 316350
rect 318778 316294 347154 316350
rect 347210 316294 347278 316350
rect 347334 316294 347402 316350
rect 347458 316294 347526 316350
rect 347582 316294 377874 316350
rect 377930 316294 377998 316350
rect 378054 316294 378122 316350
rect 378178 316294 378246 316350
rect 378302 316294 408594 316350
rect 408650 316294 408718 316350
rect 408774 316294 408842 316350
rect 408898 316294 408966 316350
rect 409022 316294 439314 316350
rect 439370 316294 439438 316350
rect 439494 316294 439562 316350
rect 439618 316294 439686 316350
rect 439742 316294 470034 316350
rect 470090 316294 470158 316350
rect 470214 316294 470282 316350
rect 470338 316294 470406 316350
rect 470462 316294 500754 316350
rect 500810 316294 500878 316350
rect 500934 316294 501002 316350
rect 501058 316294 501126 316350
rect 501182 316294 531474 316350
rect 531530 316294 531598 316350
rect 531654 316294 531722 316350
rect 531778 316294 531846 316350
rect 531902 316294 562194 316350
rect 562250 316294 562318 316350
rect 562374 316294 562442 316350
rect 562498 316294 562566 316350
rect 562622 316294 592914 316350
rect 592970 316294 593038 316350
rect 593094 316294 593162 316350
rect 593218 316294 593286 316350
rect 593342 316294 597456 316350
rect 597512 316294 597580 316350
rect 597636 316294 597704 316350
rect 597760 316294 597828 316350
rect 597884 316294 597980 316350
rect -1916 316226 597980 316294
rect -1916 316170 -1820 316226
rect -1764 316170 -1696 316226
rect -1640 316170 -1572 316226
rect -1516 316170 -1448 316226
rect -1392 316170 9234 316226
rect 9290 316170 9358 316226
rect 9414 316170 9482 316226
rect 9538 316170 9606 316226
rect 9662 316170 70674 316226
rect 70730 316170 70798 316226
rect 70854 316170 70922 316226
rect 70978 316170 71046 316226
rect 71102 316170 132114 316226
rect 132170 316170 132238 316226
rect 132294 316170 132362 316226
rect 132418 316170 132486 316226
rect 132542 316170 162834 316226
rect 162890 316170 162958 316226
rect 163014 316170 163082 316226
rect 163138 316170 163206 316226
rect 163262 316170 193554 316226
rect 193610 316170 193678 316226
rect 193734 316170 193802 316226
rect 193858 316170 193926 316226
rect 193982 316170 224274 316226
rect 224330 316170 224398 316226
rect 224454 316170 224522 316226
rect 224578 316170 224646 316226
rect 224702 316170 254994 316226
rect 255050 316170 255118 316226
rect 255174 316170 255242 316226
rect 255298 316170 255366 316226
rect 255422 316170 287878 316226
rect 287934 316170 288002 316226
rect 288058 316170 318598 316226
rect 318654 316170 318722 316226
rect 318778 316170 347154 316226
rect 347210 316170 347278 316226
rect 347334 316170 347402 316226
rect 347458 316170 347526 316226
rect 347582 316170 377874 316226
rect 377930 316170 377998 316226
rect 378054 316170 378122 316226
rect 378178 316170 378246 316226
rect 378302 316170 408594 316226
rect 408650 316170 408718 316226
rect 408774 316170 408842 316226
rect 408898 316170 408966 316226
rect 409022 316170 439314 316226
rect 439370 316170 439438 316226
rect 439494 316170 439562 316226
rect 439618 316170 439686 316226
rect 439742 316170 470034 316226
rect 470090 316170 470158 316226
rect 470214 316170 470282 316226
rect 470338 316170 470406 316226
rect 470462 316170 500754 316226
rect 500810 316170 500878 316226
rect 500934 316170 501002 316226
rect 501058 316170 501126 316226
rect 501182 316170 531474 316226
rect 531530 316170 531598 316226
rect 531654 316170 531722 316226
rect 531778 316170 531846 316226
rect 531902 316170 562194 316226
rect 562250 316170 562318 316226
rect 562374 316170 562442 316226
rect 562498 316170 562566 316226
rect 562622 316170 592914 316226
rect 592970 316170 593038 316226
rect 593094 316170 593162 316226
rect 593218 316170 593286 316226
rect 593342 316170 597456 316226
rect 597512 316170 597580 316226
rect 597636 316170 597704 316226
rect 597760 316170 597828 316226
rect 597884 316170 597980 316226
rect -1916 316102 597980 316170
rect -1916 316046 -1820 316102
rect -1764 316046 -1696 316102
rect -1640 316046 -1572 316102
rect -1516 316046 -1448 316102
rect -1392 316046 9234 316102
rect 9290 316046 9358 316102
rect 9414 316046 9482 316102
rect 9538 316046 9606 316102
rect 9662 316046 70674 316102
rect 70730 316046 70798 316102
rect 70854 316046 70922 316102
rect 70978 316046 71046 316102
rect 71102 316046 132114 316102
rect 132170 316046 132238 316102
rect 132294 316046 132362 316102
rect 132418 316046 132486 316102
rect 132542 316046 162834 316102
rect 162890 316046 162958 316102
rect 163014 316046 163082 316102
rect 163138 316046 163206 316102
rect 163262 316046 193554 316102
rect 193610 316046 193678 316102
rect 193734 316046 193802 316102
rect 193858 316046 193926 316102
rect 193982 316046 224274 316102
rect 224330 316046 224398 316102
rect 224454 316046 224522 316102
rect 224578 316046 224646 316102
rect 224702 316046 254994 316102
rect 255050 316046 255118 316102
rect 255174 316046 255242 316102
rect 255298 316046 255366 316102
rect 255422 316046 287878 316102
rect 287934 316046 288002 316102
rect 288058 316046 318598 316102
rect 318654 316046 318722 316102
rect 318778 316046 347154 316102
rect 347210 316046 347278 316102
rect 347334 316046 347402 316102
rect 347458 316046 347526 316102
rect 347582 316046 377874 316102
rect 377930 316046 377998 316102
rect 378054 316046 378122 316102
rect 378178 316046 378246 316102
rect 378302 316046 408594 316102
rect 408650 316046 408718 316102
rect 408774 316046 408842 316102
rect 408898 316046 408966 316102
rect 409022 316046 439314 316102
rect 439370 316046 439438 316102
rect 439494 316046 439562 316102
rect 439618 316046 439686 316102
rect 439742 316046 470034 316102
rect 470090 316046 470158 316102
rect 470214 316046 470282 316102
rect 470338 316046 470406 316102
rect 470462 316046 500754 316102
rect 500810 316046 500878 316102
rect 500934 316046 501002 316102
rect 501058 316046 501126 316102
rect 501182 316046 531474 316102
rect 531530 316046 531598 316102
rect 531654 316046 531722 316102
rect 531778 316046 531846 316102
rect 531902 316046 562194 316102
rect 562250 316046 562318 316102
rect 562374 316046 562442 316102
rect 562498 316046 562566 316102
rect 562622 316046 592914 316102
rect 592970 316046 593038 316102
rect 593094 316046 593162 316102
rect 593218 316046 593286 316102
rect 593342 316046 597456 316102
rect 597512 316046 597580 316102
rect 597636 316046 597704 316102
rect 597760 316046 597828 316102
rect 597884 316046 597980 316102
rect -1916 315978 597980 316046
rect -1916 315922 -1820 315978
rect -1764 315922 -1696 315978
rect -1640 315922 -1572 315978
rect -1516 315922 -1448 315978
rect -1392 315922 9234 315978
rect 9290 315922 9358 315978
rect 9414 315922 9482 315978
rect 9538 315922 9606 315978
rect 9662 315922 70674 315978
rect 70730 315922 70798 315978
rect 70854 315922 70922 315978
rect 70978 315922 71046 315978
rect 71102 315922 132114 315978
rect 132170 315922 132238 315978
rect 132294 315922 132362 315978
rect 132418 315922 132486 315978
rect 132542 315922 162834 315978
rect 162890 315922 162958 315978
rect 163014 315922 163082 315978
rect 163138 315922 163206 315978
rect 163262 315922 193554 315978
rect 193610 315922 193678 315978
rect 193734 315922 193802 315978
rect 193858 315922 193926 315978
rect 193982 315922 224274 315978
rect 224330 315922 224398 315978
rect 224454 315922 224522 315978
rect 224578 315922 224646 315978
rect 224702 315922 254994 315978
rect 255050 315922 255118 315978
rect 255174 315922 255242 315978
rect 255298 315922 255366 315978
rect 255422 315922 287878 315978
rect 287934 315922 288002 315978
rect 288058 315922 318598 315978
rect 318654 315922 318722 315978
rect 318778 315922 347154 315978
rect 347210 315922 347278 315978
rect 347334 315922 347402 315978
rect 347458 315922 347526 315978
rect 347582 315922 377874 315978
rect 377930 315922 377998 315978
rect 378054 315922 378122 315978
rect 378178 315922 378246 315978
rect 378302 315922 408594 315978
rect 408650 315922 408718 315978
rect 408774 315922 408842 315978
rect 408898 315922 408966 315978
rect 409022 315922 439314 315978
rect 439370 315922 439438 315978
rect 439494 315922 439562 315978
rect 439618 315922 439686 315978
rect 439742 315922 470034 315978
rect 470090 315922 470158 315978
rect 470214 315922 470282 315978
rect 470338 315922 470406 315978
rect 470462 315922 500754 315978
rect 500810 315922 500878 315978
rect 500934 315922 501002 315978
rect 501058 315922 501126 315978
rect 501182 315922 531474 315978
rect 531530 315922 531598 315978
rect 531654 315922 531722 315978
rect 531778 315922 531846 315978
rect 531902 315922 562194 315978
rect 562250 315922 562318 315978
rect 562374 315922 562442 315978
rect 562498 315922 562566 315978
rect 562622 315922 592914 315978
rect 592970 315922 593038 315978
rect 593094 315922 593162 315978
rect 593218 315922 593286 315978
rect 593342 315922 597456 315978
rect 597512 315922 597580 315978
rect 597636 315922 597704 315978
rect 597760 315922 597828 315978
rect 597884 315922 597980 315978
rect -1916 315826 597980 315922
rect 351916 314038 563012 314054
rect 351916 313982 351932 314038
rect 351988 313982 562940 314038
rect 562996 313982 563012 314038
rect 351916 313966 563012 313982
rect -1916 310350 597980 310446
rect -1916 310294 -860 310350
rect -804 310294 -736 310350
rect -680 310294 -612 310350
rect -556 310294 -488 310350
rect -432 310294 5514 310350
rect 5570 310294 5638 310350
rect 5694 310294 5762 310350
rect 5818 310294 5886 310350
rect 5942 310294 36234 310350
rect 36290 310294 36358 310350
rect 36414 310294 36482 310350
rect 36538 310294 36606 310350
rect 36662 310294 66954 310350
rect 67010 310294 67078 310350
rect 67134 310294 67202 310350
rect 67258 310294 67326 310350
rect 67382 310294 97674 310350
rect 97730 310294 97798 310350
rect 97854 310294 97922 310350
rect 97978 310294 98046 310350
rect 98102 310294 128394 310350
rect 128450 310294 128518 310350
rect 128574 310294 128642 310350
rect 128698 310294 128766 310350
rect 128822 310294 159114 310350
rect 159170 310294 159238 310350
rect 159294 310294 159362 310350
rect 159418 310294 159486 310350
rect 159542 310294 189834 310350
rect 189890 310294 189958 310350
rect 190014 310294 190082 310350
rect 190138 310294 190206 310350
rect 190262 310294 220554 310350
rect 220610 310294 220678 310350
rect 220734 310294 220802 310350
rect 220858 310294 220926 310350
rect 220982 310294 251274 310350
rect 251330 310294 251398 310350
rect 251454 310294 251522 310350
rect 251578 310294 251646 310350
rect 251702 310294 272518 310350
rect 272574 310294 272642 310350
rect 272698 310294 303238 310350
rect 303294 310294 303362 310350
rect 303418 310294 343434 310350
rect 343490 310294 343558 310350
rect 343614 310294 343682 310350
rect 343738 310294 343806 310350
rect 343862 310294 374154 310350
rect 374210 310294 374278 310350
rect 374334 310294 374402 310350
rect 374458 310294 374526 310350
rect 374582 310294 404874 310350
rect 404930 310294 404998 310350
rect 405054 310294 405122 310350
rect 405178 310294 405246 310350
rect 405302 310294 435594 310350
rect 435650 310294 435718 310350
rect 435774 310294 435842 310350
rect 435898 310294 435966 310350
rect 436022 310294 466314 310350
rect 466370 310294 466438 310350
rect 466494 310294 466562 310350
rect 466618 310294 466686 310350
rect 466742 310294 497034 310350
rect 497090 310294 497158 310350
rect 497214 310294 497282 310350
rect 497338 310294 497406 310350
rect 497462 310294 527754 310350
rect 527810 310294 527878 310350
rect 527934 310294 528002 310350
rect 528058 310294 528126 310350
rect 528182 310294 558474 310350
rect 558530 310294 558598 310350
rect 558654 310294 558722 310350
rect 558778 310294 558846 310350
rect 558902 310294 589194 310350
rect 589250 310294 589318 310350
rect 589374 310294 589442 310350
rect 589498 310294 589566 310350
rect 589622 310294 596496 310350
rect 596552 310294 596620 310350
rect 596676 310294 596744 310350
rect 596800 310294 596868 310350
rect 596924 310294 597980 310350
rect -1916 310226 597980 310294
rect -1916 310170 -860 310226
rect -804 310170 -736 310226
rect -680 310170 -612 310226
rect -556 310170 -488 310226
rect -432 310170 5514 310226
rect 5570 310170 5638 310226
rect 5694 310170 5762 310226
rect 5818 310170 5886 310226
rect 5942 310170 36234 310226
rect 36290 310170 36358 310226
rect 36414 310170 36482 310226
rect 36538 310170 36606 310226
rect 36662 310170 66954 310226
rect 67010 310170 67078 310226
rect 67134 310170 67202 310226
rect 67258 310170 67326 310226
rect 67382 310170 97674 310226
rect 97730 310170 97798 310226
rect 97854 310170 97922 310226
rect 97978 310170 98046 310226
rect 98102 310170 128394 310226
rect 128450 310170 128518 310226
rect 128574 310170 128642 310226
rect 128698 310170 128766 310226
rect 128822 310170 159114 310226
rect 159170 310170 159238 310226
rect 159294 310170 159362 310226
rect 159418 310170 159486 310226
rect 159542 310170 189834 310226
rect 189890 310170 189958 310226
rect 190014 310170 190082 310226
rect 190138 310170 190206 310226
rect 190262 310170 220554 310226
rect 220610 310170 220678 310226
rect 220734 310170 220802 310226
rect 220858 310170 220926 310226
rect 220982 310170 251274 310226
rect 251330 310170 251398 310226
rect 251454 310170 251522 310226
rect 251578 310170 251646 310226
rect 251702 310170 272518 310226
rect 272574 310170 272642 310226
rect 272698 310170 303238 310226
rect 303294 310170 303362 310226
rect 303418 310170 343434 310226
rect 343490 310170 343558 310226
rect 343614 310170 343682 310226
rect 343738 310170 343806 310226
rect 343862 310170 374154 310226
rect 374210 310170 374278 310226
rect 374334 310170 374402 310226
rect 374458 310170 374526 310226
rect 374582 310170 404874 310226
rect 404930 310170 404998 310226
rect 405054 310170 405122 310226
rect 405178 310170 405246 310226
rect 405302 310170 435594 310226
rect 435650 310170 435718 310226
rect 435774 310170 435842 310226
rect 435898 310170 435966 310226
rect 436022 310170 466314 310226
rect 466370 310170 466438 310226
rect 466494 310170 466562 310226
rect 466618 310170 466686 310226
rect 466742 310170 497034 310226
rect 497090 310170 497158 310226
rect 497214 310170 497282 310226
rect 497338 310170 497406 310226
rect 497462 310170 527754 310226
rect 527810 310170 527878 310226
rect 527934 310170 528002 310226
rect 528058 310170 528126 310226
rect 528182 310170 558474 310226
rect 558530 310170 558598 310226
rect 558654 310170 558722 310226
rect 558778 310170 558846 310226
rect 558902 310170 589194 310226
rect 589250 310170 589318 310226
rect 589374 310170 589442 310226
rect 589498 310170 589566 310226
rect 589622 310170 596496 310226
rect 596552 310170 596620 310226
rect 596676 310170 596744 310226
rect 596800 310170 596868 310226
rect 596924 310170 597980 310226
rect -1916 310102 597980 310170
rect -1916 310046 -860 310102
rect -804 310046 -736 310102
rect -680 310046 -612 310102
rect -556 310046 -488 310102
rect -432 310046 5514 310102
rect 5570 310046 5638 310102
rect 5694 310046 5762 310102
rect 5818 310046 5886 310102
rect 5942 310046 36234 310102
rect 36290 310046 36358 310102
rect 36414 310046 36482 310102
rect 36538 310046 36606 310102
rect 36662 310046 66954 310102
rect 67010 310046 67078 310102
rect 67134 310046 67202 310102
rect 67258 310046 67326 310102
rect 67382 310046 97674 310102
rect 97730 310046 97798 310102
rect 97854 310046 97922 310102
rect 97978 310046 98046 310102
rect 98102 310046 128394 310102
rect 128450 310046 128518 310102
rect 128574 310046 128642 310102
rect 128698 310046 128766 310102
rect 128822 310046 159114 310102
rect 159170 310046 159238 310102
rect 159294 310046 159362 310102
rect 159418 310046 159486 310102
rect 159542 310046 189834 310102
rect 189890 310046 189958 310102
rect 190014 310046 190082 310102
rect 190138 310046 190206 310102
rect 190262 310046 220554 310102
rect 220610 310046 220678 310102
rect 220734 310046 220802 310102
rect 220858 310046 220926 310102
rect 220982 310046 251274 310102
rect 251330 310046 251398 310102
rect 251454 310046 251522 310102
rect 251578 310046 251646 310102
rect 251702 310046 272518 310102
rect 272574 310046 272642 310102
rect 272698 310046 303238 310102
rect 303294 310046 303362 310102
rect 303418 310046 343434 310102
rect 343490 310046 343558 310102
rect 343614 310046 343682 310102
rect 343738 310046 343806 310102
rect 343862 310046 374154 310102
rect 374210 310046 374278 310102
rect 374334 310046 374402 310102
rect 374458 310046 374526 310102
rect 374582 310046 404874 310102
rect 404930 310046 404998 310102
rect 405054 310046 405122 310102
rect 405178 310046 405246 310102
rect 405302 310046 435594 310102
rect 435650 310046 435718 310102
rect 435774 310046 435842 310102
rect 435898 310046 435966 310102
rect 436022 310046 466314 310102
rect 466370 310046 466438 310102
rect 466494 310046 466562 310102
rect 466618 310046 466686 310102
rect 466742 310046 497034 310102
rect 497090 310046 497158 310102
rect 497214 310046 497282 310102
rect 497338 310046 497406 310102
rect 497462 310046 527754 310102
rect 527810 310046 527878 310102
rect 527934 310046 528002 310102
rect 528058 310046 528126 310102
rect 528182 310046 558474 310102
rect 558530 310046 558598 310102
rect 558654 310046 558722 310102
rect 558778 310046 558846 310102
rect 558902 310046 589194 310102
rect 589250 310046 589318 310102
rect 589374 310046 589442 310102
rect 589498 310046 589566 310102
rect 589622 310046 596496 310102
rect 596552 310046 596620 310102
rect 596676 310046 596744 310102
rect 596800 310046 596868 310102
rect 596924 310046 597980 310102
rect -1916 309978 597980 310046
rect -1916 309922 -860 309978
rect -804 309922 -736 309978
rect -680 309922 -612 309978
rect -556 309922 -488 309978
rect -432 309922 5514 309978
rect 5570 309922 5638 309978
rect 5694 309922 5762 309978
rect 5818 309922 5886 309978
rect 5942 309922 36234 309978
rect 36290 309922 36358 309978
rect 36414 309922 36482 309978
rect 36538 309922 36606 309978
rect 36662 309922 66954 309978
rect 67010 309922 67078 309978
rect 67134 309922 67202 309978
rect 67258 309922 67326 309978
rect 67382 309922 97674 309978
rect 97730 309922 97798 309978
rect 97854 309922 97922 309978
rect 97978 309922 98046 309978
rect 98102 309922 128394 309978
rect 128450 309922 128518 309978
rect 128574 309922 128642 309978
rect 128698 309922 128766 309978
rect 128822 309922 159114 309978
rect 159170 309922 159238 309978
rect 159294 309922 159362 309978
rect 159418 309922 159486 309978
rect 159542 309922 189834 309978
rect 189890 309922 189958 309978
rect 190014 309922 190082 309978
rect 190138 309922 190206 309978
rect 190262 309922 220554 309978
rect 220610 309922 220678 309978
rect 220734 309922 220802 309978
rect 220858 309922 220926 309978
rect 220982 309922 251274 309978
rect 251330 309922 251398 309978
rect 251454 309922 251522 309978
rect 251578 309922 251646 309978
rect 251702 309922 272518 309978
rect 272574 309922 272642 309978
rect 272698 309922 303238 309978
rect 303294 309922 303362 309978
rect 303418 309922 343434 309978
rect 343490 309922 343558 309978
rect 343614 309922 343682 309978
rect 343738 309922 343806 309978
rect 343862 309922 374154 309978
rect 374210 309922 374278 309978
rect 374334 309922 374402 309978
rect 374458 309922 374526 309978
rect 374582 309922 404874 309978
rect 404930 309922 404998 309978
rect 405054 309922 405122 309978
rect 405178 309922 405246 309978
rect 405302 309922 435594 309978
rect 435650 309922 435718 309978
rect 435774 309922 435842 309978
rect 435898 309922 435966 309978
rect 436022 309922 466314 309978
rect 466370 309922 466438 309978
rect 466494 309922 466562 309978
rect 466618 309922 466686 309978
rect 466742 309922 497034 309978
rect 497090 309922 497158 309978
rect 497214 309922 497282 309978
rect 497338 309922 497406 309978
rect 497462 309922 527754 309978
rect 527810 309922 527878 309978
rect 527934 309922 528002 309978
rect 528058 309922 528126 309978
rect 528182 309922 558474 309978
rect 558530 309922 558598 309978
rect 558654 309922 558722 309978
rect 558778 309922 558846 309978
rect 558902 309922 589194 309978
rect 589250 309922 589318 309978
rect 589374 309922 589442 309978
rect 589498 309922 589566 309978
rect 589622 309922 596496 309978
rect 596552 309922 596620 309978
rect 596676 309922 596744 309978
rect 596800 309922 596868 309978
rect 596924 309922 597980 309978
rect -1916 309826 597980 309922
rect -1916 298350 597980 298446
rect -1916 298294 -1820 298350
rect -1764 298294 -1696 298350
rect -1640 298294 -1572 298350
rect -1516 298294 -1448 298350
rect -1392 298294 9234 298350
rect 9290 298294 9358 298350
rect 9414 298294 9482 298350
rect 9538 298294 9606 298350
rect 9662 298294 70674 298350
rect 70730 298294 70798 298350
rect 70854 298294 70922 298350
rect 70978 298294 71046 298350
rect 71102 298294 132114 298350
rect 132170 298294 132238 298350
rect 132294 298294 132362 298350
rect 132418 298294 132486 298350
rect 132542 298294 162834 298350
rect 162890 298294 162958 298350
rect 163014 298294 163082 298350
rect 163138 298294 163206 298350
rect 163262 298294 193554 298350
rect 193610 298294 193678 298350
rect 193734 298294 193802 298350
rect 193858 298294 193926 298350
rect 193982 298294 224274 298350
rect 224330 298294 224398 298350
rect 224454 298294 224522 298350
rect 224578 298294 224646 298350
rect 224702 298294 254994 298350
rect 255050 298294 255118 298350
rect 255174 298294 255242 298350
rect 255298 298294 255366 298350
rect 255422 298294 287878 298350
rect 287934 298294 288002 298350
rect 288058 298294 318598 298350
rect 318654 298294 318722 298350
rect 318778 298294 347154 298350
rect 347210 298294 347278 298350
rect 347334 298294 347402 298350
rect 347458 298294 347526 298350
rect 347582 298294 377874 298350
rect 377930 298294 377998 298350
rect 378054 298294 378122 298350
rect 378178 298294 378246 298350
rect 378302 298294 408594 298350
rect 408650 298294 408718 298350
rect 408774 298294 408842 298350
rect 408898 298294 408966 298350
rect 409022 298294 439314 298350
rect 439370 298294 439438 298350
rect 439494 298294 439562 298350
rect 439618 298294 439686 298350
rect 439742 298294 470034 298350
rect 470090 298294 470158 298350
rect 470214 298294 470282 298350
rect 470338 298294 470406 298350
rect 470462 298294 500754 298350
rect 500810 298294 500878 298350
rect 500934 298294 501002 298350
rect 501058 298294 501126 298350
rect 501182 298294 531474 298350
rect 531530 298294 531598 298350
rect 531654 298294 531722 298350
rect 531778 298294 531846 298350
rect 531902 298294 562194 298350
rect 562250 298294 562318 298350
rect 562374 298294 562442 298350
rect 562498 298294 562566 298350
rect 562622 298294 592914 298350
rect 592970 298294 593038 298350
rect 593094 298294 593162 298350
rect 593218 298294 593286 298350
rect 593342 298294 597456 298350
rect 597512 298294 597580 298350
rect 597636 298294 597704 298350
rect 597760 298294 597828 298350
rect 597884 298294 597980 298350
rect -1916 298226 597980 298294
rect -1916 298170 -1820 298226
rect -1764 298170 -1696 298226
rect -1640 298170 -1572 298226
rect -1516 298170 -1448 298226
rect -1392 298170 9234 298226
rect 9290 298170 9358 298226
rect 9414 298170 9482 298226
rect 9538 298170 9606 298226
rect 9662 298170 70674 298226
rect 70730 298170 70798 298226
rect 70854 298170 70922 298226
rect 70978 298170 71046 298226
rect 71102 298170 132114 298226
rect 132170 298170 132238 298226
rect 132294 298170 132362 298226
rect 132418 298170 132486 298226
rect 132542 298170 162834 298226
rect 162890 298170 162958 298226
rect 163014 298170 163082 298226
rect 163138 298170 163206 298226
rect 163262 298170 193554 298226
rect 193610 298170 193678 298226
rect 193734 298170 193802 298226
rect 193858 298170 193926 298226
rect 193982 298170 224274 298226
rect 224330 298170 224398 298226
rect 224454 298170 224522 298226
rect 224578 298170 224646 298226
rect 224702 298170 254994 298226
rect 255050 298170 255118 298226
rect 255174 298170 255242 298226
rect 255298 298170 255366 298226
rect 255422 298170 287878 298226
rect 287934 298170 288002 298226
rect 288058 298170 318598 298226
rect 318654 298170 318722 298226
rect 318778 298170 347154 298226
rect 347210 298170 347278 298226
rect 347334 298170 347402 298226
rect 347458 298170 347526 298226
rect 347582 298170 377874 298226
rect 377930 298170 377998 298226
rect 378054 298170 378122 298226
rect 378178 298170 378246 298226
rect 378302 298170 408594 298226
rect 408650 298170 408718 298226
rect 408774 298170 408842 298226
rect 408898 298170 408966 298226
rect 409022 298170 439314 298226
rect 439370 298170 439438 298226
rect 439494 298170 439562 298226
rect 439618 298170 439686 298226
rect 439742 298170 470034 298226
rect 470090 298170 470158 298226
rect 470214 298170 470282 298226
rect 470338 298170 470406 298226
rect 470462 298170 500754 298226
rect 500810 298170 500878 298226
rect 500934 298170 501002 298226
rect 501058 298170 501126 298226
rect 501182 298170 531474 298226
rect 531530 298170 531598 298226
rect 531654 298170 531722 298226
rect 531778 298170 531846 298226
rect 531902 298170 562194 298226
rect 562250 298170 562318 298226
rect 562374 298170 562442 298226
rect 562498 298170 562566 298226
rect 562622 298170 592914 298226
rect 592970 298170 593038 298226
rect 593094 298170 593162 298226
rect 593218 298170 593286 298226
rect 593342 298170 597456 298226
rect 597512 298170 597580 298226
rect 597636 298170 597704 298226
rect 597760 298170 597828 298226
rect 597884 298170 597980 298226
rect -1916 298102 597980 298170
rect -1916 298046 -1820 298102
rect -1764 298046 -1696 298102
rect -1640 298046 -1572 298102
rect -1516 298046 -1448 298102
rect -1392 298046 9234 298102
rect 9290 298046 9358 298102
rect 9414 298046 9482 298102
rect 9538 298046 9606 298102
rect 9662 298046 70674 298102
rect 70730 298046 70798 298102
rect 70854 298046 70922 298102
rect 70978 298046 71046 298102
rect 71102 298046 132114 298102
rect 132170 298046 132238 298102
rect 132294 298046 132362 298102
rect 132418 298046 132486 298102
rect 132542 298046 162834 298102
rect 162890 298046 162958 298102
rect 163014 298046 163082 298102
rect 163138 298046 163206 298102
rect 163262 298046 193554 298102
rect 193610 298046 193678 298102
rect 193734 298046 193802 298102
rect 193858 298046 193926 298102
rect 193982 298046 224274 298102
rect 224330 298046 224398 298102
rect 224454 298046 224522 298102
rect 224578 298046 224646 298102
rect 224702 298046 254994 298102
rect 255050 298046 255118 298102
rect 255174 298046 255242 298102
rect 255298 298046 255366 298102
rect 255422 298046 287878 298102
rect 287934 298046 288002 298102
rect 288058 298046 318598 298102
rect 318654 298046 318722 298102
rect 318778 298046 347154 298102
rect 347210 298046 347278 298102
rect 347334 298046 347402 298102
rect 347458 298046 347526 298102
rect 347582 298046 377874 298102
rect 377930 298046 377998 298102
rect 378054 298046 378122 298102
rect 378178 298046 378246 298102
rect 378302 298046 408594 298102
rect 408650 298046 408718 298102
rect 408774 298046 408842 298102
rect 408898 298046 408966 298102
rect 409022 298046 439314 298102
rect 439370 298046 439438 298102
rect 439494 298046 439562 298102
rect 439618 298046 439686 298102
rect 439742 298046 470034 298102
rect 470090 298046 470158 298102
rect 470214 298046 470282 298102
rect 470338 298046 470406 298102
rect 470462 298046 500754 298102
rect 500810 298046 500878 298102
rect 500934 298046 501002 298102
rect 501058 298046 501126 298102
rect 501182 298046 531474 298102
rect 531530 298046 531598 298102
rect 531654 298046 531722 298102
rect 531778 298046 531846 298102
rect 531902 298046 562194 298102
rect 562250 298046 562318 298102
rect 562374 298046 562442 298102
rect 562498 298046 562566 298102
rect 562622 298046 592914 298102
rect 592970 298046 593038 298102
rect 593094 298046 593162 298102
rect 593218 298046 593286 298102
rect 593342 298046 597456 298102
rect 597512 298046 597580 298102
rect 597636 298046 597704 298102
rect 597760 298046 597828 298102
rect 597884 298046 597980 298102
rect -1916 297978 597980 298046
rect -1916 297922 -1820 297978
rect -1764 297922 -1696 297978
rect -1640 297922 -1572 297978
rect -1516 297922 -1448 297978
rect -1392 297922 9234 297978
rect 9290 297922 9358 297978
rect 9414 297922 9482 297978
rect 9538 297922 9606 297978
rect 9662 297922 70674 297978
rect 70730 297922 70798 297978
rect 70854 297922 70922 297978
rect 70978 297922 71046 297978
rect 71102 297922 132114 297978
rect 132170 297922 132238 297978
rect 132294 297922 132362 297978
rect 132418 297922 132486 297978
rect 132542 297922 162834 297978
rect 162890 297922 162958 297978
rect 163014 297922 163082 297978
rect 163138 297922 163206 297978
rect 163262 297922 193554 297978
rect 193610 297922 193678 297978
rect 193734 297922 193802 297978
rect 193858 297922 193926 297978
rect 193982 297922 224274 297978
rect 224330 297922 224398 297978
rect 224454 297922 224522 297978
rect 224578 297922 224646 297978
rect 224702 297922 254994 297978
rect 255050 297922 255118 297978
rect 255174 297922 255242 297978
rect 255298 297922 255366 297978
rect 255422 297922 287878 297978
rect 287934 297922 288002 297978
rect 288058 297922 318598 297978
rect 318654 297922 318722 297978
rect 318778 297922 347154 297978
rect 347210 297922 347278 297978
rect 347334 297922 347402 297978
rect 347458 297922 347526 297978
rect 347582 297922 377874 297978
rect 377930 297922 377998 297978
rect 378054 297922 378122 297978
rect 378178 297922 378246 297978
rect 378302 297922 408594 297978
rect 408650 297922 408718 297978
rect 408774 297922 408842 297978
rect 408898 297922 408966 297978
rect 409022 297922 439314 297978
rect 439370 297922 439438 297978
rect 439494 297922 439562 297978
rect 439618 297922 439686 297978
rect 439742 297922 470034 297978
rect 470090 297922 470158 297978
rect 470214 297922 470282 297978
rect 470338 297922 470406 297978
rect 470462 297922 500754 297978
rect 500810 297922 500878 297978
rect 500934 297922 501002 297978
rect 501058 297922 501126 297978
rect 501182 297922 531474 297978
rect 531530 297922 531598 297978
rect 531654 297922 531722 297978
rect 531778 297922 531846 297978
rect 531902 297922 562194 297978
rect 562250 297922 562318 297978
rect 562374 297922 562442 297978
rect 562498 297922 562566 297978
rect 562622 297922 592914 297978
rect 592970 297922 593038 297978
rect 593094 297922 593162 297978
rect 593218 297922 593286 297978
rect 593342 297922 597456 297978
rect 597512 297922 597580 297978
rect 597636 297922 597704 297978
rect 597760 297922 597828 297978
rect 597884 297922 597980 297978
rect -1916 297826 597980 297922
rect -1916 292350 597980 292446
rect -1916 292294 -860 292350
rect -804 292294 -736 292350
rect -680 292294 -612 292350
rect -556 292294 -488 292350
rect -432 292294 5514 292350
rect 5570 292294 5638 292350
rect 5694 292294 5762 292350
rect 5818 292294 5886 292350
rect 5942 292294 36234 292350
rect 36290 292294 36358 292350
rect 36414 292294 36482 292350
rect 36538 292294 36606 292350
rect 36662 292294 66954 292350
rect 67010 292294 67078 292350
rect 67134 292294 67202 292350
rect 67258 292294 67326 292350
rect 67382 292294 97674 292350
rect 97730 292294 97798 292350
rect 97854 292294 97922 292350
rect 97978 292294 98046 292350
rect 98102 292294 128394 292350
rect 128450 292294 128518 292350
rect 128574 292294 128642 292350
rect 128698 292294 128766 292350
rect 128822 292294 159114 292350
rect 159170 292294 159238 292350
rect 159294 292294 159362 292350
rect 159418 292294 159486 292350
rect 159542 292294 189834 292350
rect 189890 292294 189958 292350
rect 190014 292294 190082 292350
rect 190138 292294 190206 292350
rect 190262 292294 220554 292350
rect 220610 292294 220678 292350
rect 220734 292294 220802 292350
rect 220858 292294 220926 292350
rect 220982 292294 251274 292350
rect 251330 292294 251398 292350
rect 251454 292294 251522 292350
rect 251578 292294 251646 292350
rect 251702 292294 272518 292350
rect 272574 292294 272642 292350
rect 272698 292294 303238 292350
rect 303294 292294 303362 292350
rect 303418 292294 343434 292350
rect 343490 292294 343558 292350
rect 343614 292294 343682 292350
rect 343738 292294 343806 292350
rect 343862 292294 374154 292350
rect 374210 292294 374278 292350
rect 374334 292294 374402 292350
rect 374458 292294 374526 292350
rect 374582 292294 404874 292350
rect 404930 292294 404998 292350
rect 405054 292294 405122 292350
rect 405178 292294 405246 292350
rect 405302 292294 435594 292350
rect 435650 292294 435718 292350
rect 435774 292294 435842 292350
rect 435898 292294 435966 292350
rect 436022 292294 466314 292350
rect 466370 292294 466438 292350
rect 466494 292294 466562 292350
rect 466618 292294 466686 292350
rect 466742 292294 497034 292350
rect 497090 292294 497158 292350
rect 497214 292294 497282 292350
rect 497338 292294 497406 292350
rect 497462 292294 527754 292350
rect 527810 292294 527878 292350
rect 527934 292294 528002 292350
rect 528058 292294 528126 292350
rect 528182 292294 558474 292350
rect 558530 292294 558598 292350
rect 558654 292294 558722 292350
rect 558778 292294 558846 292350
rect 558902 292294 589194 292350
rect 589250 292294 589318 292350
rect 589374 292294 589442 292350
rect 589498 292294 589566 292350
rect 589622 292294 596496 292350
rect 596552 292294 596620 292350
rect 596676 292294 596744 292350
rect 596800 292294 596868 292350
rect 596924 292294 597980 292350
rect -1916 292226 597980 292294
rect -1916 292170 -860 292226
rect -804 292170 -736 292226
rect -680 292170 -612 292226
rect -556 292170 -488 292226
rect -432 292170 5514 292226
rect 5570 292170 5638 292226
rect 5694 292170 5762 292226
rect 5818 292170 5886 292226
rect 5942 292170 36234 292226
rect 36290 292170 36358 292226
rect 36414 292170 36482 292226
rect 36538 292170 36606 292226
rect 36662 292170 66954 292226
rect 67010 292170 67078 292226
rect 67134 292170 67202 292226
rect 67258 292170 67326 292226
rect 67382 292170 97674 292226
rect 97730 292170 97798 292226
rect 97854 292170 97922 292226
rect 97978 292170 98046 292226
rect 98102 292170 128394 292226
rect 128450 292170 128518 292226
rect 128574 292170 128642 292226
rect 128698 292170 128766 292226
rect 128822 292170 159114 292226
rect 159170 292170 159238 292226
rect 159294 292170 159362 292226
rect 159418 292170 159486 292226
rect 159542 292170 189834 292226
rect 189890 292170 189958 292226
rect 190014 292170 190082 292226
rect 190138 292170 190206 292226
rect 190262 292170 220554 292226
rect 220610 292170 220678 292226
rect 220734 292170 220802 292226
rect 220858 292170 220926 292226
rect 220982 292170 251274 292226
rect 251330 292170 251398 292226
rect 251454 292170 251522 292226
rect 251578 292170 251646 292226
rect 251702 292170 272518 292226
rect 272574 292170 272642 292226
rect 272698 292170 303238 292226
rect 303294 292170 303362 292226
rect 303418 292170 343434 292226
rect 343490 292170 343558 292226
rect 343614 292170 343682 292226
rect 343738 292170 343806 292226
rect 343862 292170 374154 292226
rect 374210 292170 374278 292226
rect 374334 292170 374402 292226
rect 374458 292170 374526 292226
rect 374582 292170 404874 292226
rect 404930 292170 404998 292226
rect 405054 292170 405122 292226
rect 405178 292170 405246 292226
rect 405302 292170 435594 292226
rect 435650 292170 435718 292226
rect 435774 292170 435842 292226
rect 435898 292170 435966 292226
rect 436022 292170 466314 292226
rect 466370 292170 466438 292226
rect 466494 292170 466562 292226
rect 466618 292170 466686 292226
rect 466742 292170 497034 292226
rect 497090 292170 497158 292226
rect 497214 292170 497282 292226
rect 497338 292170 497406 292226
rect 497462 292170 527754 292226
rect 527810 292170 527878 292226
rect 527934 292170 528002 292226
rect 528058 292170 528126 292226
rect 528182 292170 558474 292226
rect 558530 292170 558598 292226
rect 558654 292170 558722 292226
rect 558778 292170 558846 292226
rect 558902 292170 589194 292226
rect 589250 292170 589318 292226
rect 589374 292170 589442 292226
rect 589498 292170 589566 292226
rect 589622 292170 596496 292226
rect 596552 292170 596620 292226
rect 596676 292170 596744 292226
rect 596800 292170 596868 292226
rect 596924 292170 597980 292226
rect -1916 292102 597980 292170
rect -1916 292046 -860 292102
rect -804 292046 -736 292102
rect -680 292046 -612 292102
rect -556 292046 -488 292102
rect -432 292046 5514 292102
rect 5570 292046 5638 292102
rect 5694 292046 5762 292102
rect 5818 292046 5886 292102
rect 5942 292046 36234 292102
rect 36290 292046 36358 292102
rect 36414 292046 36482 292102
rect 36538 292046 36606 292102
rect 36662 292046 66954 292102
rect 67010 292046 67078 292102
rect 67134 292046 67202 292102
rect 67258 292046 67326 292102
rect 67382 292046 97674 292102
rect 97730 292046 97798 292102
rect 97854 292046 97922 292102
rect 97978 292046 98046 292102
rect 98102 292046 128394 292102
rect 128450 292046 128518 292102
rect 128574 292046 128642 292102
rect 128698 292046 128766 292102
rect 128822 292046 159114 292102
rect 159170 292046 159238 292102
rect 159294 292046 159362 292102
rect 159418 292046 159486 292102
rect 159542 292046 189834 292102
rect 189890 292046 189958 292102
rect 190014 292046 190082 292102
rect 190138 292046 190206 292102
rect 190262 292046 220554 292102
rect 220610 292046 220678 292102
rect 220734 292046 220802 292102
rect 220858 292046 220926 292102
rect 220982 292046 251274 292102
rect 251330 292046 251398 292102
rect 251454 292046 251522 292102
rect 251578 292046 251646 292102
rect 251702 292046 272518 292102
rect 272574 292046 272642 292102
rect 272698 292046 303238 292102
rect 303294 292046 303362 292102
rect 303418 292046 343434 292102
rect 343490 292046 343558 292102
rect 343614 292046 343682 292102
rect 343738 292046 343806 292102
rect 343862 292046 374154 292102
rect 374210 292046 374278 292102
rect 374334 292046 374402 292102
rect 374458 292046 374526 292102
rect 374582 292046 404874 292102
rect 404930 292046 404998 292102
rect 405054 292046 405122 292102
rect 405178 292046 405246 292102
rect 405302 292046 435594 292102
rect 435650 292046 435718 292102
rect 435774 292046 435842 292102
rect 435898 292046 435966 292102
rect 436022 292046 466314 292102
rect 466370 292046 466438 292102
rect 466494 292046 466562 292102
rect 466618 292046 466686 292102
rect 466742 292046 497034 292102
rect 497090 292046 497158 292102
rect 497214 292046 497282 292102
rect 497338 292046 497406 292102
rect 497462 292046 527754 292102
rect 527810 292046 527878 292102
rect 527934 292046 528002 292102
rect 528058 292046 528126 292102
rect 528182 292046 558474 292102
rect 558530 292046 558598 292102
rect 558654 292046 558722 292102
rect 558778 292046 558846 292102
rect 558902 292046 589194 292102
rect 589250 292046 589318 292102
rect 589374 292046 589442 292102
rect 589498 292046 589566 292102
rect 589622 292046 596496 292102
rect 596552 292046 596620 292102
rect 596676 292046 596744 292102
rect 596800 292046 596868 292102
rect 596924 292046 597980 292102
rect -1916 291978 597980 292046
rect -1916 291922 -860 291978
rect -804 291922 -736 291978
rect -680 291922 -612 291978
rect -556 291922 -488 291978
rect -432 291922 5514 291978
rect 5570 291922 5638 291978
rect 5694 291922 5762 291978
rect 5818 291922 5886 291978
rect 5942 291922 36234 291978
rect 36290 291922 36358 291978
rect 36414 291922 36482 291978
rect 36538 291922 36606 291978
rect 36662 291922 66954 291978
rect 67010 291922 67078 291978
rect 67134 291922 67202 291978
rect 67258 291922 67326 291978
rect 67382 291922 97674 291978
rect 97730 291922 97798 291978
rect 97854 291922 97922 291978
rect 97978 291922 98046 291978
rect 98102 291922 128394 291978
rect 128450 291922 128518 291978
rect 128574 291922 128642 291978
rect 128698 291922 128766 291978
rect 128822 291922 159114 291978
rect 159170 291922 159238 291978
rect 159294 291922 159362 291978
rect 159418 291922 159486 291978
rect 159542 291922 189834 291978
rect 189890 291922 189958 291978
rect 190014 291922 190082 291978
rect 190138 291922 190206 291978
rect 190262 291922 220554 291978
rect 220610 291922 220678 291978
rect 220734 291922 220802 291978
rect 220858 291922 220926 291978
rect 220982 291922 251274 291978
rect 251330 291922 251398 291978
rect 251454 291922 251522 291978
rect 251578 291922 251646 291978
rect 251702 291922 272518 291978
rect 272574 291922 272642 291978
rect 272698 291922 303238 291978
rect 303294 291922 303362 291978
rect 303418 291922 343434 291978
rect 343490 291922 343558 291978
rect 343614 291922 343682 291978
rect 343738 291922 343806 291978
rect 343862 291922 374154 291978
rect 374210 291922 374278 291978
rect 374334 291922 374402 291978
rect 374458 291922 374526 291978
rect 374582 291922 404874 291978
rect 404930 291922 404998 291978
rect 405054 291922 405122 291978
rect 405178 291922 405246 291978
rect 405302 291922 435594 291978
rect 435650 291922 435718 291978
rect 435774 291922 435842 291978
rect 435898 291922 435966 291978
rect 436022 291922 466314 291978
rect 466370 291922 466438 291978
rect 466494 291922 466562 291978
rect 466618 291922 466686 291978
rect 466742 291922 497034 291978
rect 497090 291922 497158 291978
rect 497214 291922 497282 291978
rect 497338 291922 497406 291978
rect 497462 291922 527754 291978
rect 527810 291922 527878 291978
rect 527934 291922 528002 291978
rect 528058 291922 528126 291978
rect 528182 291922 558474 291978
rect 558530 291922 558598 291978
rect 558654 291922 558722 291978
rect 558778 291922 558846 291978
rect 558902 291922 589194 291978
rect 589250 291922 589318 291978
rect 589374 291922 589442 291978
rect 589498 291922 589566 291978
rect 589622 291922 596496 291978
rect 596552 291922 596620 291978
rect 596676 291922 596744 291978
rect 596800 291922 596868 291978
rect 596924 291922 597980 291978
rect -1916 291826 597980 291922
rect -1916 280350 597980 280446
rect -1916 280294 -1820 280350
rect -1764 280294 -1696 280350
rect -1640 280294 -1572 280350
rect -1516 280294 -1448 280350
rect -1392 280294 9234 280350
rect 9290 280294 9358 280350
rect 9414 280294 9482 280350
rect 9538 280294 9606 280350
rect 9662 280294 39878 280350
rect 39934 280294 40002 280350
rect 40058 280294 70674 280350
rect 70730 280294 70798 280350
rect 70854 280294 70922 280350
rect 70978 280294 71046 280350
rect 71102 280294 101878 280350
rect 101934 280294 102002 280350
rect 102058 280294 132114 280350
rect 132170 280294 132238 280350
rect 132294 280294 132362 280350
rect 132418 280294 132486 280350
rect 132542 280294 162834 280350
rect 162890 280294 162958 280350
rect 163014 280294 163082 280350
rect 163138 280294 163206 280350
rect 163262 280294 163878 280350
rect 163934 280294 164002 280350
rect 164058 280294 193554 280350
rect 193610 280294 193678 280350
rect 193734 280294 193802 280350
rect 193858 280294 193926 280350
rect 193982 280294 224274 280350
rect 224330 280294 224398 280350
rect 224454 280294 224522 280350
rect 224578 280294 224646 280350
rect 224702 280294 225878 280350
rect 225934 280294 226002 280350
rect 226058 280294 254994 280350
rect 255050 280294 255118 280350
rect 255174 280294 255242 280350
rect 255298 280294 255366 280350
rect 255422 280294 287878 280350
rect 287934 280294 288002 280350
rect 288058 280294 318598 280350
rect 318654 280294 318722 280350
rect 318778 280294 347154 280350
rect 347210 280294 347278 280350
rect 347334 280294 347402 280350
rect 347458 280294 347526 280350
rect 347582 280294 371878 280350
rect 371934 280294 372002 280350
rect 372058 280294 377874 280350
rect 377930 280294 377998 280350
rect 378054 280294 378122 280350
rect 378178 280294 378246 280350
rect 378302 280294 408594 280350
rect 408650 280294 408718 280350
rect 408774 280294 408842 280350
rect 408898 280294 408966 280350
rect 409022 280294 433878 280350
rect 433934 280294 434002 280350
rect 434058 280294 439314 280350
rect 439370 280294 439438 280350
rect 439494 280294 439562 280350
rect 439618 280294 439686 280350
rect 439742 280294 470034 280350
rect 470090 280294 470158 280350
rect 470214 280294 470282 280350
rect 470338 280294 470406 280350
rect 470462 280294 495878 280350
rect 495934 280294 496002 280350
rect 496058 280294 500754 280350
rect 500810 280294 500878 280350
rect 500934 280294 501002 280350
rect 501058 280294 501126 280350
rect 501182 280294 531474 280350
rect 531530 280294 531598 280350
rect 531654 280294 531722 280350
rect 531778 280294 531846 280350
rect 531902 280294 557878 280350
rect 557934 280294 558002 280350
rect 558058 280294 562194 280350
rect 562250 280294 562318 280350
rect 562374 280294 562442 280350
rect 562498 280294 562566 280350
rect 562622 280294 592914 280350
rect 592970 280294 593038 280350
rect 593094 280294 593162 280350
rect 593218 280294 593286 280350
rect 593342 280294 597456 280350
rect 597512 280294 597580 280350
rect 597636 280294 597704 280350
rect 597760 280294 597828 280350
rect 597884 280294 597980 280350
rect -1916 280226 597980 280294
rect -1916 280170 -1820 280226
rect -1764 280170 -1696 280226
rect -1640 280170 -1572 280226
rect -1516 280170 -1448 280226
rect -1392 280170 9234 280226
rect 9290 280170 9358 280226
rect 9414 280170 9482 280226
rect 9538 280170 9606 280226
rect 9662 280170 39878 280226
rect 39934 280170 40002 280226
rect 40058 280170 70674 280226
rect 70730 280170 70798 280226
rect 70854 280170 70922 280226
rect 70978 280170 71046 280226
rect 71102 280170 101878 280226
rect 101934 280170 102002 280226
rect 102058 280170 132114 280226
rect 132170 280170 132238 280226
rect 132294 280170 132362 280226
rect 132418 280170 132486 280226
rect 132542 280170 162834 280226
rect 162890 280170 162958 280226
rect 163014 280170 163082 280226
rect 163138 280170 163206 280226
rect 163262 280170 163878 280226
rect 163934 280170 164002 280226
rect 164058 280170 193554 280226
rect 193610 280170 193678 280226
rect 193734 280170 193802 280226
rect 193858 280170 193926 280226
rect 193982 280170 224274 280226
rect 224330 280170 224398 280226
rect 224454 280170 224522 280226
rect 224578 280170 224646 280226
rect 224702 280170 225878 280226
rect 225934 280170 226002 280226
rect 226058 280170 254994 280226
rect 255050 280170 255118 280226
rect 255174 280170 255242 280226
rect 255298 280170 255366 280226
rect 255422 280170 287878 280226
rect 287934 280170 288002 280226
rect 288058 280170 318598 280226
rect 318654 280170 318722 280226
rect 318778 280170 347154 280226
rect 347210 280170 347278 280226
rect 347334 280170 347402 280226
rect 347458 280170 347526 280226
rect 347582 280170 371878 280226
rect 371934 280170 372002 280226
rect 372058 280170 377874 280226
rect 377930 280170 377998 280226
rect 378054 280170 378122 280226
rect 378178 280170 378246 280226
rect 378302 280170 408594 280226
rect 408650 280170 408718 280226
rect 408774 280170 408842 280226
rect 408898 280170 408966 280226
rect 409022 280170 433878 280226
rect 433934 280170 434002 280226
rect 434058 280170 439314 280226
rect 439370 280170 439438 280226
rect 439494 280170 439562 280226
rect 439618 280170 439686 280226
rect 439742 280170 470034 280226
rect 470090 280170 470158 280226
rect 470214 280170 470282 280226
rect 470338 280170 470406 280226
rect 470462 280170 495878 280226
rect 495934 280170 496002 280226
rect 496058 280170 500754 280226
rect 500810 280170 500878 280226
rect 500934 280170 501002 280226
rect 501058 280170 501126 280226
rect 501182 280170 531474 280226
rect 531530 280170 531598 280226
rect 531654 280170 531722 280226
rect 531778 280170 531846 280226
rect 531902 280170 557878 280226
rect 557934 280170 558002 280226
rect 558058 280170 562194 280226
rect 562250 280170 562318 280226
rect 562374 280170 562442 280226
rect 562498 280170 562566 280226
rect 562622 280170 592914 280226
rect 592970 280170 593038 280226
rect 593094 280170 593162 280226
rect 593218 280170 593286 280226
rect 593342 280170 597456 280226
rect 597512 280170 597580 280226
rect 597636 280170 597704 280226
rect 597760 280170 597828 280226
rect 597884 280170 597980 280226
rect -1916 280102 597980 280170
rect -1916 280046 -1820 280102
rect -1764 280046 -1696 280102
rect -1640 280046 -1572 280102
rect -1516 280046 -1448 280102
rect -1392 280046 9234 280102
rect 9290 280046 9358 280102
rect 9414 280046 9482 280102
rect 9538 280046 9606 280102
rect 9662 280046 39878 280102
rect 39934 280046 40002 280102
rect 40058 280046 70674 280102
rect 70730 280046 70798 280102
rect 70854 280046 70922 280102
rect 70978 280046 71046 280102
rect 71102 280046 101878 280102
rect 101934 280046 102002 280102
rect 102058 280046 132114 280102
rect 132170 280046 132238 280102
rect 132294 280046 132362 280102
rect 132418 280046 132486 280102
rect 132542 280046 162834 280102
rect 162890 280046 162958 280102
rect 163014 280046 163082 280102
rect 163138 280046 163206 280102
rect 163262 280046 163878 280102
rect 163934 280046 164002 280102
rect 164058 280046 193554 280102
rect 193610 280046 193678 280102
rect 193734 280046 193802 280102
rect 193858 280046 193926 280102
rect 193982 280046 224274 280102
rect 224330 280046 224398 280102
rect 224454 280046 224522 280102
rect 224578 280046 224646 280102
rect 224702 280046 225878 280102
rect 225934 280046 226002 280102
rect 226058 280046 254994 280102
rect 255050 280046 255118 280102
rect 255174 280046 255242 280102
rect 255298 280046 255366 280102
rect 255422 280046 287878 280102
rect 287934 280046 288002 280102
rect 288058 280046 318598 280102
rect 318654 280046 318722 280102
rect 318778 280046 347154 280102
rect 347210 280046 347278 280102
rect 347334 280046 347402 280102
rect 347458 280046 347526 280102
rect 347582 280046 371878 280102
rect 371934 280046 372002 280102
rect 372058 280046 377874 280102
rect 377930 280046 377998 280102
rect 378054 280046 378122 280102
rect 378178 280046 378246 280102
rect 378302 280046 408594 280102
rect 408650 280046 408718 280102
rect 408774 280046 408842 280102
rect 408898 280046 408966 280102
rect 409022 280046 433878 280102
rect 433934 280046 434002 280102
rect 434058 280046 439314 280102
rect 439370 280046 439438 280102
rect 439494 280046 439562 280102
rect 439618 280046 439686 280102
rect 439742 280046 470034 280102
rect 470090 280046 470158 280102
rect 470214 280046 470282 280102
rect 470338 280046 470406 280102
rect 470462 280046 495878 280102
rect 495934 280046 496002 280102
rect 496058 280046 500754 280102
rect 500810 280046 500878 280102
rect 500934 280046 501002 280102
rect 501058 280046 501126 280102
rect 501182 280046 531474 280102
rect 531530 280046 531598 280102
rect 531654 280046 531722 280102
rect 531778 280046 531846 280102
rect 531902 280046 557878 280102
rect 557934 280046 558002 280102
rect 558058 280046 562194 280102
rect 562250 280046 562318 280102
rect 562374 280046 562442 280102
rect 562498 280046 562566 280102
rect 562622 280046 592914 280102
rect 592970 280046 593038 280102
rect 593094 280046 593162 280102
rect 593218 280046 593286 280102
rect 593342 280046 597456 280102
rect 597512 280046 597580 280102
rect 597636 280046 597704 280102
rect 597760 280046 597828 280102
rect 597884 280046 597980 280102
rect -1916 279978 597980 280046
rect -1916 279922 -1820 279978
rect -1764 279922 -1696 279978
rect -1640 279922 -1572 279978
rect -1516 279922 -1448 279978
rect -1392 279922 9234 279978
rect 9290 279922 9358 279978
rect 9414 279922 9482 279978
rect 9538 279922 9606 279978
rect 9662 279922 39878 279978
rect 39934 279922 40002 279978
rect 40058 279922 70674 279978
rect 70730 279922 70798 279978
rect 70854 279922 70922 279978
rect 70978 279922 71046 279978
rect 71102 279922 101878 279978
rect 101934 279922 102002 279978
rect 102058 279922 132114 279978
rect 132170 279922 132238 279978
rect 132294 279922 132362 279978
rect 132418 279922 132486 279978
rect 132542 279922 162834 279978
rect 162890 279922 162958 279978
rect 163014 279922 163082 279978
rect 163138 279922 163206 279978
rect 163262 279922 163878 279978
rect 163934 279922 164002 279978
rect 164058 279922 193554 279978
rect 193610 279922 193678 279978
rect 193734 279922 193802 279978
rect 193858 279922 193926 279978
rect 193982 279922 224274 279978
rect 224330 279922 224398 279978
rect 224454 279922 224522 279978
rect 224578 279922 224646 279978
rect 224702 279922 225878 279978
rect 225934 279922 226002 279978
rect 226058 279922 254994 279978
rect 255050 279922 255118 279978
rect 255174 279922 255242 279978
rect 255298 279922 255366 279978
rect 255422 279922 287878 279978
rect 287934 279922 288002 279978
rect 288058 279922 318598 279978
rect 318654 279922 318722 279978
rect 318778 279922 347154 279978
rect 347210 279922 347278 279978
rect 347334 279922 347402 279978
rect 347458 279922 347526 279978
rect 347582 279922 371878 279978
rect 371934 279922 372002 279978
rect 372058 279922 377874 279978
rect 377930 279922 377998 279978
rect 378054 279922 378122 279978
rect 378178 279922 378246 279978
rect 378302 279922 408594 279978
rect 408650 279922 408718 279978
rect 408774 279922 408842 279978
rect 408898 279922 408966 279978
rect 409022 279922 433878 279978
rect 433934 279922 434002 279978
rect 434058 279922 439314 279978
rect 439370 279922 439438 279978
rect 439494 279922 439562 279978
rect 439618 279922 439686 279978
rect 439742 279922 470034 279978
rect 470090 279922 470158 279978
rect 470214 279922 470282 279978
rect 470338 279922 470406 279978
rect 470462 279922 495878 279978
rect 495934 279922 496002 279978
rect 496058 279922 500754 279978
rect 500810 279922 500878 279978
rect 500934 279922 501002 279978
rect 501058 279922 501126 279978
rect 501182 279922 531474 279978
rect 531530 279922 531598 279978
rect 531654 279922 531722 279978
rect 531778 279922 531846 279978
rect 531902 279922 557878 279978
rect 557934 279922 558002 279978
rect 558058 279922 562194 279978
rect 562250 279922 562318 279978
rect 562374 279922 562442 279978
rect 562498 279922 562566 279978
rect 562622 279922 592914 279978
rect 592970 279922 593038 279978
rect 593094 279922 593162 279978
rect 593218 279922 593286 279978
rect 593342 279922 597456 279978
rect 597512 279922 597580 279978
rect 597636 279922 597704 279978
rect 597760 279922 597828 279978
rect 597884 279922 597980 279978
rect -1916 279826 597980 279922
rect 195676 278218 263860 278234
rect 195676 278162 195692 278218
rect 195748 278162 263788 278218
rect 263844 278162 263860 278218
rect 195676 278146 263860 278162
rect 126796 278038 263412 278054
rect 126796 277982 126812 278038
rect 126868 277982 263340 278038
rect 263396 277982 263412 278038
rect 126796 277966 263412 277982
rect 334332 278038 455492 278054
rect 334332 277982 334348 278038
rect 334404 277982 455420 278038
rect 455476 277982 455492 278038
rect 334332 277966 455492 277982
rect 334444 277318 396524 277334
rect 334444 277262 334460 277318
rect 334516 277262 396524 277318
rect 334444 277246 396524 277262
rect 396436 277154 396524 277246
rect 396436 277138 455380 277154
rect 396436 277082 455308 277138
rect 455364 277082 455380 277138
rect 396436 277066 455380 277082
rect 127580 276418 262180 276434
rect 127580 276362 127596 276418
rect 127652 276362 262108 276418
rect 262164 276362 262180 276418
rect 127580 276346 262180 276362
rect 64188 275698 124420 275714
rect 64188 275642 64204 275698
rect 64260 275642 124348 275698
rect 124404 275642 124420 275698
rect 64188 275626 124420 275642
rect 133516 275698 263860 275714
rect 133516 275642 133532 275698
rect 133588 275642 263788 275698
rect 263844 275642 263860 275698
rect 133516 275626 263860 275642
rect 334444 275698 394900 275714
rect 334444 275642 334460 275698
rect 334516 275642 394828 275698
rect 394884 275642 394900 275698
rect 334444 275626 394900 275642
rect -1916 274350 597980 274446
rect -1916 274294 -860 274350
rect -804 274294 -736 274350
rect -680 274294 -612 274350
rect -556 274294 -488 274350
rect -432 274294 5514 274350
rect 5570 274294 5638 274350
rect 5694 274294 5762 274350
rect 5818 274294 5886 274350
rect 5942 274294 24518 274350
rect 24574 274294 24642 274350
rect 24698 274294 36234 274350
rect 36290 274294 36358 274350
rect 36414 274294 36482 274350
rect 36538 274294 36606 274350
rect 36662 274294 55238 274350
rect 55294 274294 55362 274350
rect 55418 274294 66954 274350
rect 67010 274294 67078 274350
rect 67134 274294 67202 274350
rect 67258 274294 67326 274350
rect 67382 274294 86518 274350
rect 86574 274294 86642 274350
rect 86698 274294 97674 274350
rect 97730 274294 97798 274350
rect 97854 274294 97922 274350
rect 97978 274294 98046 274350
rect 98102 274294 117238 274350
rect 117294 274294 117362 274350
rect 117418 274294 128394 274350
rect 128450 274294 128518 274350
rect 128574 274294 128642 274350
rect 128698 274294 128766 274350
rect 128822 274294 148518 274350
rect 148574 274294 148642 274350
rect 148698 274294 159114 274350
rect 159170 274294 159238 274350
rect 159294 274294 159362 274350
rect 159418 274294 159486 274350
rect 159542 274294 179238 274350
rect 179294 274294 179362 274350
rect 179418 274294 189834 274350
rect 189890 274294 189958 274350
rect 190014 274294 190082 274350
rect 190138 274294 190206 274350
rect 190262 274294 210518 274350
rect 210574 274294 210642 274350
rect 210698 274294 220554 274350
rect 220610 274294 220678 274350
rect 220734 274294 220802 274350
rect 220858 274294 220926 274350
rect 220982 274294 241238 274350
rect 241294 274294 241362 274350
rect 241418 274294 251274 274350
rect 251330 274294 251398 274350
rect 251454 274294 251522 274350
rect 251578 274294 251646 274350
rect 251702 274294 272518 274350
rect 272574 274294 272642 274350
rect 272698 274294 303238 274350
rect 303294 274294 303362 274350
rect 303418 274294 343434 274350
rect 343490 274294 343558 274350
rect 343614 274294 343682 274350
rect 343738 274294 343806 274350
rect 343862 274294 356518 274350
rect 356574 274294 356642 274350
rect 356698 274294 374154 274350
rect 374210 274294 374278 274350
rect 374334 274294 374402 274350
rect 374458 274294 374526 274350
rect 374582 274294 387238 274350
rect 387294 274294 387362 274350
rect 387418 274294 404874 274350
rect 404930 274294 404998 274350
rect 405054 274294 405122 274350
rect 405178 274294 405246 274350
rect 405302 274294 418518 274350
rect 418574 274294 418642 274350
rect 418698 274294 435594 274350
rect 435650 274294 435718 274350
rect 435774 274294 435842 274350
rect 435898 274294 435966 274350
rect 436022 274294 449238 274350
rect 449294 274294 449362 274350
rect 449418 274294 466314 274350
rect 466370 274294 466438 274350
rect 466494 274294 466562 274350
rect 466618 274294 466686 274350
rect 466742 274294 480518 274350
rect 480574 274294 480642 274350
rect 480698 274294 497034 274350
rect 497090 274294 497158 274350
rect 497214 274294 497282 274350
rect 497338 274294 497406 274350
rect 497462 274294 511238 274350
rect 511294 274294 511362 274350
rect 511418 274294 527754 274350
rect 527810 274294 527878 274350
rect 527934 274294 528002 274350
rect 528058 274294 528126 274350
rect 528182 274294 542518 274350
rect 542574 274294 542642 274350
rect 542698 274294 558474 274350
rect 558530 274294 558598 274350
rect 558654 274294 558722 274350
rect 558778 274294 558846 274350
rect 558902 274294 573238 274350
rect 573294 274294 573362 274350
rect 573418 274294 589194 274350
rect 589250 274294 589318 274350
rect 589374 274294 589442 274350
rect 589498 274294 589566 274350
rect 589622 274294 596496 274350
rect 596552 274294 596620 274350
rect 596676 274294 596744 274350
rect 596800 274294 596868 274350
rect 596924 274294 597980 274350
rect -1916 274226 597980 274294
rect -1916 274170 -860 274226
rect -804 274170 -736 274226
rect -680 274170 -612 274226
rect -556 274170 -488 274226
rect -432 274170 5514 274226
rect 5570 274170 5638 274226
rect 5694 274170 5762 274226
rect 5818 274170 5886 274226
rect 5942 274170 24518 274226
rect 24574 274170 24642 274226
rect 24698 274170 36234 274226
rect 36290 274170 36358 274226
rect 36414 274170 36482 274226
rect 36538 274170 36606 274226
rect 36662 274170 55238 274226
rect 55294 274170 55362 274226
rect 55418 274170 66954 274226
rect 67010 274170 67078 274226
rect 67134 274170 67202 274226
rect 67258 274170 67326 274226
rect 67382 274170 86518 274226
rect 86574 274170 86642 274226
rect 86698 274170 97674 274226
rect 97730 274170 97798 274226
rect 97854 274170 97922 274226
rect 97978 274170 98046 274226
rect 98102 274170 117238 274226
rect 117294 274170 117362 274226
rect 117418 274170 128394 274226
rect 128450 274170 128518 274226
rect 128574 274170 128642 274226
rect 128698 274170 128766 274226
rect 128822 274170 148518 274226
rect 148574 274170 148642 274226
rect 148698 274170 159114 274226
rect 159170 274170 159238 274226
rect 159294 274170 159362 274226
rect 159418 274170 159486 274226
rect 159542 274170 179238 274226
rect 179294 274170 179362 274226
rect 179418 274170 189834 274226
rect 189890 274170 189958 274226
rect 190014 274170 190082 274226
rect 190138 274170 190206 274226
rect 190262 274170 210518 274226
rect 210574 274170 210642 274226
rect 210698 274170 220554 274226
rect 220610 274170 220678 274226
rect 220734 274170 220802 274226
rect 220858 274170 220926 274226
rect 220982 274170 241238 274226
rect 241294 274170 241362 274226
rect 241418 274170 251274 274226
rect 251330 274170 251398 274226
rect 251454 274170 251522 274226
rect 251578 274170 251646 274226
rect 251702 274170 272518 274226
rect 272574 274170 272642 274226
rect 272698 274170 303238 274226
rect 303294 274170 303362 274226
rect 303418 274170 343434 274226
rect 343490 274170 343558 274226
rect 343614 274170 343682 274226
rect 343738 274170 343806 274226
rect 343862 274170 356518 274226
rect 356574 274170 356642 274226
rect 356698 274170 374154 274226
rect 374210 274170 374278 274226
rect 374334 274170 374402 274226
rect 374458 274170 374526 274226
rect 374582 274170 387238 274226
rect 387294 274170 387362 274226
rect 387418 274170 404874 274226
rect 404930 274170 404998 274226
rect 405054 274170 405122 274226
rect 405178 274170 405246 274226
rect 405302 274170 418518 274226
rect 418574 274170 418642 274226
rect 418698 274170 435594 274226
rect 435650 274170 435718 274226
rect 435774 274170 435842 274226
rect 435898 274170 435966 274226
rect 436022 274170 449238 274226
rect 449294 274170 449362 274226
rect 449418 274170 466314 274226
rect 466370 274170 466438 274226
rect 466494 274170 466562 274226
rect 466618 274170 466686 274226
rect 466742 274170 480518 274226
rect 480574 274170 480642 274226
rect 480698 274170 497034 274226
rect 497090 274170 497158 274226
rect 497214 274170 497282 274226
rect 497338 274170 497406 274226
rect 497462 274170 511238 274226
rect 511294 274170 511362 274226
rect 511418 274170 527754 274226
rect 527810 274170 527878 274226
rect 527934 274170 528002 274226
rect 528058 274170 528126 274226
rect 528182 274170 542518 274226
rect 542574 274170 542642 274226
rect 542698 274170 558474 274226
rect 558530 274170 558598 274226
rect 558654 274170 558722 274226
rect 558778 274170 558846 274226
rect 558902 274170 573238 274226
rect 573294 274170 573362 274226
rect 573418 274170 589194 274226
rect 589250 274170 589318 274226
rect 589374 274170 589442 274226
rect 589498 274170 589566 274226
rect 589622 274170 596496 274226
rect 596552 274170 596620 274226
rect 596676 274170 596744 274226
rect 596800 274170 596868 274226
rect 596924 274170 597980 274226
rect -1916 274102 597980 274170
rect -1916 274046 -860 274102
rect -804 274046 -736 274102
rect -680 274046 -612 274102
rect -556 274046 -488 274102
rect -432 274046 5514 274102
rect 5570 274046 5638 274102
rect 5694 274046 5762 274102
rect 5818 274046 5886 274102
rect 5942 274046 24518 274102
rect 24574 274046 24642 274102
rect 24698 274046 36234 274102
rect 36290 274046 36358 274102
rect 36414 274046 36482 274102
rect 36538 274046 36606 274102
rect 36662 274046 55238 274102
rect 55294 274046 55362 274102
rect 55418 274046 66954 274102
rect 67010 274046 67078 274102
rect 67134 274046 67202 274102
rect 67258 274046 67326 274102
rect 67382 274046 86518 274102
rect 86574 274046 86642 274102
rect 86698 274046 97674 274102
rect 97730 274046 97798 274102
rect 97854 274046 97922 274102
rect 97978 274046 98046 274102
rect 98102 274046 117238 274102
rect 117294 274046 117362 274102
rect 117418 274046 128394 274102
rect 128450 274046 128518 274102
rect 128574 274046 128642 274102
rect 128698 274046 128766 274102
rect 128822 274046 148518 274102
rect 148574 274046 148642 274102
rect 148698 274046 159114 274102
rect 159170 274046 159238 274102
rect 159294 274046 159362 274102
rect 159418 274046 159486 274102
rect 159542 274046 179238 274102
rect 179294 274046 179362 274102
rect 179418 274046 189834 274102
rect 189890 274046 189958 274102
rect 190014 274046 190082 274102
rect 190138 274046 190206 274102
rect 190262 274046 210518 274102
rect 210574 274046 210642 274102
rect 210698 274046 220554 274102
rect 220610 274046 220678 274102
rect 220734 274046 220802 274102
rect 220858 274046 220926 274102
rect 220982 274046 241238 274102
rect 241294 274046 241362 274102
rect 241418 274046 251274 274102
rect 251330 274046 251398 274102
rect 251454 274046 251522 274102
rect 251578 274046 251646 274102
rect 251702 274046 272518 274102
rect 272574 274046 272642 274102
rect 272698 274046 303238 274102
rect 303294 274046 303362 274102
rect 303418 274046 343434 274102
rect 343490 274046 343558 274102
rect 343614 274046 343682 274102
rect 343738 274046 343806 274102
rect 343862 274046 356518 274102
rect 356574 274046 356642 274102
rect 356698 274046 374154 274102
rect 374210 274046 374278 274102
rect 374334 274046 374402 274102
rect 374458 274046 374526 274102
rect 374582 274046 387238 274102
rect 387294 274046 387362 274102
rect 387418 274046 404874 274102
rect 404930 274046 404998 274102
rect 405054 274046 405122 274102
rect 405178 274046 405246 274102
rect 405302 274046 418518 274102
rect 418574 274046 418642 274102
rect 418698 274046 435594 274102
rect 435650 274046 435718 274102
rect 435774 274046 435842 274102
rect 435898 274046 435966 274102
rect 436022 274046 449238 274102
rect 449294 274046 449362 274102
rect 449418 274046 466314 274102
rect 466370 274046 466438 274102
rect 466494 274046 466562 274102
rect 466618 274046 466686 274102
rect 466742 274046 480518 274102
rect 480574 274046 480642 274102
rect 480698 274046 497034 274102
rect 497090 274046 497158 274102
rect 497214 274046 497282 274102
rect 497338 274046 497406 274102
rect 497462 274046 511238 274102
rect 511294 274046 511362 274102
rect 511418 274046 527754 274102
rect 527810 274046 527878 274102
rect 527934 274046 528002 274102
rect 528058 274046 528126 274102
rect 528182 274046 542518 274102
rect 542574 274046 542642 274102
rect 542698 274046 558474 274102
rect 558530 274046 558598 274102
rect 558654 274046 558722 274102
rect 558778 274046 558846 274102
rect 558902 274046 573238 274102
rect 573294 274046 573362 274102
rect 573418 274046 589194 274102
rect 589250 274046 589318 274102
rect 589374 274046 589442 274102
rect 589498 274046 589566 274102
rect 589622 274046 596496 274102
rect 596552 274046 596620 274102
rect 596676 274046 596744 274102
rect 596800 274046 596868 274102
rect 596924 274046 597980 274102
rect -1916 273978 597980 274046
rect -1916 273922 -860 273978
rect -804 273922 -736 273978
rect -680 273922 -612 273978
rect -556 273922 -488 273978
rect -432 273922 5514 273978
rect 5570 273922 5638 273978
rect 5694 273922 5762 273978
rect 5818 273922 5886 273978
rect 5942 273922 24518 273978
rect 24574 273922 24642 273978
rect 24698 273922 36234 273978
rect 36290 273922 36358 273978
rect 36414 273922 36482 273978
rect 36538 273922 36606 273978
rect 36662 273922 55238 273978
rect 55294 273922 55362 273978
rect 55418 273922 66954 273978
rect 67010 273922 67078 273978
rect 67134 273922 67202 273978
rect 67258 273922 67326 273978
rect 67382 273922 86518 273978
rect 86574 273922 86642 273978
rect 86698 273922 97674 273978
rect 97730 273922 97798 273978
rect 97854 273922 97922 273978
rect 97978 273922 98046 273978
rect 98102 273922 117238 273978
rect 117294 273922 117362 273978
rect 117418 273922 128394 273978
rect 128450 273922 128518 273978
rect 128574 273922 128642 273978
rect 128698 273922 128766 273978
rect 128822 273922 148518 273978
rect 148574 273922 148642 273978
rect 148698 273922 159114 273978
rect 159170 273922 159238 273978
rect 159294 273922 159362 273978
rect 159418 273922 159486 273978
rect 159542 273922 179238 273978
rect 179294 273922 179362 273978
rect 179418 273922 189834 273978
rect 189890 273922 189958 273978
rect 190014 273922 190082 273978
rect 190138 273922 190206 273978
rect 190262 273922 210518 273978
rect 210574 273922 210642 273978
rect 210698 273922 220554 273978
rect 220610 273922 220678 273978
rect 220734 273922 220802 273978
rect 220858 273922 220926 273978
rect 220982 273922 241238 273978
rect 241294 273922 241362 273978
rect 241418 273922 251274 273978
rect 251330 273922 251398 273978
rect 251454 273922 251522 273978
rect 251578 273922 251646 273978
rect 251702 273922 272518 273978
rect 272574 273922 272642 273978
rect 272698 273922 303238 273978
rect 303294 273922 303362 273978
rect 303418 273922 343434 273978
rect 343490 273922 343558 273978
rect 343614 273922 343682 273978
rect 343738 273922 343806 273978
rect 343862 273922 356518 273978
rect 356574 273922 356642 273978
rect 356698 273922 374154 273978
rect 374210 273922 374278 273978
rect 374334 273922 374402 273978
rect 374458 273922 374526 273978
rect 374582 273922 387238 273978
rect 387294 273922 387362 273978
rect 387418 273922 404874 273978
rect 404930 273922 404998 273978
rect 405054 273922 405122 273978
rect 405178 273922 405246 273978
rect 405302 273922 418518 273978
rect 418574 273922 418642 273978
rect 418698 273922 435594 273978
rect 435650 273922 435718 273978
rect 435774 273922 435842 273978
rect 435898 273922 435966 273978
rect 436022 273922 449238 273978
rect 449294 273922 449362 273978
rect 449418 273922 466314 273978
rect 466370 273922 466438 273978
rect 466494 273922 466562 273978
rect 466618 273922 466686 273978
rect 466742 273922 480518 273978
rect 480574 273922 480642 273978
rect 480698 273922 497034 273978
rect 497090 273922 497158 273978
rect 497214 273922 497282 273978
rect 497338 273922 497406 273978
rect 497462 273922 511238 273978
rect 511294 273922 511362 273978
rect 511418 273922 527754 273978
rect 527810 273922 527878 273978
rect 527934 273922 528002 273978
rect 528058 273922 528126 273978
rect 528182 273922 542518 273978
rect 542574 273922 542642 273978
rect 542698 273922 558474 273978
rect 558530 273922 558598 273978
rect 558654 273922 558722 273978
rect 558778 273922 558846 273978
rect 558902 273922 573238 273978
rect 573294 273922 573362 273978
rect 573418 273922 589194 273978
rect 589250 273922 589318 273978
rect 589374 273922 589442 273978
rect 589498 273922 589566 273978
rect 589622 273922 596496 273978
rect 596552 273922 596620 273978
rect 596676 273922 596744 273978
rect 596800 273922 596868 273978
rect 596924 273922 597980 273978
rect -1916 273826 597980 273922
rect 127580 272998 262292 273014
rect 127580 272942 127596 272998
rect 127652 272942 262220 272998
rect 262276 272942 262292 272998
rect 127580 272926 262292 272942
rect 334444 272998 396692 273014
rect 334444 272942 334460 272998
rect 334516 272942 396620 272998
rect 396676 272942 396692 272998
rect 334444 272926 396692 272942
rect 334332 272278 395684 272294
rect 334332 272222 334348 272278
rect 334404 272222 395612 272278
rect 395668 272222 395684 272278
rect 334332 272206 395684 272222
rect 351020 271738 396916 271754
rect 351020 271682 351036 271738
rect 351092 271682 396844 271738
rect 396900 271682 396916 271738
rect 351020 271666 396916 271682
rect 194892 271558 263860 271574
rect 194892 271502 194908 271558
rect 194964 271502 263788 271558
rect 263844 271502 263860 271558
rect 194892 271486 263860 271502
rect 334444 271558 397028 271574
rect 334444 271502 334460 271558
rect 334516 271502 396956 271558
rect 397012 271502 397028 271558
rect 334444 271486 397028 271502
rect 149476 271378 201700 271394
rect 149476 271322 201628 271378
rect 201684 271322 201700 271378
rect 149476 271306 201700 271322
rect 394812 271378 455604 271394
rect 394812 271322 394828 271378
rect 394884 271322 455604 271378
rect 394812 271306 455604 271322
rect 149476 271214 149564 271306
rect 144044 271198 149564 271214
rect 144044 271142 144060 271198
rect 144116 271142 149564 271198
rect 144044 271126 149564 271142
rect 455516 271018 455604 271306
rect 455516 270962 455532 271018
rect 455588 270962 455604 271018
rect 455516 270946 455604 270962
rect 64636 270838 263972 270854
rect 64636 270782 64652 270838
rect 64708 270782 263900 270838
rect 263956 270782 263972 270838
rect 64636 270766 263972 270782
rect 78916 270658 141108 270674
rect 78916 270602 82460 270658
rect 82516 270602 141036 270658
rect 141092 270602 141108 270658
rect 78916 270586 141108 270602
rect 78916 270494 79004 270586
rect 20060 270478 79004 270494
rect 20060 270422 20076 270478
rect 20132 270422 79004 270478
rect 20060 270406 79004 270422
rect 64188 270298 262180 270314
rect 64188 270242 64204 270298
rect 64260 270242 262108 270298
rect 262164 270242 262180 270298
rect 64188 270226 262180 270242
rect 64188 270118 194980 270134
rect 64188 270062 64204 270118
rect 64260 270062 194908 270118
rect 194964 270062 194980 270118
rect 64188 270046 194980 270062
rect 334556 269758 394900 269774
rect 334556 269702 334572 269758
rect 334628 269702 394828 269758
rect 394884 269702 394900 269758
rect 334556 269686 394900 269702
rect 352700 269578 534340 269594
rect 352700 269522 352716 269578
rect 352772 269522 414652 269578
rect 414708 269522 473676 269578
rect 473732 269522 534268 269578
rect 534324 269522 534340 269578
rect 352700 269506 534340 269522
rect 393804 269038 472180 269054
rect 393804 268982 393820 269038
rect 393876 268982 472108 269038
rect 472164 268982 472180 269038
rect 393804 268966 472180 268982
rect 198252 268858 263860 268874
rect 198252 268802 198268 268858
rect 198324 268802 263788 268858
rect 263844 268802 263860 268858
rect 198252 268786 263860 268802
rect 334444 268858 393556 268874
rect 334444 268802 334460 268858
rect 334516 268802 393484 268858
rect 393540 268802 393556 268858
rect 334444 268786 393556 268802
rect 428300 268858 583060 268874
rect 428300 268802 428316 268858
rect 428372 268802 582988 268858
rect 583044 268802 583060 268858
rect 428300 268786 583060 268802
rect 64188 268678 249524 268694
rect 64188 268622 64204 268678
rect 64260 268622 249452 268678
rect 249508 268622 249524 268678
rect 64188 268606 249524 268622
rect 124332 268498 263860 268514
rect 124332 268442 124348 268498
rect 124404 268442 263788 268498
rect 263844 268442 263860 268498
rect 124332 268426 263860 268442
rect 334444 267958 534340 267974
rect 334444 267902 334460 267958
rect 334516 267902 534268 267958
rect 534324 267902 534340 267958
rect 334444 267886 534340 267902
rect 334332 267418 393332 267434
rect 334332 267362 334348 267418
rect 334404 267362 393260 267418
rect 393316 267362 393332 267418
rect 334332 267346 393332 267362
rect 429196 267418 472180 267434
rect 429196 267362 429212 267418
rect 429268 267362 472108 267418
rect 472164 267362 472180 267418
rect 429196 267346 472180 267362
rect 206428 267238 229364 267254
rect 206428 267182 206444 267238
rect 206500 267182 229364 267238
rect 206428 267166 229364 267182
rect 351916 267238 517540 267254
rect 351916 267182 351932 267238
rect 351988 267182 517468 267238
rect 517524 267182 517540 267238
rect 351916 267166 517540 267182
rect 229276 267074 229364 267166
rect 82444 267058 195764 267074
rect 82444 267002 82460 267058
rect 82516 267002 195692 267058
rect 195748 267002 195764 267058
rect 82444 266986 195764 267002
rect 229276 267058 263860 267074
rect 229276 267002 263788 267058
rect 263844 267002 263860 267058
rect 229276 266986 263860 267002
rect 336908 267058 384764 267074
rect 336908 267002 336924 267058
rect 336980 267002 384764 267058
rect 336908 266986 384764 267002
rect 384676 266714 384764 266986
rect 579276 267058 579364 267074
rect 579276 267002 579292 267058
rect 579348 267002 579364 267058
rect 384676 266698 393444 266714
rect 384676 266642 393372 266698
rect 393428 266642 393444 266698
rect 384676 266626 393444 266642
rect 393580 266698 579140 266714
rect 393580 266642 393596 266698
rect 393652 266642 579068 266698
rect 579124 266642 579140 266698
rect 393580 266626 579140 266642
rect 579276 266534 579364 267002
rect 206316 266518 263860 266534
rect 206316 266462 206332 266518
rect 206388 266462 263788 266518
rect 263844 266462 263860 266518
rect 206316 266446 263860 266462
rect 334444 266518 579364 266534
rect 334444 266462 334460 266518
rect 334516 266462 579364 266518
rect 334444 266446 579364 266462
rect 334556 266338 429284 266354
rect 334556 266282 334572 266338
rect 334628 266282 429212 266338
rect 429268 266282 429284 266338
rect 334556 266266 429284 266282
rect 334444 265438 428388 265454
rect 334444 265382 334460 265438
rect 334516 265382 428316 265438
rect 428372 265382 428388 265438
rect 334444 265366 428388 265382
rect 347772 265258 393444 265274
rect 347772 265202 347788 265258
rect 347844 265202 393444 265258
rect 347772 265186 393444 265202
rect 189516 264898 262628 264914
rect 189516 264842 189532 264898
rect 189588 264842 262556 264898
rect 262612 264842 262628 264898
rect 189516 264826 262628 264842
rect 393356 264898 393444 265186
rect 393356 264842 393372 264898
rect 393428 264842 393444 264898
rect 393356 264826 393444 264842
rect 141020 264718 260052 264734
rect 141020 264662 141036 264718
rect 141092 264662 259980 264718
rect 260036 264662 260052 264718
rect 141020 264646 260052 264662
rect 64188 264538 198340 264554
rect 64188 264482 64204 264538
rect 64260 264482 198268 264538
rect 198324 264482 198340 264538
rect 64188 264466 198340 264482
rect 334444 263818 428500 263834
rect 334444 263762 334460 263818
rect 334516 263762 428428 263818
rect 428484 263762 428500 263818
rect 334444 263746 428500 263762
rect 334444 263638 393668 263654
rect 334444 263582 334460 263638
rect 334516 263582 393596 263638
rect 393652 263582 393668 263638
rect 334444 263566 393668 263582
rect -1916 262350 597980 262446
rect -1916 262294 -1820 262350
rect -1764 262294 -1696 262350
rect -1640 262294 -1572 262350
rect -1516 262294 -1448 262350
rect -1392 262294 9234 262350
rect 9290 262294 9358 262350
rect 9414 262294 9482 262350
rect 9538 262294 9606 262350
rect 9662 262294 39878 262350
rect 39934 262294 40002 262350
rect 40058 262294 70674 262350
rect 70730 262294 70798 262350
rect 70854 262294 70922 262350
rect 70978 262294 71046 262350
rect 71102 262294 101878 262350
rect 101934 262294 102002 262350
rect 102058 262294 132114 262350
rect 132170 262294 132238 262350
rect 132294 262294 132362 262350
rect 132418 262294 132486 262350
rect 132542 262294 163878 262350
rect 163934 262294 164002 262350
rect 164058 262294 193554 262350
rect 193610 262294 193678 262350
rect 193734 262294 193802 262350
rect 193858 262294 193926 262350
rect 193982 262294 224274 262350
rect 224330 262294 224398 262350
rect 224454 262294 224522 262350
rect 224578 262294 224646 262350
rect 224702 262294 225878 262350
rect 225934 262294 226002 262350
rect 226058 262294 254994 262350
rect 255050 262294 255118 262350
rect 255174 262294 255242 262350
rect 255298 262294 255366 262350
rect 255422 262294 287878 262350
rect 287934 262294 288002 262350
rect 288058 262294 318598 262350
rect 318654 262294 318722 262350
rect 318778 262294 347154 262350
rect 347210 262294 347278 262350
rect 347334 262294 347402 262350
rect 347458 262294 347526 262350
rect 347582 262294 371878 262350
rect 371934 262294 372002 262350
rect 372058 262294 377874 262350
rect 377930 262294 377998 262350
rect 378054 262294 378122 262350
rect 378178 262294 378246 262350
rect 378302 262294 408594 262350
rect 408650 262294 408718 262350
rect 408774 262294 408842 262350
rect 408898 262294 408966 262350
rect 409022 262294 433878 262350
rect 433934 262294 434002 262350
rect 434058 262294 439314 262350
rect 439370 262294 439438 262350
rect 439494 262294 439562 262350
rect 439618 262294 439686 262350
rect 439742 262294 470034 262350
rect 470090 262294 470158 262350
rect 470214 262294 470282 262350
rect 470338 262294 470406 262350
rect 470462 262294 495878 262350
rect 495934 262294 496002 262350
rect 496058 262294 500754 262350
rect 500810 262294 500878 262350
rect 500934 262294 501002 262350
rect 501058 262294 501126 262350
rect 501182 262294 531474 262350
rect 531530 262294 531598 262350
rect 531654 262294 531722 262350
rect 531778 262294 531846 262350
rect 531902 262294 557878 262350
rect 557934 262294 558002 262350
rect 558058 262294 562194 262350
rect 562250 262294 562318 262350
rect 562374 262294 562442 262350
rect 562498 262294 562566 262350
rect 562622 262294 592914 262350
rect 592970 262294 593038 262350
rect 593094 262294 593162 262350
rect 593218 262294 593286 262350
rect 593342 262294 597456 262350
rect 597512 262294 597580 262350
rect 597636 262294 597704 262350
rect 597760 262294 597828 262350
rect 597884 262294 597980 262350
rect -1916 262226 597980 262294
rect -1916 262170 -1820 262226
rect -1764 262170 -1696 262226
rect -1640 262170 -1572 262226
rect -1516 262170 -1448 262226
rect -1392 262170 9234 262226
rect 9290 262170 9358 262226
rect 9414 262170 9482 262226
rect 9538 262170 9606 262226
rect 9662 262170 39878 262226
rect 39934 262170 40002 262226
rect 40058 262170 70674 262226
rect 70730 262170 70798 262226
rect 70854 262170 70922 262226
rect 70978 262170 71046 262226
rect 71102 262170 101878 262226
rect 101934 262170 102002 262226
rect 102058 262170 132114 262226
rect 132170 262170 132238 262226
rect 132294 262170 132362 262226
rect 132418 262170 132486 262226
rect 132542 262170 163878 262226
rect 163934 262170 164002 262226
rect 164058 262170 193554 262226
rect 193610 262170 193678 262226
rect 193734 262170 193802 262226
rect 193858 262170 193926 262226
rect 193982 262170 224274 262226
rect 224330 262170 224398 262226
rect 224454 262170 224522 262226
rect 224578 262170 224646 262226
rect 224702 262170 225878 262226
rect 225934 262170 226002 262226
rect 226058 262170 254994 262226
rect 255050 262170 255118 262226
rect 255174 262170 255242 262226
rect 255298 262170 255366 262226
rect 255422 262170 287878 262226
rect 287934 262170 288002 262226
rect 288058 262170 318598 262226
rect 318654 262170 318722 262226
rect 318778 262170 347154 262226
rect 347210 262170 347278 262226
rect 347334 262170 347402 262226
rect 347458 262170 347526 262226
rect 347582 262170 371878 262226
rect 371934 262170 372002 262226
rect 372058 262170 377874 262226
rect 377930 262170 377998 262226
rect 378054 262170 378122 262226
rect 378178 262170 378246 262226
rect 378302 262170 408594 262226
rect 408650 262170 408718 262226
rect 408774 262170 408842 262226
rect 408898 262170 408966 262226
rect 409022 262170 433878 262226
rect 433934 262170 434002 262226
rect 434058 262170 439314 262226
rect 439370 262170 439438 262226
rect 439494 262170 439562 262226
rect 439618 262170 439686 262226
rect 439742 262170 470034 262226
rect 470090 262170 470158 262226
rect 470214 262170 470282 262226
rect 470338 262170 470406 262226
rect 470462 262170 495878 262226
rect 495934 262170 496002 262226
rect 496058 262170 500754 262226
rect 500810 262170 500878 262226
rect 500934 262170 501002 262226
rect 501058 262170 501126 262226
rect 501182 262170 531474 262226
rect 531530 262170 531598 262226
rect 531654 262170 531722 262226
rect 531778 262170 531846 262226
rect 531902 262170 557878 262226
rect 557934 262170 558002 262226
rect 558058 262170 562194 262226
rect 562250 262170 562318 262226
rect 562374 262170 562442 262226
rect 562498 262170 562566 262226
rect 562622 262170 592914 262226
rect 592970 262170 593038 262226
rect 593094 262170 593162 262226
rect 593218 262170 593286 262226
rect 593342 262170 597456 262226
rect 597512 262170 597580 262226
rect 597636 262170 597704 262226
rect 597760 262170 597828 262226
rect 597884 262170 597980 262226
rect -1916 262102 597980 262170
rect -1916 262046 -1820 262102
rect -1764 262046 -1696 262102
rect -1640 262046 -1572 262102
rect -1516 262046 -1448 262102
rect -1392 262046 9234 262102
rect 9290 262046 9358 262102
rect 9414 262046 9482 262102
rect 9538 262046 9606 262102
rect 9662 262046 39878 262102
rect 39934 262046 40002 262102
rect 40058 262046 70674 262102
rect 70730 262046 70798 262102
rect 70854 262046 70922 262102
rect 70978 262046 71046 262102
rect 71102 262046 101878 262102
rect 101934 262046 102002 262102
rect 102058 262046 132114 262102
rect 132170 262046 132238 262102
rect 132294 262046 132362 262102
rect 132418 262046 132486 262102
rect 132542 262052 163878 262102
rect 132542 262046 162834 262052
rect -1916 261996 162834 262046
rect 162890 261996 162958 262052
rect 163014 261996 163082 262052
rect 163138 261996 163206 262052
rect 163262 262046 163878 262052
rect 163934 262046 164002 262102
rect 164058 262046 193554 262102
rect 193610 262046 193678 262102
rect 193734 262046 193802 262102
rect 193858 262046 193926 262102
rect 193982 262046 224274 262102
rect 224330 262046 224398 262102
rect 224454 262046 224522 262102
rect 224578 262046 224646 262102
rect 224702 262046 225878 262102
rect 225934 262046 226002 262102
rect 226058 262046 254994 262102
rect 255050 262046 255118 262102
rect 255174 262046 255242 262102
rect 255298 262046 255366 262102
rect 255422 262046 287878 262102
rect 287934 262046 288002 262102
rect 288058 262046 318598 262102
rect 318654 262046 318722 262102
rect 318778 262046 347154 262102
rect 347210 262046 347278 262102
rect 347334 262046 347402 262102
rect 347458 262046 347526 262102
rect 347582 262046 371878 262102
rect 371934 262046 372002 262102
rect 372058 262046 377874 262102
rect 377930 262046 377998 262102
rect 378054 262046 378122 262102
rect 378178 262046 378246 262102
rect 378302 262046 408594 262102
rect 408650 262046 408718 262102
rect 408774 262046 408842 262102
rect 408898 262046 408966 262102
rect 409022 262046 433878 262102
rect 433934 262046 434002 262102
rect 434058 262046 439314 262102
rect 439370 262046 439438 262102
rect 439494 262046 439562 262102
rect 439618 262046 439686 262102
rect 439742 262046 470034 262102
rect 470090 262046 470158 262102
rect 470214 262046 470282 262102
rect 470338 262046 470406 262102
rect 470462 262046 495878 262102
rect 495934 262046 496002 262102
rect 496058 262046 500754 262102
rect 500810 262046 500878 262102
rect 500934 262046 501002 262102
rect 501058 262046 501126 262102
rect 501182 262046 531474 262102
rect 531530 262046 531598 262102
rect 531654 262046 531722 262102
rect 531778 262046 531846 262102
rect 531902 262046 557878 262102
rect 557934 262046 558002 262102
rect 558058 262046 562194 262102
rect 562250 262046 562318 262102
rect 562374 262046 562442 262102
rect 562498 262046 562566 262102
rect 562622 262046 592914 262102
rect 592970 262046 593038 262102
rect 593094 262046 593162 262102
rect 593218 262046 593286 262102
rect 593342 262046 597456 262102
rect 597512 262046 597580 262102
rect 597636 262046 597704 262102
rect 597760 262046 597828 262102
rect 597884 262046 597980 262102
rect 163262 261996 597980 262046
rect -1916 261978 597980 261996
rect -1916 261922 -1820 261978
rect -1764 261922 -1696 261978
rect -1640 261922 -1572 261978
rect -1516 261922 -1448 261978
rect -1392 261922 9234 261978
rect 9290 261922 9358 261978
rect 9414 261922 9482 261978
rect 9538 261922 9606 261978
rect 9662 261922 39878 261978
rect 39934 261922 40002 261978
rect 40058 261922 70674 261978
rect 70730 261922 70798 261978
rect 70854 261922 70922 261978
rect 70978 261922 71046 261978
rect 71102 261922 101878 261978
rect 101934 261922 102002 261978
rect 102058 261922 132114 261978
rect 132170 261922 132238 261978
rect 132294 261922 132362 261978
rect 132418 261922 132486 261978
rect 132542 261928 163878 261978
rect 132542 261922 162834 261928
rect -1916 261872 162834 261922
rect 162890 261872 162958 261928
rect 163014 261872 163082 261928
rect 163138 261872 163206 261928
rect 163262 261922 163878 261928
rect 163934 261922 164002 261978
rect 164058 261922 193554 261978
rect 193610 261922 193678 261978
rect 193734 261922 193802 261978
rect 193858 261922 193926 261978
rect 193982 261922 224274 261978
rect 224330 261922 224398 261978
rect 224454 261922 224522 261978
rect 224578 261922 224646 261978
rect 224702 261922 225878 261978
rect 225934 261922 226002 261978
rect 226058 261922 254994 261978
rect 255050 261922 255118 261978
rect 255174 261922 255242 261978
rect 255298 261922 255366 261978
rect 255422 261922 287878 261978
rect 287934 261922 288002 261978
rect 288058 261922 318598 261978
rect 318654 261922 318722 261978
rect 318778 261922 347154 261978
rect 347210 261922 347278 261978
rect 347334 261922 347402 261978
rect 347458 261922 347526 261978
rect 347582 261922 371878 261978
rect 371934 261922 372002 261978
rect 372058 261922 377874 261978
rect 377930 261922 377998 261978
rect 378054 261922 378122 261978
rect 378178 261922 378246 261978
rect 378302 261922 408594 261978
rect 408650 261922 408718 261978
rect 408774 261922 408842 261978
rect 408898 261922 408966 261978
rect 409022 261922 433878 261978
rect 433934 261922 434002 261978
rect 434058 261922 439314 261978
rect 439370 261922 439438 261978
rect 439494 261922 439562 261978
rect 439618 261922 439686 261978
rect 439742 261922 470034 261978
rect 470090 261922 470158 261978
rect 470214 261922 470282 261978
rect 470338 261922 470406 261978
rect 470462 261922 495878 261978
rect 495934 261922 496002 261978
rect 496058 261922 500754 261978
rect 500810 261922 500878 261978
rect 500934 261922 501002 261978
rect 501058 261922 501126 261978
rect 501182 261922 531474 261978
rect 531530 261922 531598 261978
rect 531654 261922 531722 261978
rect 531778 261922 531846 261978
rect 531902 261922 557878 261978
rect 557934 261922 558002 261978
rect 558058 261922 562194 261978
rect 562250 261922 562318 261978
rect 562374 261922 562442 261978
rect 562498 261922 562566 261978
rect 562622 261922 592914 261978
rect 592970 261922 593038 261978
rect 593094 261922 593162 261978
rect 593218 261922 593286 261978
rect 593342 261922 597456 261978
rect 597512 261922 597580 261978
rect 597636 261922 597704 261978
rect 597760 261922 597828 261978
rect 597884 261922 597980 261978
rect 163262 261872 597980 261922
rect -1916 261826 597980 261872
rect 206428 261658 260388 261674
rect 206428 261602 206444 261658
rect 206500 261602 260316 261658
rect 260372 261602 260388 261658
rect 206428 261586 260388 261602
rect 572836 260938 579364 260954
rect 572836 260882 579292 260938
rect 579348 260882 579364 260938
rect 572836 260866 579364 260882
rect 572836 260774 572924 260866
rect 334444 260758 572924 260774
rect 334444 260702 334460 260758
rect 334516 260702 572924 260758
rect 334444 260686 572924 260702
rect 334444 260578 396524 260594
rect 334444 260522 334460 260578
rect 334516 260522 396524 260578
rect 334444 260506 396524 260522
rect 144268 260398 263860 260414
rect 144268 260342 144284 260398
rect 144340 260342 263788 260398
rect 263844 260342 263860 260398
rect 144268 260326 263860 260342
rect 334444 260398 393892 260414
rect 334444 260342 334460 260398
rect 334516 260342 393820 260398
rect 393876 260342 393892 260398
rect 334444 260326 393892 260342
rect 396436 260234 396524 260506
rect 428412 260398 579700 260414
rect 428412 260342 428428 260398
rect 428484 260342 579628 260398
rect 579684 260342 579700 260398
rect 428412 260326 579700 260342
rect 199820 260218 263972 260234
rect 199820 260162 199836 260218
rect 199892 260162 263900 260218
rect 263956 260162 263972 260218
rect 199820 260146 263972 260162
rect 396436 260218 534340 260234
rect 396436 260162 534268 260218
rect 534324 260162 534340 260218
rect 396436 260146 534340 260162
rect 82668 259498 125204 259514
rect 82668 259442 82684 259498
rect 82740 259442 125132 259498
rect 125188 259442 125204 259498
rect 82668 259426 125204 259442
rect 334444 258958 393220 258974
rect 334444 258902 334460 258958
rect 334516 258902 393148 258958
rect 393204 258902 393220 258958
rect 334444 258886 393220 258902
rect 351020 258778 472180 258794
rect 351020 258722 351036 258778
rect 351092 258722 472108 258778
rect 472164 258722 472180 258778
rect 351020 258706 472180 258722
rect 142700 258598 263860 258614
rect 142700 258542 142716 258598
rect 142772 258542 263788 258598
rect 263844 258542 263860 258598
rect 142700 258526 263860 258542
rect 334444 258598 468708 258614
rect 334444 258542 334460 258598
rect 334516 258542 468636 258598
rect 468692 258542 468708 258598
rect 334444 258526 468708 258542
rect 194892 258418 263972 258434
rect 194892 258362 194908 258418
rect 194964 258362 263900 258418
rect 263956 258362 263972 258418
rect 194892 258346 263972 258362
rect 393132 258418 502364 258434
rect 393132 258362 393148 258418
rect 393204 258362 502364 258418
rect 393132 258346 502364 258362
rect 502276 258254 502364 258346
rect 334444 258238 456948 258254
rect 334444 258182 334460 258238
rect 334516 258182 456876 258238
rect 456932 258182 456948 258238
rect 334444 258166 456948 258182
rect 502276 258238 517540 258254
rect 502276 258182 517468 258238
rect 517524 258182 517540 258238
rect 502276 258166 517540 258182
rect -1916 256350 597980 256446
rect -1916 256294 -860 256350
rect -804 256294 -736 256350
rect -680 256294 -612 256350
rect -556 256294 -488 256350
rect -432 256294 5514 256350
rect 5570 256294 5638 256350
rect 5694 256294 5762 256350
rect 5818 256294 5886 256350
rect 5942 256294 24518 256350
rect 24574 256294 24642 256350
rect 24698 256294 36234 256350
rect 36290 256294 36358 256350
rect 36414 256294 36482 256350
rect 36538 256294 36606 256350
rect 36662 256294 55238 256350
rect 55294 256294 55362 256350
rect 55418 256294 66954 256350
rect 67010 256294 67078 256350
rect 67134 256294 67202 256350
rect 67258 256294 67326 256350
rect 67382 256294 86518 256350
rect 86574 256294 86642 256350
rect 86698 256294 97674 256350
rect 97730 256294 97798 256350
rect 97854 256294 97922 256350
rect 97978 256294 98046 256350
rect 98102 256294 117238 256350
rect 117294 256294 117362 256350
rect 117418 256294 128394 256350
rect 128450 256294 128518 256350
rect 128574 256294 128642 256350
rect 128698 256294 128766 256350
rect 128822 256294 148518 256350
rect 148574 256294 148642 256350
rect 148698 256294 159114 256350
rect 159170 256294 159238 256350
rect 159294 256294 159362 256350
rect 159418 256294 159486 256350
rect 159542 256294 179238 256350
rect 179294 256294 179362 256350
rect 179418 256294 189834 256350
rect 189890 256294 189958 256350
rect 190014 256294 190082 256350
rect 190138 256294 190206 256350
rect 190262 256294 210518 256350
rect 210574 256294 210642 256350
rect 210698 256294 220554 256350
rect 220610 256294 220678 256350
rect 220734 256294 220802 256350
rect 220858 256294 220926 256350
rect 220982 256294 241238 256350
rect 241294 256294 241362 256350
rect 241418 256294 251274 256350
rect 251330 256294 251398 256350
rect 251454 256294 251522 256350
rect 251578 256294 251646 256350
rect 251702 256294 272518 256350
rect 272574 256294 272642 256350
rect 272698 256294 303238 256350
rect 303294 256294 303362 256350
rect 303418 256294 343434 256350
rect 343490 256294 343558 256350
rect 343614 256294 343682 256350
rect 343738 256294 343806 256350
rect 343862 256294 356518 256350
rect 356574 256294 356642 256350
rect 356698 256294 374154 256350
rect 374210 256294 374278 256350
rect 374334 256294 374402 256350
rect 374458 256294 374526 256350
rect 374582 256294 387238 256350
rect 387294 256294 387362 256350
rect 387418 256294 404874 256350
rect 404930 256294 404998 256350
rect 405054 256294 405122 256350
rect 405178 256294 405246 256350
rect 405302 256294 418518 256350
rect 418574 256294 418642 256350
rect 418698 256294 435594 256350
rect 435650 256294 435718 256350
rect 435774 256294 435842 256350
rect 435898 256294 435966 256350
rect 436022 256294 449238 256350
rect 449294 256294 449362 256350
rect 449418 256294 466314 256350
rect 466370 256294 466438 256350
rect 466494 256294 466562 256350
rect 466618 256294 466686 256350
rect 466742 256294 480518 256350
rect 480574 256294 480642 256350
rect 480698 256294 497034 256350
rect 497090 256294 497158 256350
rect 497214 256294 497282 256350
rect 497338 256294 497406 256350
rect 497462 256294 511238 256350
rect 511294 256294 511362 256350
rect 511418 256294 527754 256350
rect 527810 256294 527878 256350
rect 527934 256294 528002 256350
rect 528058 256294 528126 256350
rect 528182 256294 542518 256350
rect 542574 256294 542642 256350
rect 542698 256294 558474 256350
rect 558530 256294 558598 256350
rect 558654 256294 558722 256350
rect 558778 256294 558846 256350
rect 558902 256294 573238 256350
rect 573294 256294 573362 256350
rect 573418 256294 589194 256350
rect 589250 256294 589318 256350
rect 589374 256294 589442 256350
rect 589498 256294 589566 256350
rect 589622 256294 596496 256350
rect 596552 256294 596620 256350
rect 596676 256294 596744 256350
rect 596800 256294 596868 256350
rect 596924 256294 597980 256350
rect -1916 256226 597980 256294
rect -1916 256170 -860 256226
rect -804 256170 -736 256226
rect -680 256170 -612 256226
rect -556 256170 -488 256226
rect -432 256170 5514 256226
rect 5570 256170 5638 256226
rect 5694 256170 5762 256226
rect 5818 256170 5886 256226
rect 5942 256170 24518 256226
rect 24574 256170 24642 256226
rect 24698 256170 36234 256226
rect 36290 256170 36358 256226
rect 36414 256170 36482 256226
rect 36538 256170 36606 256226
rect 36662 256170 55238 256226
rect 55294 256170 55362 256226
rect 55418 256170 66954 256226
rect 67010 256170 67078 256226
rect 67134 256170 67202 256226
rect 67258 256170 67326 256226
rect 67382 256170 86518 256226
rect 86574 256170 86642 256226
rect 86698 256170 97674 256226
rect 97730 256170 97798 256226
rect 97854 256170 97922 256226
rect 97978 256170 98046 256226
rect 98102 256170 117238 256226
rect 117294 256170 117362 256226
rect 117418 256170 128394 256226
rect 128450 256170 128518 256226
rect 128574 256170 128642 256226
rect 128698 256170 128766 256226
rect 128822 256170 148518 256226
rect 148574 256170 148642 256226
rect 148698 256170 159114 256226
rect 159170 256170 159238 256226
rect 159294 256170 159362 256226
rect 159418 256170 159486 256226
rect 159542 256170 179238 256226
rect 179294 256170 179362 256226
rect 179418 256170 189834 256226
rect 189890 256170 189958 256226
rect 190014 256170 190082 256226
rect 190138 256170 190206 256226
rect 190262 256170 210518 256226
rect 210574 256170 210642 256226
rect 210698 256170 220554 256226
rect 220610 256170 220678 256226
rect 220734 256170 220802 256226
rect 220858 256170 220926 256226
rect 220982 256170 241238 256226
rect 241294 256170 241362 256226
rect 241418 256170 251274 256226
rect 251330 256170 251398 256226
rect 251454 256170 251522 256226
rect 251578 256170 251646 256226
rect 251702 256170 272518 256226
rect 272574 256170 272642 256226
rect 272698 256170 303238 256226
rect 303294 256170 303362 256226
rect 303418 256170 343434 256226
rect 343490 256170 343558 256226
rect 343614 256170 343682 256226
rect 343738 256170 343806 256226
rect 343862 256170 356518 256226
rect 356574 256170 356642 256226
rect 356698 256170 374154 256226
rect 374210 256170 374278 256226
rect 374334 256170 374402 256226
rect 374458 256170 374526 256226
rect 374582 256170 387238 256226
rect 387294 256170 387362 256226
rect 387418 256170 404874 256226
rect 404930 256170 404998 256226
rect 405054 256170 405122 256226
rect 405178 256170 405246 256226
rect 405302 256170 418518 256226
rect 418574 256170 418642 256226
rect 418698 256170 435594 256226
rect 435650 256170 435718 256226
rect 435774 256170 435842 256226
rect 435898 256170 435966 256226
rect 436022 256170 449238 256226
rect 449294 256170 449362 256226
rect 449418 256170 466314 256226
rect 466370 256170 466438 256226
rect 466494 256170 466562 256226
rect 466618 256170 466686 256226
rect 466742 256170 480518 256226
rect 480574 256170 480642 256226
rect 480698 256170 497034 256226
rect 497090 256170 497158 256226
rect 497214 256170 497282 256226
rect 497338 256170 497406 256226
rect 497462 256170 511238 256226
rect 511294 256170 511362 256226
rect 511418 256170 527754 256226
rect 527810 256170 527878 256226
rect 527934 256170 528002 256226
rect 528058 256170 528126 256226
rect 528182 256170 542518 256226
rect 542574 256170 542642 256226
rect 542698 256170 558474 256226
rect 558530 256170 558598 256226
rect 558654 256170 558722 256226
rect 558778 256170 558846 256226
rect 558902 256170 573238 256226
rect 573294 256170 573362 256226
rect 573418 256170 589194 256226
rect 589250 256170 589318 256226
rect 589374 256170 589442 256226
rect 589498 256170 589566 256226
rect 589622 256170 596496 256226
rect 596552 256170 596620 256226
rect 596676 256170 596744 256226
rect 596800 256170 596868 256226
rect 596924 256170 597980 256226
rect -1916 256102 597980 256170
rect -1916 256046 -860 256102
rect -804 256046 -736 256102
rect -680 256046 -612 256102
rect -556 256046 -488 256102
rect -432 256046 5514 256102
rect 5570 256046 5638 256102
rect 5694 256046 5762 256102
rect 5818 256046 5886 256102
rect 5942 256046 24518 256102
rect 24574 256046 24642 256102
rect 24698 256046 36234 256102
rect 36290 256046 36358 256102
rect 36414 256046 36482 256102
rect 36538 256046 36606 256102
rect 36662 256046 55238 256102
rect 55294 256046 55362 256102
rect 55418 256046 66954 256102
rect 67010 256046 67078 256102
rect 67134 256046 67202 256102
rect 67258 256046 67326 256102
rect 67382 256046 86518 256102
rect 86574 256046 86642 256102
rect 86698 256046 97674 256102
rect 97730 256046 97798 256102
rect 97854 256046 97922 256102
rect 97978 256046 98046 256102
rect 98102 256046 117238 256102
rect 117294 256046 117362 256102
rect 117418 256046 128394 256102
rect 128450 256046 128518 256102
rect 128574 256046 128642 256102
rect 128698 256046 128766 256102
rect 128822 256046 148518 256102
rect 148574 256046 148642 256102
rect 148698 256046 159114 256102
rect 159170 256046 159238 256102
rect 159294 256046 159362 256102
rect 159418 256046 159486 256102
rect 159542 256046 179238 256102
rect 179294 256046 179362 256102
rect 179418 256046 189834 256102
rect 189890 256046 189958 256102
rect 190014 256046 190082 256102
rect 190138 256046 190206 256102
rect 190262 256046 210518 256102
rect 210574 256046 210642 256102
rect 210698 256046 220554 256102
rect 220610 256046 220678 256102
rect 220734 256046 220802 256102
rect 220858 256046 220926 256102
rect 220982 256046 241238 256102
rect 241294 256046 241362 256102
rect 241418 256046 251274 256102
rect 251330 256046 251398 256102
rect 251454 256046 251522 256102
rect 251578 256046 251646 256102
rect 251702 256046 272518 256102
rect 272574 256046 272642 256102
rect 272698 256046 303238 256102
rect 303294 256046 303362 256102
rect 303418 256046 343434 256102
rect 343490 256046 343558 256102
rect 343614 256046 343682 256102
rect 343738 256046 343806 256102
rect 343862 256046 356518 256102
rect 356574 256046 356642 256102
rect 356698 256046 374154 256102
rect 374210 256046 374278 256102
rect 374334 256046 374402 256102
rect 374458 256046 374526 256102
rect 374582 256046 387238 256102
rect 387294 256046 387362 256102
rect 387418 256046 404874 256102
rect 404930 256046 404998 256102
rect 405054 256046 405122 256102
rect 405178 256046 405246 256102
rect 405302 256046 418518 256102
rect 418574 256046 418642 256102
rect 418698 256046 435594 256102
rect 435650 256046 435718 256102
rect 435774 256046 435842 256102
rect 435898 256046 435966 256102
rect 436022 256046 449238 256102
rect 449294 256046 449362 256102
rect 449418 256046 466314 256102
rect 466370 256046 466438 256102
rect 466494 256046 466562 256102
rect 466618 256046 466686 256102
rect 466742 256046 480518 256102
rect 480574 256046 480642 256102
rect 480698 256046 497034 256102
rect 497090 256046 497158 256102
rect 497214 256046 497282 256102
rect 497338 256046 497406 256102
rect 497462 256046 511238 256102
rect 511294 256046 511362 256102
rect 511418 256046 527754 256102
rect 527810 256046 527878 256102
rect 527934 256046 528002 256102
rect 528058 256046 528126 256102
rect 528182 256046 542518 256102
rect 542574 256046 542642 256102
rect 542698 256046 558474 256102
rect 558530 256046 558598 256102
rect 558654 256046 558722 256102
rect 558778 256046 558846 256102
rect 558902 256046 573238 256102
rect 573294 256046 573362 256102
rect 573418 256046 589194 256102
rect 589250 256046 589318 256102
rect 589374 256046 589442 256102
rect 589498 256046 589566 256102
rect 589622 256046 596496 256102
rect 596552 256046 596620 256102
rect 596676 256046 596744 256102
rect 596800 256046 596868 256102
rect 596924 256046 597980 256102
rect -1916 255978 597980 256046
rect -1916 255922 -860 255978
rect -804 255922 -736 255978
rect -680 255922 -612 255978
rect -556 255922 -488 255978
rect -432 255922 5514 255978
rect 5570 255922 5638 255978
rect 5694 255922 5762 255978
rect 5818 255922 5886 255978
rect 5942 255922 24518 255978
rect 24574 255922 24642 255978
rect 24698 255922 36234 255978
rect 36290 255922 36358 255978
rect 36414 255922 36482 255978
rect 36538 255922 36606 255978
rect 36662 255922 55238 255978
rect 55294 255922 55362 255978
rect 55418 255922 66954 255978
rect 67010 255922 67078 255978
rect 67134 255922 67202 255978
rect 67258 255922 67326 255978
rect 67382 255922 86518 255978
rect 86574 255922 86642 255978
rect 86698 255922 97674 255978
rect 97730 255922 97798 255978
rect 97854 255922 97922 255978
rect 97978 255922 98046 255978
rect 98102 255922 117238 255978
rect 117294 255922 117362 255978
rect 117418 255922 128394 255978
rect 128450 255922 128518 255978
rect 128574 255922 128642 255978
rect 128698 255922 128766 255978
rect 128822 255922 148518 255978
rect 148574 255922 148642 255978
rect 148698 255922 159114 255978
rect 159170 255922 159238 255978
rect 159294 255922 159362 255978
rect 159418 255922 159486 255978
rect 159542 255922 179238 255978
rect 179294 255922 179362 255978
rect 179418 255922 189834 255978
rect 189890 255922 189958 255978
rect 190014 255922 190082 255978
rect 190138 255922 190206 255978
rect 190262 255922 210518 255978
rect 210574 255922 210642 255978
rect 210698 255922 220554 255978
rect 220610 255922 220678 255978
rect 220734 255922 220802 255978
rect 220858 255922 220926 255978
rect 220982 255922 241238 255978
rect 241294 255922 241362 255978
rect 241418 255922 251274 255978
rect 251330 255922 251398 255978
rect 251454 255922 251522 255978
rect 251578 255922 251646 255978
rect 251702 255922 272518 255978
rect 272574 255922 272642 255978
rect 272698 255922 303238 255978
rect 303294 255922 303362 255978
rect 303418 255922 343434 255978
rect 343490 255922 343558 255978
rect 343614 255922 343682 255978
rect 343738 255922 343806 255978
rect 343862 255922 356518 255978
rect 356574 255922 356642 255978
rect 356698 255922 374154 255978
rect 374210 255922 374278 255978
rect 374334 255922 374402 255978
rect 374458 255922 374526 255978
rect 374582 255922 387238 255978
rect 387294 255922 387362 255978
rect 387418 255922 404874 255978
rect 404930 255922 404998 255978
rect 405054 255922 405122 255978
rect 405178 255922 405246 255978
rect 405302 255922 418518 255978
rect 418574 255922 418642 255978
rect 418698 255922 435594 255978
rect 435650 255922 435718 255978
rect 435774 255922 435842 255978
rect 435898 255922 435966 255978
rect 436022 255922 449238 255978
rect 449294 255922 449362 255978
rect 449418 255922 466314 255978
rect 466370 255922 466438 255978
rect 466494 255922 466562 255978
rect 466618 255922 466686 255978
rect 466742 255922 480518 255978
rect 480574 255922 480642 255978
rect 480698 255922 497034 255978
rect 497090 255922 497158 255978
rect 497214 255922 497282 255978
rect 497338 255922 497406 255978
rect 497462 255922 511238 255978
rect 511294 255922 511362 255978
rect 511418 255922 527754 255978
rect 527810 255922 527878 255978
rect 527934 255922 528002 255978
rect 528058 255922 528126 255978
rect 528182 255922 542518 255978
rect 542574 255922 542642 255978
rect 542698 255922 558474 255978
rect 558530 255922 558598 255978
rect 558654 255922 558722 255978
rect 558778 255922 558846 255978
rect 558902 255922 573238 255978
rect 573294 255922 573362 255978
rect 573418 255922 589194 255978
rect 589250 255922 589318 255978
rect 589374 255922 589442 255978
rect 589498 255922 589566 255978
rect 589622 255922 596496 255978
rect 596552 255922 596620 255978
rect 596676 255922 596744 255978
rect 596800 255922 596868 255978
rect 596924 255922 597980 255978
rect -1916 255826 597980 255922
rect 135196 255358 263860 255374
rect 135196 255302 135212 255358
rect 135268 255302 263788 255358
rect 263844 255302 263860 255358
rect 135196 255286 263860 255302
rect 334668 255358 464564 255374
rect 334668 255302 334684 255358
rect 334740 255302 464492 255358
rect 464548 255302 464564 255358
rect 334668 255286 464564 255302
rect 334444 255178 461204 255194
rect 334444 255122 334460 255178
rect 334516 255122 461132 255178
rect 461188 255122 461204 255178
rect 334444 255106 461204 255122
rect 334332 254998 399044 255014
rect 334332 254942 334348 254998
rect 334404 254942 398972 254998
rect 399028 254942 399044 254998
rect 334332 254926 399044 254942
rect 126796 254458 260388 254474
rect 126796 254402 126812 254458
rect 126868 254402 260316 254458
rect 260372 254402 260388 254458
rect 126796 254386 260388 254402
rect 80428 253558 263860 253574
rect 80428 253502 80444 253558
rect 80500 253502 263788 253558
rect 263844 253502 263860 253558
rect 80428 253486 263860 253502
rect 334444 253558 457172 253574
rect 334444 253502 334460 253558
rect 334516 253502 457100 253558
rect 457156 253502 457172 253558
rect 334444 253486 457172 253502
rect 125116 253378 263972 253394
rect 125116 253322 125132 253378
rect 125188 253322 263900 253378
rect 263956 253322 263972 253378
rect 125116 253306 263972 253322
rect 133516 251938 263860 251954
rect 133516 251882 133532 251938
rect 133588 251882 263788 251938
rect 263844 251882 263860 251938
rect 133516 251866 263860 251882
rect 334444 251938 457284 251954
rect 334444 251882 334460 251938
rect 334516 251882 457212 251938
rect 457268 251882 457284 251938
rect 334444 251866 457284 251882
rect 334332 251758 407444 251774
rect 334332 251702 334348 251758
rect 334404 251702 407372 251758
rect 407428 251702 407444 251758
rect 334332 251686 407444 251702
rect 130156 250318 263860 250334
rect 130156 250262 130172 250318
rect 130228 250262 263788 250318
rect 263844 250262 263860 250318
rect 130156 250246 263860 250262
rect 351020 250318 458964 250334
rect 351020 250262 351036 250318
rect 351092 250262 458892 250318
rect 458948 250262 458964 250318
rect 351020 250246 458964 250262
rect 334444 250138 404084 250154
rect 334444 250082 334460 250138
rect 334516 250082 404012 250138
rect 404068 250082 404084 250138
rect 334444 250066 404084 250082
rect 334444 248518 402404 248534
rect 334444 248462 334460 248518
rect 334516 248462 402332 248518
rect 402388 248462 402404 248518
rect 334444 248446 402404 248462
rect -1916 244350 597980 244446
rect -1916 244294 -1820 244350
rect -1764 244294 -1696 244350
rect -1640 244294 -1572 244350
rect -1516 244294 -1448 244350
rect -1392 244294 9234 244350
rect 9290 244294 9358 244350
rect 9414 244294 9482 244350
rect 9538 244294 9606 244350
rect 9662 244294 70674 244350
rect 70730 244294 70798 244350
rect 70854 244294 70922 244350
rect 70978 244294 71046 244350
rect 71102 244294 132114 244350
rect 132170 244294 132238 244350
rect 132294 244294 132362 244350
rect 132418 244294 132486 244350
rect 132542 244294 162834 244350
rect 162890 244294 162958 244350
rect 163014 244294 163082 244350
rect 163138 244294 163206 244350
rect 163262 244294 193554 244350
rect 193610 244294 193678 244350
rect 193734 244294 193802 244350
rect 193858 244294 193926 244350
rect 193982 244294 224274 244350
rect 224330 244294 224398 244350
rect 224454 244294 224522 244350
rect 224578 244294 224646 244350
rect 224702 244294 254994 244350
rect 255050 244294 255118 244350
rect 255174 244294 255242 244350
rect 255298 244294 255366 244350
rect 255422 244294 287878 244350
rect 287934 244294 288002 244350
rect 288058 244294 318598 244350
rect 318654 244294 318722 244350
rect 318778 244294 347154 244350
rect 347210 244294 347278 244350
rect 347334 244294 347402 244350
rect 347458 244294 347526 244350
rect 347582 244294 377874 244350
rect 377930 244294 377998 244350
rect 378054 244294 378122 244350
rect 378178 244294 378246 244350
rect 378302 244294 408594 244350
rect 408650 244294 408718 244350
rect 408774 244294 408842 244350
rect 408898 244294 408966 244350
rect 409022 244294 439314 244350
rect 439370 244294 439438 244350
rect 439494 244294 439562 244350
rect 439618 244294 439686 244350
rect 439742 244294 470034 244350
rect 470090 244294 470158 244350
rect 470214 244294 470282 244350
rect 470338 244294 470406 244350
rect 470462 244294 500754 244350
rect 500810 244294 500878 244350
rect 500934 244294 501002 244350
rect 501058 244294 501126 244350
rect 501182 244294 531474 244350
rect 531530 244294 531598 244350
rect 531654 244294 531722 244350
rect 531778 244294 531846 244350
rect 531902 244294 562194 244350
rect 562250 244294 562318 244350
rect 562374 244294 562442 244350
rect 562498 244294 562566 244350
rect 562622 244294 592914 244350
rect 592970 244294 593038 244350
rect 593094 244294 593162 244350
rect 593218 244294 593286 244350
rect 593342 244294 597456 244350
rect 597512 244294 597580 244350
rect 597636 244294 597704 244350
rect 597760 244294 597828 244350
rect 597884 244294 597980 244350
rect -1916 244226 597980 244294
rect -1916 244170 -1820 244226
rect -1764 244170 -1696 244226
rect -1640 244170 -1572 244226
rect -1516 244170 -1448 244226
rect -1392 244170 9234 244226
rect 9290 244170 9358 244226
rect 9414 244170 9482 244226
rect 9538 244170 9606 244226
rect 9662 244170 70674 244226
rect 70730 244170 70798 244226
rect 70854 244170 70922 244226
rect 70978 244170 71046 244226
rect 71102 244170 132114 244226
rect 132170 244170 132238 244226
rect 132294 244170 132362 244226
rect 132418 244170 132486 244226
rect 132542 244170 162834 244226
rect 162890 244170 162958 244226
rect 163014 244170 163082 244226
rect 163138 244170 163206 244226
rect 163262 244170 193554 244226
rect 193610 244170 193678 244226
rect 193734 244170 193802 244226
rect 193858 244170 193926 244226
rect 193982 244170 224274 244226
rect 224330 244170 224398 244226
rect 224454 244170 224522 244226
rect 224578 244170 224646 244226
rect 224702 244170 254994 244226
rect 255050 244170 255118 244226
rect 255174 244170 255242 244226
rect 255298 244170 255366 244226
rect 255422 244170 287878 244226
rect 287934 244170 288002 244226
rect 288058 244170 318598 244226
rect 318654 244170 318722 244226
rect 318778 244170 347154 244226
rect 347210 244170 347278 244226
rect 347334 244170 347402 244226
rect 347458 244170 347526 244226
rect 347582 244170 377874 244226
rect 377930 244170 377998 244226
rect 378054 244170 378122 244226
rect 378178 244170 378246 244226
rect 378302 244170 408594 244226
rect 408650 244170 408718 244226
rect 408774 244170 408842 244226
rect 408898 244170 408966 244226
rect 409022 244170 439314 244226
rect 439370 244170 439438 244226
rect 439494 244170 439562 244226
rect 439618 244170 439686 244226
rect 439742 244170 470034 244226
rect 470090 244170 470158 244226
rect 470214 244170 470282 244226
rect 470338 244170 470406 244226
rect 470462 244170 500754 244226
rect 500810 244170 500878 244226
rect 500934 244170 501002 244226
rect 501058 244170 501126 244226
rect 501182 244170 531474 244226
rect 531530 244170 531598 244226
rect 531654 244170 531722 244226
rect 531778 244170 531846 244226
rect 531902 244170 562194 244226
rect 562250 244170 562318 244226
rect 562374 244170 562442 244226
rect 562498 244170 562566 244226
rect 562622 244170 592914 244226
rect 592970 244170 593038 244226
rect 593094 244170 593162 244226
rect 593218 244170 593286 244226
rect 593342 244170 597456 244226
rect 597512 244170 597580 244226
rect 597636 244170 597704 244226
rect 597760 244170 597828 244226
rect 597884 244170 597980 244226
rect -1916 244102 597980 244170
rect -1916 244046 -1820 244102
rect -1764 244046 -1696 244102
rect -1640 244046 -1572 244102
rect -1516 244046 -1448 244102
rect -1392 244046 9234 244102
rect 9290 244046 9358 244102
rect 9414 244046 9482 244102
rect 9538 244046 9606 244102
rect 9662 244046 70674 244102
rect 70730 244046 70798 244102
rect 70854 244046 70922 244102
rect 70978 244046 71046 244102
rect 71102 244046 132114 244102
rect 132170 244046 132238 244102
rect 132294 244046 132362 244102
rect 132418 244046 132486 244102
rect 132542 244046 162834 244102
rect 162890 244046 162958 244102
rect 163014 244046 163082 244102
rect 163138 244046 163206 244102
rect 163262 244046 193554 244102
rect 193610 244046 193678 244102
rect 193734 244046 193802 244102
rect 193858 244046 193926 244102
rect 193982 244046 224274 244102
rect 224330 244046 224398 244102
rect 224454 244046 224522 244102
rect 224578 244046 224646 244102
rect 224702 244046 254994 244102
rect 255050 244046 255118 244102
rect 255174 244046 255242 244102
rect 255298 244046 255366 244102
rect 255422 244046 287878 244102
rect 287934 244046 288002 244102
rect 288058 244046 318598 244102
rect 318654 244046 318722 244102
rect 318778 244046 347154 244102
rect 347210 244046 347278 244102
rect 347334 244046 347402 244102
rect 347458 244046 347526 244102
rect 347582 244046 377874 244102
rect 377930 244046 377998 244102
rect 378054 244046 378122 244102
rect 378178 244046 378246 244102
rect 378302 244046 408594 244102
rect 408650 244046 408718 244102
rect 408774 244046 408842 244102
rect 408898 244046 408966 244102
rect 409022 244046 439314 244102
rect 439370 244046 439438 244102
rect 439494 244046 439562 244102
rect 439618 244046 439686 244102
rect 439742 244046 470034 244102
rect 470090 244046 470158 244102
rect 470214 244046 470282 244102
rect 470338 244046 470406 244102
rect 470462 244046 500754 244102
rect 500810 244046 500878 244102
rect 500934 244046 501002 244102
rect 501058 244046 501126 244102
rect 501182 244046 531474 244102
rect 531530 244046 531598 244102
rect 531654 244046 531722 244102
rect 531778 244046 531846 244102
rect 531902 244046 562194 244102
rect 562250 244046 562318 244102
rect 562374 244046 562442 244102
rect 562498 244046 562566 244102
rect 562622 244046 592914 244102
rect 592970 244046 593038 244102
rect 593094 244046 593162 244102
rect 593218 244046 593286 244102
rect 593342 244046 597456 244102
rect 597512 244046 597580 244102
rect 597636 244046 597704 244102
rect 597760 244046 597828 244102
rect 597884 244046 597980 244102
rect -1916 243978 597980 244046
rect -1916 243922 -1820 243978
rect -1764 243922 -1696 243978
rect -1640 243922 -1572 243978
rect -1516 243922 -1448 243978
rect -1392 243922 9234 243978
rect 9290 243922 9358 243978
rect 9414 243922 9482 243978
rect 9538 243922 9606 243978
rect 9662 243922 70674 243978
rect 70730 243922 70798 243978
rect 70854 243922 70922 243978
rect 70978 243922 71046 243978
rect 71102 243922 132114 243978
rect 132170 243922 132238 243978
rect 132294 243922 132362 243978
rect 132418 243922 132486 243978
rect 132542 243922 162834 243978
rect 162890 243922 162958 243978
rect 163014 243922 163082 243978
rect 163138 243922 163206 243978
rect 163262 243922 193554 243978
rect 193610 243922 193678 243978
rect 193734 243922 193802 243978
rect 193858 243922 193926 243978
rect 193982 243922 224274 243978
rect 224330 243922 224398 243978
rect 224454 243922 224522 243978
rect 224578 243922 224646 243978
rect 224702 243922 254994 243978
rect 255050 243922 255118 243978
rect 255174 243922 255242 243978
rect 255298 243922 255366 243978
rect 255422 243922 287878 243978
rect 287934 243922 288002 243978
rect 288058 243922 318598 243978
rect 318654 243922 318722 243978
rect 318778 243922 347154 243978
rect 347210 243922 347278 243978
rect 347334 243922 347402 243978
rect 347458 243922 347526 243978
rect 347582 243922 377874 243978
rect 377930 243922 377998 243978
rect 378054 243922 378122 243978
rect 378178 243922 378246 243978
rect 378302 243922 408594 243978
rect 408650 243922 408718 243978
rect 408774 243922 408842 243978
rect 408898 243922 408966 243978
rect 409022 243922 439314 243978
rect 439370 243922 439438 243978
rect 439494 243922 439562 243978
rect 439618 243922 439686 243978
rect 439742 243922 470034 243978
rect 470090 243922 470158 243978
rect 470214 243922 470282 243978
rect 470338 243922 470406 243978
rect 470462 243922 500754 243978
rect 500810 243922 500878 243978
rect 500934 243922 501002 243978
rect 501058 243922 501126 243978
rect 501182 243922 531474 243978
rect 531530 243922 531598 243978
rect 531654 243922 531722 243978
rect 531778 243922 531846 243978
rect 531902 243922 562194 243978
rect 562250 243922 562318 243978
rect 562374 243922 562442 243978
rect 562498 243922 562566 243978
rect 562622 243922 592914 243978
rect 592970 243922 593038 243978
rect 593094 243922 593162 243978
rect 593218 243922 593286 243978
rect 593342 243922 597456 243978
rect 597512 243922 597580 243978
rect 597636 243922 597704 243978
rect 597760 243922 597828 243978
rect 597884 243922 597980 243978
rect -1916 243826 597980 243922
rect -1916 238350 597980 238446
rect -1916 238294 -860 238350
rect -804 238294 -736 238350
rect -680 238294 -612 238350
rect -556 238294 -488 238350
rect -432 238294 5514 238350
rect 5570 238294 5638 238350
rect 5694 238294 5762 238350
rect 5818 238294 5886 238350
rect 5942 238294 36234 238350
rect 36290 238294 36358 238350
rect 36414 238294 36482 238350
rect 36538 238294 36606 238350
rect 36662 238294 66954 238350
rect 67010 238294 67078 238350
rect 67134 238294 67202 238350
rect 67258 238294 67326 238350
rect 67382 238294 97674 238350
rect 97730 238294 97798 238350
rect 97854 238294 97922 238350
rect 97978 238294 98046 238350
rect 98102 238294 128394 238350
rect 128450 238294 128518 238350
rect 128574 238294 128642 238350
rect 128698 238294 128766 238350
rect 128822 238294 159114 238350
rect 159170 238294 159238 238350
rect 159294 238294 159362 238350
rect 159418 238294 159486 238350
rect 159542 238294 189834 238350
rect 189890 238294 189958 238350
rect 190014 238294 190082 238350
rect 190138 238294 190206 238350
rect 190262 238294 220554 238350
rect 220610 238294 220678 238350
rect 220734 238294 220802 238350
rect 220858 238294 220926 238350
rect 220982 238294 251274 238350
rect 251330 238294 251398 238350
rect 251454 238294 251522 238350
rect 251578 238294 251646 238350
rect 251702 238294 272518 238350
rect 272574 238294 272642 238350
rect 272698 238294 303238 238350
rect 303294 238294 303362 238350
rect 303418 238294 343434 238350
rect 343490 238294 343558 238350
rect 343614 238294 343682 238350
rect 343738 238294 343806 238350
rect 343862 238294 374154 238350
rect 374210 238294 374278 238350
rect 374334 238294 374402 238350
rect 374458 238294 374526 238350
rect 374582 238294 404874 238350
rect 404930 238294 404998 238350
rect 405054 238294 405122 238350
rect 405178 238294 405246 238350
rect 405302 238294 435594 238350
rect 435650 238294 435718 238350
rect 435774 238294 435842 238350
rect 435898 238294 435966 238350
rect 436022 238294 466314 238350
rect 466370 238294 466438 238350
rect 466494 238294 466562 238350
rect 466618 238294 466686 238350
rect 466742 238294 497034 238350
rect 497090 238294 497158 238350
rect 497214 238294 497282 238350
rect 497338 238294 497406 238350
rect 497462 238294 527754 238350
rect 527810 238294 527878 238350
rect 527934 238294 528002 238350
rect 528058 238294 528126 238350
rect 528182 238294 558474 238350
rect 558530 238294 558598 238350
rect 558654 238294 558722 238350
rect 558778 238294 558846 238350
rect 558902 238294 589194 238350
rect 589250 238294 589318 238350
rect 589374 238294 589442 238350
rect 589498 238294 589566 238350
rect 589622 238294 596496 238350
rect 596552 238294 596620 238350
rect 596676 238294 596744 238350
rect 596800 238294 596868 238350
rect 596924 238294 597980 238350
rect -1916 238226 597980 238294
rect -1916 238170 -860 238226
rect -804 238170 -736 238226
rect -680 238170 -612 238226
rect -556 238170 -488 238226
rect -432 238170 5514 238226
rect 5570 238170 5638 238226
rect 5694 238170 5762 238226
rect 5818 238170 5886 238226
rect 5942 238170 36234 238226
rect 36290 238170 36358 238226
rect 36414 238170 36482 238226
rect 36538 238170 36606 238226
rect 36662 238170 66954 238226
rect 67010 238170 67078 238226
rect 67134 238170 67202 238226
rect 67258 238170 67326 238226
rect 67382 238170 97674 238226
rect 97730 238170 97798 238226
rect 97854 238170 97922 238226
rect 97978 238170 98046 238226
rect 98102 238170 128394 238226
rect 128450 238170 128518 238226
rect 128574 238170 128642 238226
rect 128698 238170 128766 238226
rect 128822 238170 159114 238226
rect 159170 238170 159238 238226
rect 159294 238170 159362 238226
rect 159418 238170 159486 238226
rect 159542 238170 189834 238226
rect 189890 238170 189958 238226
rect 190014 238170 190082 238226
rect 190138 238170 190206 238226
rect 190262 238170 220554 238226
rect 220610 238170 220678 238226
rect 220734 238170 220802 238226
rect 220858 238170 220926 238226
rect 220982 238170 251274 238226
rect 251330 238170 251398 238226
rect 251454 238170 251522 238226
rect 251578 238170 251646 238226
rect 251702 238170 272518 238226
rect 272574 238170 272642 238226
rect 272698 238170 303238 238226
rect 303294 238170 303362 238226
rect 303418 238170 343434 238226
rect 343490 238170 343558 238226
rect 343614 238170 343682 238226
rect 343738 238170 343806 238226
rect 343862 238170 374154 238226
rect 374210 238170 374278 238226
rect 374334 238170 374402 238226
rect 374458 238170 374526 238226
rect 374582 238170 404874 238226
rect 404930 238170 404998 238226
rect 405054 238170 405122 238226
rect 405178 238170 405246 238226
rect 405302 238170 435594 238226
rect 435650 238170 435718 238226
rect 435774 238170 435842 238226
rect 435898 238170 435966 238226
rect 436022 238170 466314 238226
rect 466370 238170 466438 238226
rect 466494 238170 466562 238226
rect 466618 238170 466686 238226
rect 466742 238170 497034 238226
rect 497090 238170 497158 238226
rect 497214 238170 497282 238226
rect 497338 238170 497406 238226
rect 497462 238170 527754 238226
rect 527810 238170 527878 238226
rect 527934 238170 528002 238226
rect 528058 238170 528126 238226
rect 528182 238170 558474 238226
rect 558530 238170 558598 238226
rect 558654 238170 558722 238226
rect 558778 238170 558846 238226
rect 558902 238170 589194 238226
rect 589250 238170 589318 238226
rect 589374 238170 589442 238226
rect 589498 238170 589566 238226
rect 589622 238170 596496 238226
rect 596552 238170 596620 238226
rect 596676 238170 596744 238226
rect 596800 238170 596868 238226
rect 596924 238170 597980 238226
rect -1916 238102 597980 238170
rect -1916 238046 -860 238102
rect -804 238046 -736 238102
rect -680 238046 -612 238102
rect -556 238046 -488 238102
rect -432 238046 5514 238102
rect 5570 238046 5638 238102
rect 5694 238046 5762 238102
rect 5818 238046 5886 238102
rect 5942 238046 36234 238102
rect 36290 238046 36358 238102
rect 36414 238046 36482 238102
rect 36538 238046 36606 238102
rect 36662 238046 66954 238102
rect 67010 238046 67078 238102
rect 67134 238046 67202 238102
rect 67258 238046 67326 238102
rect 67382 238046 97674 238102
rect 97730 238046 97798 238102
rect 97854 238046 97922 238102
rect 97978 238046 98046 238102
rect 98102 238046 128394 238102
rect 128450 238046 128518 238102
rect 128574 238046 128642 238102
rect 128698 238046 128766 238102
rect 128822 238046 159114 238102
rect 159170 238046 159238 238102
rect 159294 238046 159362 238102
rect 159418 238046 159486 238102
rect 159542 238046 189834 238102
rect 189890 238046 189958 238102
rect 190014 238046 190082 238102
rect 190138 238046 190206 238102
rect 190262 238046 220554 238102
rect 220610 238046 220678 238102
rect 220734 238046 220802 238102
rect 220858 238046 220926 238102
rect 220982 238046 251274 238102
rect 251330 238046 251398 238102
rect 251454 238046 251522 238102
rect 251578 238046 251646 238102
rect 251702 238046 272518 238102
rect 272574 238046 272642 238102
rect 272698 238046 303238 238102
rect 303294 238046 303362 238102
rect 303418 238046 343434 238102
rect 343490 238046 343558 238102
rect 343614 238046 343682 238102
rect 343738 238046 343806 238102
rect 343862 238046 374154 238102
rect 374210 238046 374278 238102
rect 374334 238046 374402 238102
rect 374458 238046 374526 238102
rect 374582 238046 404874 238102
rect 404930 238046 404998 238102
rect 405054 238046 405122 238102
rect 405178 238046 405246 238102
rect 405302 238046 435594 238102
rect 435650 238046 435718 238102
rect 435774 238046 435842 238102
rect 435898 238046 435966 238102
rect 436022 238046 466314 238102
rect 466370 238046 466438 238102
rect 466494 238046 466562 238102
rect 466618 238046 466686 238102
rect 466742 238046 497034 238102
rect 497090 238046 497158 238102
rect 497214 238046 497282 238102
rect 497338 238046 497406 238102
rect 497462 238046 527754 238102
rect 527810 238046 527878 238102
rect 527934 238046 528002 238102
rect 528058 238046 528126 238102
rect 528182 238046 558474 238102
rect 558530 238046 558598 238102
rect 558654 238046 558722 238102
rect 558778 238046 558846 238102
rect 558902 238046 589194 238102
rect 589250 238046 589318 238102
rect 589374 238046 589442 238102
rect 589498 238046 589566 238102
rect 589622 238046 596496 238102
rect 596552 238046 596620 238102
rect 596676 238046 596744 238102
rect 596800 238046 596868 238102
rect 596924 238046 597980 238102
rect -1916 237978 597980 238046
rect -1916 237922 -860 237978
rect -804 237922 -736 237978
rect -680 237922 -612 237978
rect -556 237922 -488 237978
rect -432 237922 5514 237978
rect 5570 237922 5638 237978
rect 5694 237922 5762 237978
rect 5818 237922 5886 237978
rect 5942 237922 36234 237978
rect 36290 237922 36358 237978
rect 36414 237922 36482 237978
rect 36538 237922 36606 237978
rect 36662 237922 66954 237978
rect 67010 237922 67078 237978
rect 67134 237922 67202 237978
rect 67258 237922 67326 237978
rect 67382 237922 97674 237978
rect 97730 237922 97798 237978
rect 97854 237922 97922 237978
rect 97978 237922 98046 237978
rect 98102 237922 128394 237978
rect 128450 237922 128518 237978
rect 128574 237922 128642 237978
rect 128698 237922 128766 237978
rect 128822 237922 159114 237978
rect 159170 237922 159238 237978
rect 159294 237922 159362 237978
rect 159418 237922 159486 237978
rect 159542 237922 189834 237978
rect 189890 237922 189958 237978
rect 190014 237922 190082 237978
rect 190138 237922 190206 237978
rect 190262 237922 220554 237978
rect 220610 237922 220678 237978
rect 220734 237922 220802 237978
rect 220858 237922 220926 237978
rect 220982 237922 251274 237978
rect 251330 237922 251398 237978
rect 251454 237922 251522 237978
rect 251578 237922 251646 237978
rect 251702 237922 272518 237978
rect 272574 237922 272642 237978
rect 272698 237922 303238 237978
rect 303294 237922 303362 237978
rect 303418 237922 343434 237978
rect 343490 237922 343558 237978
rect 343614 237922 343682 237978
rect 343738 237922 343806 237978
rect 343862 237922 374154 237978
rect 374210 237922 374278 237978
rect 374334 237922 374402 237978
rect 374458 237922 374526 237978
rect 374582 237922 404874 237978
rect 404930 237922 404998 237978
rect 405054 237922 405122 237978
rect 405178 237922 405246 237978
rect 405302 237922 435594 237978
rect 435650 237922 435718 237978
rect 435774 237922 435842 237978
rect 435898 237922 435966 237978
rect 436022 237922 466314 237978
rect 466370 237922 466438 237978
rect 466494 237922 466562 237978
rect 466618 237922 466686 237978
rect 466742 237922 497034 237978
rect 497090 237922 497158 237978
rect 497214 237922 497282 237978
rect 497338 237922 497406 237978
rect 497462 237922 527754 237978
rect 527810 237922 527878 237978
rect 527934 237922 528002 237978
rect 528058 237922 528126 237978
rect 528182 237922 558474 237978
rect 558530 237922 558598 237978
rect 558654 237922 558722 237978
rect 558778 237922 558846 237978
rect 558902 237922 589194 237978
rect 589250 237922 589318 237978
rect 589374 237922 589442 237978
rect 589498 237922 589566 237978
rect 589622 237922 596496 237978
rect 596552 237922 596620 237978
rect 596676 237922 596744 237978
rect 596800 237922 596868 237978
rect 596924 237922 597980 237978
rect -1916 237826 597980 237922
rect -1916 226350 597980 226446
rect -1916 226294 -1820 226350
rect -1764 226294 -1696 226350
rect -1640 226294 -1572 226350
rect -1516 226294 -1448 226350
rect -1392 226294 9234 226350
rect 9290 226294 9358 226350
rect 9414 226294 9482 226350
rect 9538 226294 9606 226350
rect 9662 226294 70674 226350
rect 70730 226294 70798 226350
rect 70854 226294 70922 226350
rect 70978 226294 71046 226350
rect 71102 226294 132114 226350
rect 132170 226294 132238 226350
rect 132294 226294 132362 226350
rect 132418 226294 132486 226350
rect 132542 226294 162834 226350
rect 162890 226294 162958 226350
rect 163014 226294 163082 226350
rect 163138 226294 163206 226350
rect 163262 226294 193554 226350
rect 193610 226294 193678 226350
rect 193734 226294 193802 226350
rect 193858 226294 193926 226350
rect 193982 226294 224274 226350
rect 224330 226294 224398 226350
rect 224454 226294 224522 226350
rect 224578 226294 224646 226350
rect 224702 226294 254994 226350
rect 255050 226294 255118 226350
rect 255174 226294 255242 226350
rect 255298 226294 255366 226350
rect 255422 226294 287878 226350
rect 287934 226294 288002 226350
rect 288058 226294 318598 226350
rect 318654 226294 318722 226350
rect 318778 226294 347154 226350
rect 347210 226294 347278 226350
rect 347334 226294 347402 226350
rect 347458 226294 347526 226350
rect 347582 226294 377874 226350
rect 377930 226294 377998 226350
rect 378054 226294 378122 226350
rect 378178 226294 378246 226350
rect 378302 226294 408594 226350
rect 408650 226294 408718 226350
rect 408774 226294 408842 226350
rect 408898 226294 408966 226350
rect 409022 226294 439314 226350
rect 439370 226294 439438 226350
rect 439494 226294 439562 226350
rect 439618 226294 439686 226350
rect 439742 226294 470034 226350
rect 470090 226294 470158 226350
rect 470214 226294 470282 226350
rect 470338 226294 470406 226350
rect 470462 226294 500754 226350
rect 500810 226294 500878 226350
rect 500934 226294 501002 226350
rect 501058 226294 501126 226350
rect 501182 226294 531474 226350
rect 531530 226294 531598 226350
rect 531654 226294 531722 226350
rect 531778 226294 531846 226350
rect 531902 226294 562194 226350
rect 562250 226294 562318 226350
rect 562374 226294 562442 226350
rect 562498 226294 562566 226350
rect 562622 226294 592914 226350
rect 592970 226294 593038 226350
rect 593094 226294 593162 226350
rect 593218 226294 593286 226350
rect 593342 226294 597456 226350
rect 597512 226294 597580 226350
rect 597636 226294 597704 226350
rect 597760 226294 597828 226350
rect 597884 226294 597980 226350
rect -1916 226226 597980 226294
rect -1916 226170 -1820 226226
rect -1764 226170 -1696 226226
rect -1640 226170 -1572 226226
rect -1516 226170 -1448 226226
rect -1392 226170 9234 226226
rect 9290 226170 9358 226226
rect 9414 226170 9482 226226
rect 9538 226170 9606 226226
rect 9662 226170 70674 226226
rect 70730 226170 70798 226226
rect 70854 226170 70922 226226
rect 70978 226170 71046 226226
rect 71102 226170 132114 226226
rect 132170 226170 132238 226226
rect 132294 226170 132362 226226
rect 132418 226170 132486 226226
rect 132542 226170 162834 226226
rect 162890 226170 162958 226226
rect 163014 226170 163082 226226
rect 163138 226170 163206 226226
rect 163262 226170 193554 226226
rect 193610 226170 193678 226226
rect 193734 226170 193802 226226
rect 193858 226170 193926 226226
rect 193982 226170 224274 226226
rect 224330 226170 224398 226226
rect 224454 226170 224522 226226
rect 224578 226170 224646 226226
rect 224702 226170 254994 226226
rect 255050 226170 255118 226226
rect 255174 226170 255242 226226
rect 255298 226170 255366 226226
rect 255422 226170 287878 226226
rect 287934 226170 288002 226226
rect 288058 226170 318598 226226
rect 318654 226170 318722 226226
rect 318778 226170 347154 226226
rect 347210 226170 347278 226226
rect 347334 226170 347402 226226
rect 347458 226170 347526 226226
rect 347582 226170 377874 226226
rect 377930 226170 377998 226226
rect 378054 226170 378122 226226
rect 378178 226170 378246 226226
rect 378302 226170 408594 226226
rect 408650 226170 408718 226226
rect 408774 226170 408842 226226
rect 408898 226170 408966 226226
rect 409022 226170 439314 226226
rect 439370 226170 439438 226226
rect 439494 226170 439562 226226
rect 439618 226170 439686 226226
rect 439742 226170 470034 226226
rect 470090 226170 470158 226226
rect 470214 226170 470282 226226
rect 470338 226170 470406 226226
rect 470462 226170 500754 226226
rect 500810 226170 500878 226226
rect 500934 226170 501002 226226
rect 501058 226170 501126 226226
rect 501182 226170 531474 226226
rect 531530 226170 531598 226226
rect 531654 226170 531722 226226
rect 531778 226170 531846 226226
rect 531902 226170 562194 226226
rect 562250 226170 562318 226226
rect 562374 226170 562442 226226
rect 562498 226170 562566 226226
rect 562622 226170 592914 226226
rect 592970 226170 593038 226226
rect 593094 226170 593162 226226
rect 593218 226170 593286 226226
rect 593342 226170 597456 226226
rect 597512 226170 597580 226226
rect 597636 226170 597704 226226
rect 597760 226170 597828 226226
rect 597884 226170 597980 226226
rect -1916 226102 597980 226170
rect -1916 226046 -1820 226102
rect -1764 226046 -1696 226102
rect -1640 226046 -1572 226102
rect -1516 226046 -1448 226102
rect -1392 226046 9234 226102
rect 9290 226046 9358 226102
rect 9414 226046 9482 226102
rect 9538 226046 9606 226102
rect 9662 226046 70674 226102
rect 70730 226046 70798 226102
rect 70854 226046 70922 226102
rect 70978 226046 71046 226102
rect 71102 226046 132114 226102
rect 132170 226046 132238 226102
rect 132294 226046 132362 226102
rect 132418 226046 132486 226102
rect 132542 226046 162834 226102
rect 162890 226046 162958 226102
rect 163014 226046 163082 226102
rect 163138 226046 163206 226102
rect 163262 226046 193554 226102
rect 193610 226046 193678 226102
rect 193734 226046 193802 226102
rect 193858 226046 193926 226102
rect 193982 226046 224274 226102
rect 224330 226046 224398 226102
rect 224454 226046 224522 226102
rect 224578 226046 224646 226102
rect 224702 226046 254994 226102
rect 255050 226046 255118 226102
rect 255174 226046 255242 226102
rect 255298 226046 255366 226102
rect 255422 226046 287878 226102
rect 287934 226046 288002 226102
rect 288058 226046 318598 226102
rect 318654 226046 318722 226102
rect 318778 226046 347154 226102
rect 347210 226046 347278 226102
rect 347334 226046 347402 226102
rect 347458 226046 347526 226102
rect 347582 226046 377874 226102
rect 377930 226046 377998 226102
rect 378054 226046 378122 226102
rect 378178 226046 378246 226102
rect 378302 226046 408594 226102
rect 408650 226046 408718 226102
rect 408774 226046 408842 226102
rect 408898 226046 408966 226102
rect 409022 226046 439314 226102
rect 439370 226046 439438 226102
rect 439494 226046 439562 226102
rect 439618 226046 439686 226102
rect 439742 226046 470034 226102
rect 470090 226046 470158 226102
rect 470214 226046 470282 226102
rect 470338 226046 470406 226102
rect 470462 226046 500754 226102
rect 500810 226046 500878 226102
rect 500934 226046 501002 226102
rect 501058 226046 501126 226102
rect 501182 226046 531474 226102
rect 531530 226046 531598 226102
rect 531654 226046 531722 226102
rect 531778 226046 531846 226102
rect 531902 226046 562194 226102
rect 562250 226046 562318 226102
rect 562374 226046 562442 226102
rect 562498 226046 562566 226102
rect 562622 226046 592914 226102
rect 592970 226046 593038 226102
rect 593094 226046 593162 226102
rect 593218 226046 593286 226102
rect 593342 226046 597456 226102
rect 597512 226046 597580 226102
rect 597636 226046 597704 226102
rect 597760 226046 597828 226102
rect 597884 226046 597980 226102
rect -1916 225978 597980 226046
rect -1916 225922 -1820 225978
rect -1764 225922 -1696 225978
rect -1640 225922 -1572 225978
rect -1516 225922 -1448 225978
rect -1392 225922 9234 225978
rect 9290 225922 9358 225978
rect 9414 225922 9482 225978
rect 9538 225922 9606 225978
rect 9662 225922 70674 225978
rect 70730 225922 70798 225978
rect 70854 225922 70922 225978
rect 70978 225922 71046 225978
rect 71102 225922 132114 225978
rect 132170 225922 132238 225978
rect 132294 225922 132362 225978
rect 132418 225922 132486 225978
rect 132542 225922 162834 225978
rect 162890 225922 162958 225978
rect 163014 225922 163082 225978
rect 163138 225922 163206 225978
rect 163262 225922 193554 225978
rect 193610 225922 193678 225978
rect 193734 225922 193802 225978
rect 193858 225922 193926 225978
rect 193982 225922 224274 225978
rect 224330 225922 224398 225978
rect 224454 225922 224522 225978
rect 224578 225922 224646 225978
rect 224702 225922 254994 225978
rect 255050 225922 255118 225978
rect 255174 225922 255242 225978
rect 255298 225922 255366 225978
rect 255422 225922 287878 225978
rect 287934 225922 288002 225978
rect 288058 225922 318598 225978
rect 318654 225922 318722 225978
rect 318778 225922 347154 225978
rect 347210 225922 347278 225978
rect 347334 225922 347402 225978
rect 347458 225922 347526 225978
rect 347582 225922 377874 225978
rect 377930 225922 377998 225978
rect 378054 225922 378122 225978
rect 378178 225922 378246 225978
rect 378302 225922 408594 225978
rect 408650 225922 408718 225978
rect 408774 225922 408842 225978
rect 408898 225922 408966 225978
rect 409022 225922 439314 225978
rect 439370 225922 439438 225978
rect 439494 225922 439562 225978
rect 439618 225922 439686 225978
rect 439742 225922 470034 225978
rect 470090 225922 470158 225978
rect 470214 225922 470282 225978
rect 470338 225922 470406 225978
rect 470462 225922 500754 225978
rect 500810 225922 500878 225978
rect 500934 225922 501002 225978
rect 501058 225922 501126 225978
rect 501182 225922 531474 225978
rect 531530 225922 531598 225978
rect 531654 225922 531722 225978
rect 531778 225922 531846 225978
rect 531902 225922 562194 225978
rect 562250 225922 562318 225978
rect 562374 225922 562442 225978
rect 562498 225922 562566 225978
rect 562622 225922 592914 225978
rect 592970 225922 593038 225978
rect 593094 225922 593162 225978
rect 593218 225922 593286 225978
rect 593342 225922 597456 225978
rect 597512 225922 597580 225978
rect 597636 225922 597704 225978
rect 597760 225922 597828 225978
rect 597884 225922 597980 225978
rect -1916 225826 597980 225922
rect -1916 220350 597980 220446
rect -1916 220294 -860 220350
rect -804 220294 -736 220350
rect -680 220294 -612 220350
rect -556 220294 -488 220350
rect -432 220294 5514 220350
rect 5570 220294 5638 220350
rect 5694 220294 5762 220350
rect 5818 220294 5886 220350
rect 5942 220294 36234 220350
rect 36290 220294 36358 220350
rect 36414 220294 36482 220350
rect 36538 220294 36606 220350
rect 36662 220294 66954 220350
rect 67010 220294 67078 220350
rect 67134 220294 67202 220350
rect 67258 220294 67326 220350
rect 67382 220294 97674 220350
rect 97730 220294 97798 220350
rect 97854 220294 97922 220350
rect 97978 220294 98046 220350
rect 98102 220294 128394 220350
rect 128450 220294 128518 220350
rect 128574 220294 128642 220350
rect 128698 220294 128766 220350
rect 128822 220294 159114 220350
rect 159170 220294 159238 220350
rect 159294 220294 159362 220350
rect 159418 220294 159486 220350
rect 159542 220294 189834 220350
rect 189890 220294 189958 220350
rect 190014 220294 190082 220350
rect 190138 220294 190206 220350
rect 190262 220294 220554 220350
rect 220610 220294 220678 220350
rect 220734 220294 220802 220350
rect 220858 220294 220926 220350
rect 220982 220294 251274 220350
rect 251330 220294 251398 220350
rect 251454 220294 251522 220350
rect 251578 220294 251646 220350
rect 251702 220294 272518 220350
rect 272574 220294 272642 220350
rect 272698 220294 303238 220350
rect 303294 220294 303362 220350
rect 303418 220294 343434 220350
rect 343490 220294 343558 220350
rect 343614 220294 343682 220350
rect 343738 220294 343806 220350
rect 343862 220294 374154 220350
rect 374210 220294 374278 220350
rect 374334 220294 374402 220350
rect 374458 220294 374526 220350
rect 374582 220294 404874 220350
rect 404930 220294 404998 220350
rect 405054 220294 405122 220350
rect 405178 220294 405246 220350
rect 405302 220294 435594 220350
rect 435650 220294 435718 220350
rect 435774 220294 435842 220350
rect 435898 220294 435966 220350
rect 436022 220294 466314 220350
rect 466370 220294 466438 220350
rect 466494 220294 466562 220350
rect 466618 220294 466686 220350
rect 466742 220294 497034 220350
rect 497090 220294 497158 220350
rect 497214 220294 497282 220350
rect 497338 220294 497406 220350
rect 497462 220294 527754 220350
rect 527810 220294 527878 220350
rect 527934 220294 528002 220350
rect 528058 220294 528126 220350
rect 528182 220294 558474 220350
rect 558530 220294 558598 220350
rect 558654 220294 558722 220350
rect 558778 220294 558846 220350
rect 558902 220294 589194 220350
rect 589250 220294 589318 220350
rect 589374 220294 589442 220350
rect 589498 220294 589566 220350
rect 589622 220294 596496 220350
rect 596552 220294 596620 220350
rect 596676 220294 596744 220350
rect 596800 220294 596868 220350
rect 596924 220294 597980 220350
rect -1916 220226 597980 220294
rect -1916 220170 -860 220226
rect -804 220170 -736 220226
rect -680 220170 -612 220226
rect -556 220170 -488 220226
rect -432 220170 5514 220226
rect 5570 220170 5638 220226
rect 5694 220170 5762 220226
rect 5818 220170 5886 220226
rect 5942 220170 36234 220226
rect 36290 220170 36358 220226
rect 36414 220170 36482 220226
rect 36538 220170 36606 220226
rect 36662 220170 66954 220226
rect 67010 220170 67078 220226
rect 67134 220170 67202 220226
rect 67258 220170 67326 220226
rect 67382 220170 97674 220226
rect 97730 220170 97798 220226
rect 97854 220170 97922 220226
rect 97978 220170 98046 220226
rect 98102 220170 128394 220226
rect 128450 220170 128518 220226
rect 128574 220170 128642 220226
rect 128698 220170 128766 220226
rect 128822 220170 159114 220226
rect 159170 220170 159238 220226
rect 159294 220170 159362 220226
rect 159418 220170 159486 220226
rect 159542 220170 189834 220226
rect 189890 220170 189958 220226
rect 190014 220170 190082 220226
rect 190138 220170 190206 220226
rect 190262 220170 220554 220226
rect 220610 220170 220678 220226
rect 220734 220170 220802 220226
rect 220858 220170 220926 220226
rect 220982 220170 251274 220226
rect 251330 220170 251398 220226
rect 251454 220170 251522 220226
rect 251578 220170 251646 220226
rect 251702 220170 272518 220226
rect 272574 220170 272642 220226
rect 272698 220170 303238 220226
rect 303294 220170 303362 220226
rect 303418 220170 343434 220226
rect 343490 220170 343558 220226
rect 343614 220170 343682 220226
rect 343738 220170 343806 220226
rect 343862 220170 374154 220226
rect 374210 220170 374278 220226
rect 374334 220170 374402 220226
rect 374458 220170 374526 220226
rect 374582 220170 404874 220226
rect 404930 220170 404998 220226
rect 405054 220170 405122 220226
rect 405178 220170 405246 220226
rect 405302 220170 435594 220226
rect 435650 220170 435718 220226
rect 435774 220170 435842 220226
rect 435898 220170 435966 220226
rect 436022 220170 466314 220226
rect 466370 220170 466438 220226
rect 466494 220170 466562 220226
rect 466618 220170 466686 220226
rect 466742 220170 497034 220226
rect 497090 220170 497158 220226
rect 497214 220170 497282 220226
rect 497338 220170 497406 220226
rect 497462 220170 527754 220226
rect 527810 220170 527878 220226
rect 527934 220170 528002 220226
rect 528058 220170 528126 220226
rect 528182 220170 558474 220226
rect 558530 220170 558598 220226
rect 558654 220170 558722 220226
rect 558778 220170 558846 220226
rect 558902 220170 589194 220226
rect 589250 220170 589318 220226
rect 589374 220170 589442 220226
rect 589498 220170 589566 220226
rect 589622 220170 596496 220226
rect 596552 220170 596620 220226
rect 596676 220170 596744 220226
rect 596800 220170 596868 220226
rect 596924 220170 597980 220226
rect -1916 220102 597980 220170
rect -1916 220046 -860 220102
rect -804 220046 -736 220102
rect -680 220046 -612 220102
rect -556 220046 -488 220102
rect -432 220046 5514 220102
rect 5570 220046 5638 220102
rect 5694 220046 5762 220102
rect 5818 220046 5886 220102
rect 5942 220046 36234 220102
rect 36290 220046 36358 220102
rect 36414 220046 36482 220102
rect 36538 220046 36606 220102
rect 36662 220046 66954 220102
rect 67010 220046 67078 220102
rect 67134 220046 67202 220102
rect 67258 220046 67326 220102
rect 67382 220046 97674 220102
rect 97730 220046 97798 220102
rect 97854 220046 97922 220102
rect 97978 220046 98046 220102
rect 98102 220046 128394 220102
rect 128450 220046 128518 220102
rect 128574 220046 128642 220102
rect 128698 220046 128766 220102
rect 128822 220046 159114 220102
rect 159170 220046 159238 220102
rect 159294 220046 159362 220102
rect 159418 220046 159486 220102
rect 159542 220046 189834 220102
rect 189890 220046 189958 220102
rect 190014 220046 190082 220102
rect 190138 220046 190206 220102
rect 190262 220046 220554 220102
rect 220610 220046 220678 220102
rect 220734 220046 220802 220102
rect 220858 220046 220926 220102
rect 220982 220046 251274 220102
rect 251330 220046 251398 220102
rect 251454 220046 251522 220102
rect 251578 220046 251646 220102
rect 251702 220046 272518 220102
rect 272574 220046 272642 220102
rect 272698 220046 303238 220102
rect 303294 220046 303362 220102
rect 303418 220046 343434 220102
rect 343490 220046 343558 220102
rect 343614 220046 343682 220102
rect 343738 220046 343806 220102
rect 343862 220046 374154 220102
rect 374210 220046 374278 220102
rect 374334 220046 374402 220102
rect 374458 220046 374526 220102
rect 374582 220046 404874 220102
rect 404930 220046 404998 220102
rect 405054 220046 405122 220102
rect 405178 220046 405246 220102
rect 405302 220046 435594 220102
rect 435650 220046 435718 220102
rect 435774 220046 435842 220102
rect 435898 220046 435966 220102
rect 436022 220046 466314 220102
rect 466370 220046 466438 220102
rect 466494 220046 466562 220102
rect 466618 220046 466686 220102
rect 466742 220046 497034 220102
rect 497090 220046 497158 220102
rect 497214 220046 497282 220102
rect 497338 220046 497406 220102
rect 497462 220046 527754 220102
rect 527810 220046 527878 220102
rect 527934 220046 528002 220102
rect 528058 220046 528126 220102
rect 528182 220046 558474 220102
rect 558530 220046 558598 220102
rect 558654 220046 558722 220102
rect 558778 220046 558846 220102
rect 558902 220046 589194 220102
rect 589250 220046 589318 220102
rect 589374 220046 589442 220102
rect 589498 220046 589566 220102
rect 589622 220046 596496 220102
rect 596552 220046 596620 220102
rect 596676 220046 596744 220102
rect 596800 220046 596868 220102
rect 596924 220046 597980 220102
rect -1916 219978 597980 220046
rect -1916 219922 -860 219978
rect -804 219922 -736 219978
rect -680 219922 -612 219978
rect -556 219922 -488 219978
rect -432 219922 5514 219978
rect 5570 219922 5638 219978
rect 5694 219922 5762 219978
rect 5818 219922 5886 219978
rect 5942 219922 36234 219978
rect 36290 219922 36358 219978
rect 36414 219922 36482 219978
rect 36538 219922 36606 219978
rect 36662 219922 66954 219978
rect 67010 219922 67078 219978
rect 67134 219922 67202 219978
rect 67258 219922 67326 219978
rect 67382 219922 97674 219978
rect 97730 219922 97798 219978
rect 97854 219922 97922 219978
rect 97978 219922 98046 219978
rect 98102 219922 128394 219978
rect 128450 219922 128518 219978
rect 128574 219922 128642 219978
rect 128698 219922 128766 219978
rect 128822 219922 159114 219978
rect 159170 219922 159238 219978
rect 159294 219922 159362 219978
rect 159418 219922 159486 219978
rect 159542 219922 189834 219978
rect 189890 219922 189958 219978
rect 190014 219922 190082 219978
rect 190138 219922 190206 219978
rect 190262 219922 220554 219978
rect 220610 219922 220678 219978
rect 220734 219922 220802 219978
rect 220858 219922 220926 219978
rect 220982 219922 251274 219978
rect 251330 219922 251398 219978
rect 251454 219922 251522 219978
rect 251578 219922 251646 219978
rect 251702 219922 272518 219978
rect 272574 219922 272642 219978
rect 272698 219922 303238 219978
rect 303294 219922 303362 219978
rect 303418 219922 343434 219978
rect 343490 219922 343558 219978
rect 343614 219922 343682 219978
rect 343738 219922 343806 219978
rect 343862 219922 374154 219978
rect 374210 219922 374278 219978
rect 374334 219922 374402 219978
rect 374458 219922 374526 219978
rect 374582 219922 404874 219978
rect 404930 219922 404998 219978
rect 405054 219922 405122 219978
rect 405178 219922 405246 219978
rect 405302 219922 435594 219978
rect 435650 219922 435718 219978
rect 435774 219922 435842 219978
rect 435898 219922 435966 219978
rect 436022 219922 466314 219978
rect 466370 219922 466438 219978
rect 466494 219922 466562 219978
rect 466618 219922 466686 219978
rect 466742 219922 497034 219978
rect 497090 219922 497158 219978
rect 497214 219922 497282 219978
rect 497338 219922 497406 219978
rect 497462 219922 527754 219978
rect 527810 219922 527878 219978
rect 527934 219922 528002 219978
rect 528058 219922 528126 219978
rect 528182 219922 558474 219978
rect 558530 219922 558598 219978
rect 558654 219922 558722 219978
rect 558778 219922 558846 219978
rect 558902 219922 589194 219978
rect 589250 219922 589318 219978
rect 589374 219922 589442 219978
rect 589498 219922 589566 219978
rect 589622 219922 596496 219978
rect 596552 219922 596620 219978
rect 596676 219922 596744 219978
rect 596800 219922 596868 219978
rect 596924 219922 597980 219978
rect -1916 219826 597980 219922
rect -1916 208350 597980 208446
rect -1916 208294 -1820 208350
rect -1764 208294 -1696 208350
rect -1640 208294 -1572 208350
rect -1516 208294 -1448 208350
rect -1392 208294 9234 208350
rect 9290 208294 9358 208350
rect 9414 208294 9482 208350
rect 9538 208294 9606 208350
rect 9662 208294 39878 208350
rect 39934 208294 40002 208350
rect 40058 208294 70674 208350
rect 70730 208294 70798 208350
rect 70854 208294 70922 208350
rect 70978 208294 71046 208350
rect 71102 208294 101878 208350
rect 101934 208294 102002 208350
rect 102058 208294 132114 208350
rect 132170 208294 132238 208350
rect 132294 208294 132362 208350
rect 132418 208294 132486 208350
rect 132542 208294 162834 208350
rect 162890 208294 162958 208350
rect 163014 208294 163082 208350
rect 163138 208294 163206 208350
rect 163262 208294 163878 208350
rect 163934 208294 164002 208350
rect 164058 208294 193554 208350
rect 193610 208294 193678 208350
rect 193734 208294 193802 208350
rect 193858 208294 193926 208350
rect 193982 208294 224274 208350
rect 224330 208294 224398 208350
rect 224454 208294 224522 208350
rect 224578 208294 224646 208350
rect 224702 208294 225878 208350
rect 225934 208294 226002 208350
rect 226058 208294 254994 208350
rect 255050 208294 255118 208350
rect 255174 208294 255242 208350
rect 255298 208294 255366 208350
rect 255422 208294 287878 208350
rect 287934 208294 288002 208350
rect 288058 208294 318598 208350
rect 318654 208294 318722 208350
rect 318778 208294 347154 208350
rect 347210 208294 347278 208350
rect 347334 208294 347402 208350
rect 347458 208294 347526 208350
rect 347582 208294 371878 208350
rect 371934 208294 372002 208350
rect 372058 208294 377874 208350
rect 377930 208294 377998 208350
rect 378054 208294 378122 208350
rect 378178 208294 378246 208350
rect 378302 208294 408594 208350
rect 408650 208294 408718 208350
rect 408774 208294 408842 208350
rect 408898 208294 408966 208350
rect 409022 208294 433878 208350
rect 433934 208294 434002 208350
rect 434058 208294 439314 208350
rect 439370 208294 439438 208350
rect 439494 208294 439562 208350
rect 439618 208294 439686 208350
rect 439742 208294 470034 208350
rect 470090 208294 470158 208350
rect 470214 208294 470282 208350
rect 470338 208294 470406 208350
rect 470462 208294 495878 208350
rect 495934 208294 496002 208350
rect 496058 208294 500754 208350
rect 500810 208294 500878 208350
rect 500934 208294 501002 208350
rect 501058 208294 501126 208350
rect 501182 208294 531474 208350
rect 531530 208294 531598 208350
rect 531654 208294 531722 208350
rect 531778 208294 531846 208350
rect 531902 208294 557878 208350
rect 557934 208294 558002 208350
rect 558058 208294 562194 208350
rect 562250 208294 562318 208350
rect 562374 208294 562442 208350
rect 562498 208294 562566 208350
rect 562622 208294 592914 208350
rect 592970 208294 593038 208350
rect 593094 208294 593162 208350
rect 593218 208294 593286 208350
rect 593342 208294 597456 208350
rect 597512 208294 597580 208350
rect 597636 208294 597704 208350
rect 597760 208294 597828 208350
rect 597884 208294 597980 208350
rect -1916 208226 597980 208294
rect -1916 208170 -1820 208226
rect -1764 208170 -1696 208226
rect -1640 208170 -1572 208226
rect -1516 208170 -1448 208226
rect -1392 208170 9234 208226
rect 9290 208170 9358 208226
rect 9414 208170 9482 208226
rect 9538 208170 9606 208226
rect 9662 208170 39878 208226
rect 39934 208170 40002 208226
rect 40058 208170 70674 208226
rect 70730 208170 70798 208226
rect 70854 208170 70922 208226
rect 70978 208170 71046 208226
rect 71102 208170 101878 208226
rect 101934 208170 102002 208226
rect 102058 208170 132114 208226
rect 132170 208170 132238 208226
rect 132294 208170 132362 208226
rect 132418 208170 132486 208226
rect 132542 208170 162834 208226
rect 162890 208170 162958 208226
rect 163014 208170 163082 208226
rect 163138 208170 163206 208226
rect 163262 208170 163878 208226
rect 163934 208170 164002 208226
rect 164058 208170 193554 208226
rect 193610 208170 193678 208226
rect 193734 208170 193802 208226
rect 193858 208170 193926 208226
rect 193982 208170 224274 208226
rect 224330 208170 224398 208226
rect 224454 208170 224522 208226
rect 224578 208170 224646 208226
rect 224702 208170 225878 208226
rect 225934 208170 226002 208226
rect 226058 208170 254994 208226
rect 255050 208170 255118 208226
rect 255174 208170 255242 208226
rect 255298 208170 255366 208226
rect 255422 208170 287878 208226
rect 287934 208170 288002 208226
rect 288058 208170 318598 208226
rect 318654 208170 318722 208226
rect 318778 208170 347154 208226
rect 347210 208170 347278 208226
rect 347334 208170 347402 208226
rect 347458 208170 347526 208226
rect 347582 208170 371878 208226
rect 371934 208170 372002 208226
rect 372058 208170 377874 208226
rect 377930 208170 377998 208226
rect 378054 208170 378122 208226
rect 378178 208170 378246 208226
rect 378302 208170 408594 208226
rect 408650 208170 408718 208226
rect 408774 208170 408842 208226
rect 408898 208170 408966 208226
rect 409022 208170 433878 208226
rect 433934 208170 434002 208226
rect 434058 208170 439314 208226
rect 439370 208170 439438 208226
rect 439494 208170 439562 208226
rect 439618 208170 439686 208226
rect 439742 208170 470034 208226
rect 470090 208170 470158 208226
rect 470214 208170 470282 208226
rect 470338 208170 470406 208226
rect 470462 208170 495878 208226
rect 495934 208170 496002 208226
rect 496058 208170 500754 208226
rect 500810 208170 500878 208226
rect 500934 208170 501002 208226
rect 501058 208170 501126 208226
rect 501182 208170 531474 208226
rect 531530 208170 531598 208226
rect 531654 208170 531722 208226
rect 531778 208170 531846 208226
rect 531902 208170 557878 208226
rect 557934 208170 558002 208226
rect 558058 208170 562194 208226
rect 562250 208170 562318 208226
rect 562374 208170 562442 208226
rect 562498 208170 562566 208226
rect 562622 208170 592914 208226
rect 592970 208170 593038 208226
rect 593094 208170 593162 208226
rect 593218 208170 593286 208226
rect 593342 208170 597456 208226
rect 597512 208170 597580 208226
rect 597636 208170 597704 208226
rect 597760 208170 597828 208226
rect 597884 208170 597980 208226
rect -1916 208102 597980 208170
rect -1916 208046 -1820 208102
rect -1764 208046 -1696 208102
rect -1640 208046 -1572 208102
rect -1516 208046 -1448 208102
rect -1392 208046 9234 208102
rect 9290 208046 9358 208102
rect 9414 208046 9482 208102
rect 9538 208046 9606 208102
rect 9662 208046 39878 208102
rect 39934 208046 40002 208102
rect 40058 208046 70674 208102
rect 70730 208046 70798 208102
rect 70854 208046 70922 208102
rect 70978 208046 71046 208102
rect 71102 208046 101878 208102
rect 101934 208046 102002 208102
rect 102058 208046 132114 208102
rect 132170 208046 132238 208102
rect 132294 208046 132362 208102
rect 132418 208046 132486 208102
rect 132542 208046 162834 208102
rect 162890 208046 162958 208102
rect 163014 208046 163082 208102
rect 163138 208046 163206 208102
rect 163262 208046 163878 208102
rect 163934 208046 164002 208102
rect 164058 208046 193554 208102
rect 193610 208046 193678 208102
rect 193734 208046 193802 208102
rect 193858 208046 193926 208102
rect 193982 208046 224274 208102
rect 224330 208046 224398 208102
rect 224454 208046 224522 208102
rect 224578 208046 224646 208102
rect 224702 208046 225878 208102
rect 225934 208046 226002 208102
rect 226058 208046 254994 208102
rect 255050 208046 255118 208102
rect 255174 208046 255242 208102
rect 255298 208046 255366 208102
rect 255422 208046 287878 208102
rect 287934 208046 288002 208102
rect 288058 208046 318598 208102
rect 318654 208046 318722 208102
rect 318778 208046 347154 208102
rect 347210 208046 347278 208102
rect 347334 208046 347402 208102
rect 347458 208046 347526 208102
rect 347582 208046 371878 208102
rect 371934 208046 372002 208102
rect 372058 208046 377874 208102
rect 377930 208046 377998 208102
rect 378054 208046 378122 208102
rect 378178 208046 378246 208102
rect 378302 208046 408594 208102
rect 408650 208046 408718 208102
rect 408774 208046 408842 208102
rect 408898 208046 408966 208102
rect 409022 208046 433878 208102
rect 433934 208046 434002 208102
rect 434058 208046 439314 208102
rect 439370 208046 439438 208102
rect 439494 208046 439562 208102
rect 439618 208046 439686 208102
rect 439742 208046 470034 208102
rect 470090 208046 470158 208102
rect 470214 208046 470282 208102
rect 470338 208046 470406 208102
rect 470462 208046 495878 208102
rect 495934 208046 496002 208102
rect 496058 208046 500754 208102
rect 500810 208046 500878 208102
rect 500934 208046 501002 208102
rect 501058 208046 501126 208102
rect 501182 208046 531474 208102
rect 531530 208046 531598 208102
rect 531654 208046 531722 208102
rect 531778 208046 531846 208102
rect 531902 208046 557878 208102
rect 557934 208046 558002 208102
rect 558058 208046 562194 208102
rect 562250 208046 562318 208102
rect 562374 208046 562442 208102
rect 562498 208046 562566 208102
rect 562622 208046 592914 208102
rect 592970 208046 593038 208102
rect 593094 208046 593162 208102
rect 593218 208046 593286 208102
rect 593342 208046 597456 208102
rect 597512 208046 597580 208102
rect 597636 208046 597704 208102
rect 597760 208046 597828 208102
rect 597884 208046 597980 208102
rect -1916 207978 597980 208046
rect -1916 207922 -1820 207978
rect -1764 207922 -1696 207978
rect -1640 207922 -1572 207978
rect -1516 207922 -1448 207978
rect -1392 207922 9234 207978
rect 9290 207922 9358 207978
rect 9414 207922 9482 207978
rect 9538 207922 9606 207978
rect 9662 207922 39878 207978
rect 39934 207922 40002 207978
rect 40058 207922 70674 207978
rect 70730 207922 70798 207978
rect 70854 207922 70922 207978
rect 70978 207922 71046 207978
rect 71102 207922 101878 207978
rect 101934 207922 102002 207978
rect 102058 207922 132114 207978
rect 132170 207922 132238 207978
rect 132294 207922 132362 207978
rect 132418 207922 132486 207978
rect 132542 207922 162834 207978
rect 162890 207922 162958 207978
rect 163014 207922 163082 207978
rect 163138 207922 163206 207978
rect 163262 207922 163878 207978
rect 163934 207922 164002 207978
rect 164058 207922 193554 207978
rect 193610 207922 193678 207978
rect 193734 207922 193802 207978
rect 193858 207922 193926 207978
rect 193982 207922 224274 207978
rect 224330 207922 224398 207978
rect 224454 207922 224522 207978
rect 224578 207922 224646 207978
rect 224702 207922 225878 207978
rect 225934 207922 226002 207978
rect 226058 207922 254994 207978
rect 255050 207922 255118 207978
rect 255174 207922 255242 207978
rect 255298 207922 255366 207978
rect 255422 207922 287878 207978
rect 287934 207922 288002 207978
rect 288058 207922 318598 207978
rect 318654 207922 318722 207978
rect 318778 207922 347154 207978
rect 347210 207922 347278 207978
rect 347334 207922 347402 207978
rect 347458 207922 347526 207978
rect 347582 207922 371878 207978
rect 371934 207922 372002 207978
rect 372058 207922 377874 207978
rect 377930 207922 377998 207978
rect 378054 207922 378122 207978
rect 378178 207922 378246 207978
rect 378302 207922 408594 207978
rect 408650 207922 408718 207978
rect 408774 207922 408842 207978
rect 408898 207922 408966 207978
rect 409022 207922 433878 207978
rect 433934 207922 434002 207978
rect 434058 207922 439314 207978
rect 439370 207922 439438 207978
rect 439494 207922 439562 207978
rect 439618 207922 439686 207978
rect 439742 207922 470034 207978
rect 470090 207922 470158 207978
rect 470214 207922 470282 207978
rect 470338 207922 470406 207978
rect 470462 207922 495878 207978
rect 495934 207922 496002 207978
rect 496058 207922 500754 207978
rect 500810 207922 500878 207978
rect 500934 207922 501002 207978
rect 501058 207922 501126 207978
rect 501182 207922 531474 207978
rect 531530 207922 531598 207978
rect 531654 207922 531722 207978
rect 531778 207922 531846 207978
rect 531902 207922 557878 207978
rect 557934 207922 558002 207978
rect 558058 207922 562194 207978
rect 562250 207922 562318 207978
rect 562374 207922 562442 207978
rect 562498 207922 562566 207978
rect 562622 207922 592914 207978
rect 592970 207922 593038 207978
rect 593094 207922 593162 207978
rect 593218 207922 593286 207978
rect 593342 207922 597456 207978
rect 597512 207922 597580 207978
rect 597636 207922 597704 207978
rect 597760 207922 597828 207978
rect 597884 207922 597980 207978
rect -1916 207826 597980 207922
rect 202956 205858 262180 205874
rect 202956 205802 202972 205858
rect 203028 205802 262108 205858
rect 262164 205802 262180 205858
rect 202956 205786 262180 205802
rect 334444 205138 526724 205154
rect 334444 205082 334460 205138
rect 334516 205082 526652 205138
rect 526708 205082 526724 205138
rect 334444 205066 526724 205082
rect 334444 203338 525044 203354
rect 334444 203282 334460 203338
rect 334516 203282 524972 203338
rect 525028 203282 525044 203338
rect 334444 203266 525044 203282
rect -1916 202350 597980 202446
rect -1916 202294 -860 202350
rect -804 202294 -736 202350
rect -680 202294 -612 202350
rect -556 202294 -488 202350
rect -432 202294 5514 202350
rect 5570 202294 5638 202350
rect 5694 202294 5762 202350
rect 5818 202294 5886 202350
rect 5942 202294 24518 202350
rect 24574 202294 24642 202350
rect 24698 202294 36234 202350
rect 36290 202294 36358 202350
rect 36414 202294 36482 202350
rect 36538 202294 36606 202350
rect 36662 202294 55238 202350
rect 55294 202294 55362 202350
rect 55418 202294 66954 202350
rect 67010 202294 67078 202350
rect 67134 202294 67202 202350
rect 67258 202294 67326 202350
rect 67382 202294 86518 202350
rect 86574 202294 86642 202350
rect 86698 202294 97674 202350
rect 97730 202294 97798 202350
rect 97854 202294 97922 202350
rect 97978 202294 98046 202350
rect 98102 202294 117238 202350
rect 117294 202294 117362 202350
rect 117418 202294 128394 202350
rect 128450 202294 128518 202350
rect 128574 202294 128642 202350
rect 128698 202294 128766 202350
rect 128822 202294 148518 202350
rect 148574 202294 148642 202350
rect 148698 202294 159114 202350
rect 159170 202294 159238 202350
rect 159294 202294 159362 202350
rect 159418 202294 159486 202350
rect 159542 202294 179238 202350
rect 179294 202294 179362 202350
rect 179418 202294 189834 202350
rect 189890 202294 189958 202350
rect 190014 202294 190082 202350
rect 190138 202294 190206 202350
rect 190262 202294 210518 202350
rect 210574 202294 210642 202350
rect 210698 202294 220554 202350
rect 220610 202294 220678 202350
rect 220734 202294 220802 202350
rect 220858 202294 220926 202350
rect 220982 202294 241238 202350
rect 241294 202294 241362 202350
rect 241418 202294 251274 202350
rect 251330 202294 251398 202350
rect 251454 202294 251522 202350
rect 251578 202294 251646 202350
rect 251702 202294 272518 202350
rect 272574 202294 272642 202350
rect 272698 202294 303238 202350
rect 303294 202294 303362 202350
rect 303418 202294 343434 202350
rect 343490 202294 343558 202350
rect 343614 202294 343682 202350
rect 343738 202294 343806 202350
rect 343862 202294 356518 202350
rect 356574 202294 356642 202350
rect 356698 202294 374154 202350
rect 374210 202294 374278 202350
rect 374334 202294 374402 202350
rect 374458 202294 374526 202350
rect 374582 202294 387238 202350
rect 387294 202294 387362 202350
rect 387418 202294 404874 202350
rect 404930 202294 404998 202350
rect 405054 202294 405122 202350
rect 405178 202294 405246 202350
rect 405302 202294 418518 202350
rect 418574 202294 418642 202350
rect 418698 202294 435594 202350
rect 435650 202294 435718 202350
rect 435774 202294 435842 202350
rect 435898 202294 435966 202350
rect 436022 202294 449238 202350
rect 449294 202294 449362 202350
rect 449418 202294 466314 202350
rect 466370 202294 466438 202350
rect 466494 202294 466562 202350
rect 466618 202294 466686 202350
rect 466742 202294 480518 202350
rect 480574 202294 480642 202350
rect 480698 202294 497034 202350
rect 497090 202294 497158 202350
rect 497214 202294 497282 202350
rect 497338 202294 497406 202350
rect 497462 202294 511238 202350
rect 511294 202294 511362 202350
rect 511418 202294 527754 202350
rect 527810 202294 527878 202350
rect 527934 202294 528002 202350
rect 528058 202294 528126 202350
rect 528182 202294 542518 202350
rect 542574 202294 542642 202350
rect 542698 202294 558474 202350
rect 558530 202294 558598 202350
rect 558654 202294 558722 202350
rect 558778 202294 558846 202350
rect 558902 202294 573238 202350
rect 573294 202294 573362 202350
rect 573418 202294 589194 202350
rect 589250 202294 589318 202350
rect 589374 202294 589442 202350
rect 589498 202294 589566 202350
rect 589622 202294 596496 202350
rect 596552 202294 596620 202350
rect 596676 202294 596744 202350
rect 596800 202294 596868 202350
rect 596924 202294 597980 202350
rect -1916 202226 597980 202294
rect -1916 202170 -860 202226
rect -804 202170 -736 202226
rect -680 202170 -612 202226
rect -556 202170 -488 202226
rect -432 202170 5514 202226
rect 5570 202170 5638 202226
rect 5694 202170 5762 202226
rect 5818 202170 5886 202226
rect 5942 202170 24518 202226
rect 24574 202170 24642 202226
rect 24698 202170 36234 202226
rect 36290 202170 36358 202226
rect 36414 202170 36482 202226
rect 36538 202170 36606 202226
rect 36662 202170 55238 202226
rect 55294 202170 55362 202226
rect 55418 202170 66954 202226
rect 67010 202170 67078 202226
rect 67134 202170 67202 202226
rect 67258 202170 67326 202226
rect 67382 202170 86518 202226
rect 86574 202170 86642 202226
rect 86698 202170 97674 202226
rect 97730 202170 97798 202226
rect 97854 202170 97922 202226
rect 97978 202170 98046 202226
rect 98102 202170 117238 202226
rect 117294 202170 117362 202226
rect 117418 202170 128394 202226
rect 128450 202170 128518 202226
rect 128574 202170 128642 202226
rect 128698 202170 128766 202226
rect 128822 202170 148518 202226
rect 148574 202170 148642 202226
rect 148698 202170 159114 202226
rect 159170 202170 159238 202226
rect 159294 202170 159362 202226
rect 159418 202170 159486 202226
rect 159542 202170 179238 202226
rect 179294 202170 179362 202226
rect 179418 202170 189834 202226
rect 189890 202170 189958 202226
rect 190014 202170 190082 202226
rect 190138 202170 190206 202226
rect 190262 202170 210518 202226
rect 210574 202170 210642 202226
rect 210698 202170 220554 202226
rect 220610 202170 220678 202226
rect 220734 202170 220802 202226
rect 220858 202170 220926 202226
rect 220982 202170 241238 202226
rect 241294 202170 241362 202226
rect 241418 202170 251274 202226
rect 251330 202170 251398 202226
rect 251454 202170 251522 202226
rect 251578 202170 251646 202226
rect 251702 202170 272518 202226
rect 272574 202170 272642 202226
rect 272698 202170 303238 202226
rect 303294 202170 303362 202226
rect 303418 202170 343434 202226
rect 343490 202170 343558 202226
rect 343614 202170 343682 202226
rect 343738 202170 343806 202226
rect 343862 202170 356518 202226
rect 356574 202170 356642 202226
rect 356698 202170 374154 202226
rect 374210 202170 374278 202226
rect 374334 202170 374402 202226
rect 374458 202170 374526 202226
rect 374582 202170 387238 202226
rect 387294 202170 387362 202226
rect 387418 202170 404874 202226
rect 404930 202170 404998 202226
rect 405054 202170 405122 202226
rect 405178 202170 405246 202226
rect 405302 202170 418518 202226
rect 418574 202170 418642 202226
rect 418698 202170 435594 202226
rect 435650 202170 435718 202226
rect 435774 202170 435842 202226
rect 435898 202170 435966 202226
rect 436022 202170 449238 202226
rect 449294 202170 449362 202226
rect 449418 202170 466314 202226
rect 466370 202170 466438 202226
rect 466494 202170 466562 202226
rect 466618 202170 466686 202226
rect 466742 202170 480518 202226
rect 480574 202170 480642 202226
rect 480698 202170 497034 202226
rect 497090 202170 497158 202226
rect 497214 202170 497282 202226
rect 497338 202170 497406 202226
rect 497462 202170 511238 202226
rect 511294 202170 511362 202226
rect 511418 202170 527754 202226
rect 527810 202170 527878 202226
rect 527934 202170 528002 202226
rect 528058 202170 528126 202226
rect 528182 202170 542518 202226
rect 542574 202170 542642 202226
rect 542698 202170 558474 202226
rect 558530 202170 558598 202226
rect 558654 202170 558722 202226
rect 558778 202170 558846 202226
rect 558902 202170 573238 202226
rect 573294 202170 573362 202226
rect 573418 202170 589194 202226
rect 589250 202170 589318 202226
rect 589374 202170 589442 202226
rect 589498 202170 589566 202226
rect 589622 202170 596496 202226
rect 596552 202170 596620 202226
rect 596676 202170 596744 202226
rect 596800 202170 596868 202226
rect 596924 202170 597980 202226
rect -1916 202102 597980 202170
rect -1916 202046 -860 202102
rect -804 202046 -736 202102
rect -680 202046 -612 202102
rect -556 202046 -488 202102
rect -432 202046 5514 202102
rect 5570 202046 5638 202102
rect 5694 202046 5762 202102
rect 5818 202046 5886 202102
rect 5942 202046 24518 202102
rect 24574 202046 24642 202102
rect 24698 202046 36234 202102
rect 36290 202046 36358 202102
rect 36414 202046 36482 202102
rect 36538 202046 36606 202102
rect 36662 202046 55238 202102
rect 55294 202046 55362 202102
rect 55418 202046 66954 202102
rect 67010 202046 67078 202102
rect 67134 202046 67202 202102
rect 67258 202046 67326 202102
rect 67382 202046 86518 202102
rect 86574 202046 86642 202102
rect 86698 202046 97674 202102
rect 97730 202046 97798 202102
rect 97854 202046 97922 202102
rect 97978 202046 98046 202102
rect 98102 202046 117238 202102
rect 117294 202046 117362 202102
rect 117418 202046 128394 202102
rect 128450 202046 128518 202102
rect 128574 202046 128642 202102
rect 128698 202046 128766 202102
rect 128822 202046 148518 202102
rect 148574 202046 148642 202102
rect 148698 202046 159114 202102
rect 159170 202046 159238 202102
rect 159294 202046 159362 202102
rect 159418 202046 159486 202102
rect 159542 202046 179238 202102
rect 179294 202046 179362 202102
rect 179418 202046 189834 202102
rect 189890 202046 189958 202102
rect 190014 202046 190082 202102
rect 190138 202046 190206 202102
rect 190262 202046 210518 202102
rect 210574 202046 210642 202102
rect 210698 202046 220554 202102
rect 220610 202046 220678 202102
rect 220734 202046 220802 202102
rect 220858 202046 220926 202102
rect 220982 202046 241238 202102
rect 241294 202046 241362 202102
rect 241418 202046 251274 202102
rect 251330 202046 251398 202102
rect 251454 202046 251522 202102
rect 251578 202046 251646 202102
rect 251702 202046 272518 202102
rect 272574 202046 272642 202102
rect 272698 202046 303238 202102
rect 303294 202046 303362 202102
rect 303418 202046 343434 202102
rect 343490 202046 343558 202102
rect 343614 202046 343682 202102
rect 343738 202046 343806 202102
rect 343862 202046 356518 202102
rect 356574 202046 356642 202102
rect 356698 202046 374154 202102
rect 374210 202046 374278 202102
rect 374334 202046 374402 202102
rect 374458 202046 374526 202102
rect 374582 202046 387238 202102
rect 387294 202046 387362 202102
rect 387418 202046 404874 202102
rect 404930 202046 404998 202102
rect 405054 202046 405122 202102
rect 405178 202046 405246 202102
rect 405302 202046 418518 202102
rect 418574 202046 418642 202102
rect 418698 202046 435594 202102
rect 435650 202046 435718 202102
rect 435774 202046 435842 202102
rect 435898 202046 435966 202102
rect 436022 202046 449238 202102
rect 449294 202046 449362 202102
rect 449418 202046 466314 202102
rect 466370 202046 466438 202102
rect 466494 202046 466562 202102
rect 466618 202046 466686 202102
rect 466742 202046 480518 202102
rect 480574 202046 480642 202102
rect 480698 202046 497034 202102
rect 497090 202046 497158 202102
rect 497214 202046 497282 202102
rect 497338 202046 497406 202102
rect 497462 202046 511238 202102
rect 511294 202046 511362 202102
rect 511418 202046 527754 202102
rect 527810 202046 527878 202102
rect 527934 202046 528002 202102
rect 528058 202046 528126 202102
rect 528182 202046 542518 202102
rect 542574 202046 542642 202102
rect 542698 202046 558474 202102
rect 558530 202046 558598 202102
rect 558654 202046 558722 202102
rect 558778 202046 558846 202102
rect 558902 202046 573238 202102
rect 573294 202046 573362 202102
rect 573418 202046 589194 202102
rect 589250 202046 589318 202102
rect 589374 202046 589442 202102
rect 589498 202046 589566 202102
rect 589622 202046 596496 202102
rect 596552 202046 596620 202102
rect 596676 202046 596744 202102
rect 596800 202046 596868 202102
rect 596924 202046 597980 202102
rect -1916 201978 597980 202046
rect -1916 201922 -860 201978
rect -804 201922 -736 201978
rect -680 201922 -612 201978
rect -556 201922 -488 201978
rect -432 201922 5514 201978
rect 5570 201922 5638 201978
rect 5694 201922 5762 201978
rect 5818 201922 5886 201978
rect 5942 201922 24518 201978
rect 24574 201922 24642 201978
rect 24698 201922 36234 201978
rect 36290 201922 36358 201978
rect 36414 201922 36482 201978
rect 36538 201922 36606 201978
rect 36662 201922 55238 201978
rect 55294 201922 55362 201978
rect 55418 201922 66954 201978
rect 67010 201922 67078 201978
rect 67134 201922 67202 201978
rect 67258 201922 67326 201978
rect 67382 201922 86518 201978
rect 86574 201922 86642 201978
rect 86698 201922 97674 201978
rect 97730 201922 97798 201978
rect 97854 201922 97922 201978
rect 97978 201922 98046 201978
rect 98102 201922 117238 201978
rect 117294 201922 117362 201978
rect 117418 201922 128394 201978
rect 128450 201922 128518 201978
rect 128574 201922 128642 201978
rect 128698 201922 128766 201978
rect 128822 201922 148518 201978
rect 148574 201922 148642 201978
rect 148698 201922 159114 201978
rect 159170 201922 159238 201978
rect 159294 201922 159362 201978
rect 159418 201922 159486 201978
rect 159542 201922 179238 201978
rect 179294 201922 179362 201978
rect 179418 201922 189834 201978
rect 189890 201922 189958 201978
rect 190014 201922 190082 201978
rect 190138 201922 190206 201978
rect 190262 201922 210518 201978
rect 210574 201922 210642 201978
rect 210698 201922 220554 201978
rect 220610 201922 220678 201978
rect 220734 201922 220802 201978
rect 220858 201922 220926 201978
rect 220982 201922 241238 201978
rect 241294 201922 241362 201978
rect 241418 201922 251274 201978
rect 251330 201922 251398 201978
rect 251454 201922 251522 201978
rect 251578 201922 251646 201978
rect 251702 201922 272518 201978
rect 272574 201922 272642 201978
rect 272698 201922 303238 201978
rect 303294 201922 303362 201978
rect 303418 201922 343434 201978
rect 343490 201922 343558 201978
rect 343614 201922 343682 201978
rect 343738 201922 343806 201978
rect 343862 201922 356518 201978
rect 356574 201922 356642 201978
rect 356698 201922 374154 201978
rect 374210 201922 374278 201978
rect 374334 201922 374402 201978
rect 374458 201922 374526 201978
rect 374582 201922 387238 201978
rect 387294 201922 387362 201978
rect 387418 201922 404874 201978
rect 404930 201922 404998 201978
rect 405054 201922 405122 201978
rect 405178 201922 405246 201978
rect 405302 201922 418518 201978
rect 418574 201922 418642 201978
rect 418698 201922 435594 201978
rect 435650 201922 435718 201978
rect 435774 201922 435842 201978
rect 435898 201922 435966 201978
rect 436022 201922 449238 201978
rect 449294 201922 449362 201978
rect 449418 201922 466314 201978
rect 466370 201922 466438 201978
rect 466494 201922 466562 201978
rect 466618 201922 466686 201978
rect 466742 201922 480518 201978
rect 480574 201922 480642 201978
rect 480698 201922 497034 201978
rect 497090 201922 497158 201978
rect 497214 201922 497282 201978
rect 497338 201922 497406 201978
rect 497462 201922 511238 201978
rect 511294 201922 511362 201978
rect 511418 201922 527754 201978
rect 527810 201922 527878 201978
rect 527934 201922 528002 201978
rect 528058 201922 528126 201978
rect 528182 201922 542518 201978
rect 542574 201922 542642 201978
rect 542698 201922 558474 201978
rect 558530 201922 558598 201978
rect 558654 201922 558722 201978
rect 558778 201922 558846 201978
rect 558902 201922 573238 201978
rect 573294 201922 573362 201978
rect 573418 201922 589194 201978
rect 589250 201922 589318 201978
rect 589374 201922 589442 201978
rect 589498 201922 589566 201978
rect 589622 201922 596496 201978
rect 596552 201922 596620 201978
rect 596676 201922 596744 201978
rect 596800 201922 596868 201978
rect 596924 201922 597980 201978
rect -1916 201826 597980 201922
rect 334444 200818 519220 200834
rect 334444 200762 334460 200818
rect 334516 200762 519148 200818
rect 519204 200762 519220 200818
rect 334444 200746 519220 200762
rect 334444 200098 467924 200114
rect 334444 200042 334460 200098
rect 334516 200042 467852 200098
rect 467908 200042 467924 200098
rect 334444 200026 467924 200042
rect 18380 199018 201700 199034
rect 18380 198962 18396 199018
rect 18452 198962 82684 199018
rect 82740 198962 141036 199018
rect 141092 198962 201628 199018
rect 201684 198962 201700 199018
rect 18380 198946 201700 198962
rect 352700 199018 402404 199034
rect 352700 198962 352716 199018
rect 352772 198962 402404 199018
rect 352700 198946 402404 198962
rect 402316 198314 402404 198946
rect 403100 198478 455380 198494
rect 403100 198422 403116 198478
rect 403172 198422 455308 198478
rect 455364 198422 455380 198478
rect 403100 198406 455380 198422
rect 205644 198298 263860 198314
rect 205644 198242 205660 198298
rect 205716 198242 263788 198298
rect 263844 198242 263860 198298
rect 205644 198226 263860 198242
rect 334444 198298 401508 198314
rect 334444 198242 334460 198298
rect 334516 198242 401436 198298
rect 401492 198242 401508 198298
rect 334444 198226 401508 198242
rect 402316 198298 534340 198314
rect 402316 198242 414652 198298
rect 414708 198242 473676 198298
rect 473732 198242 534268 198298
rect 534324 198242 534340 198298
rect 402316 198226 534340 198242
rect 196572 196858 263860 196874
rect 196572 196802 196588 196858
rect 196644 196802 263788 196858
rect 263844 196802 263860 196858
rect 196572 196786 263860 196802
rect 334444 196858 456164 196874
rect 334444 196802 334460 196858
rect 334516 196802 456092 196858
rect 456148 196802 456164 196858
rect 334444 196786 456164 196802
rect 64188 196678 187364 196694
rect 64188 196622 64204 196678
rect 64260 196622 187292 196678
rect 187348 196622 187364 196678
rect 64188 196606 187364 196622
rect 197468 196678 263972 196694
rect 197468 196622 197484 196678
rect 197540 196622 263900 196678
rect 263956 196622 263972 196678
rect 197468 196606 263972 196622
rect 334444 196678 463668 196694
rect 334444 196622 334460 196678
rect 334516 196622 463596 196678
rect 463652 196622 463668 196678
rect 334444 196606 463668 196622
rect 189516 196498 248628 196514
rect 189516 196442 189532 196498
rect 189588 196442 248556 196498
rect 248612 196442 248628 196498
rect 189516 196426 248628 196442
rect 401420 195778 472180 195794
rect 401420 195722 401436 195778
rect 401492 195722 472108 195778
rect 472164 195722 472180 195778
rect 401420 195706 472180 195722
rect 64188 195238 188148 195254
rect 64188 195182 64204 195238
rect 64260 195182 188076 195238
rect 188132 195182 188148 195238
rect 64188 195166 188148 195182
rect 351804 195238 411252 195254
rect 351804 195182 351820 195238
rect 351876 195182 411180 195238
rect 411236 195182 411252 195238
rect 351804 195166 411252 195182
rect 20620 195058 191620 195074
rect 20620 195002 20636 195058
rect 20692 195002 191548 195058
rect 191604 195002 191620 195058
rect 20620 194986 191620 195002
rect 204972 195058 263860 195074
rect 204972 195002 204988 195058
rect 205044 195002 263788 195058
rect 263844 195002 263860 195058
rect 204972 194986 263860 195002
rect 334444 195058 403300 195074
rect 334444 195002 334460 195058
rect 334516 195002 403228 195058
rect 403284 195002 403300 195058
rect 334444 194986 403300 195002
rect 334444 194878 403188 194894
rect 334444 194822 334460 194878
rect 334516 194822 403116 194878
rect 403172 194822 403188 194878
rect 334444 194806 403188 194822
rect 20284 194158 248628 194174
rect 20284 194102 20300 194158
rect 20356 194102 248556 194158
rect 248612 194102 248628 194158
rect 20284 194086 248628 194102
rect 127468 193978 169780 193994
rect 127468 193922 127484 193978
rect 127540 193922 169708 193978
rect 169764 193922 169780 193978
rect 127468 193906 169780 193922
rect 334444 193978 455380 193994
rect 334444 193922 334460 193978
rect 334516 193922 455308 193978
rect 455364 193922 455380 193978
rect 334444 193906 455380 193922
rect 127580 193258 262180 193274
rect 127580 193202 127596 193258
rect 127652 193202 262108 193258
rect 262164 193202 262180 193258
rect 127580 193186 262180 193202
rect 334444 193258 401508 193274
rect 334444 193202 334460 193258
rect 334516 193202 401508 193258
rect 334444 193186 401508 193202
rect 401420 193094 401508 193186
rect 401420 193006 408284 193094
rect 408196 192734 408284 193006
rect 408196 192646 455492 192734
rect 347772 192538 411364 192554
rect 347772 192482 347788 192538
rect 347844 192482 411292 192538
rect 411348 192482 411364 192538
rect 347772 192466 411364 192482
rect 334444 192358 411252 192374
rect 334444 192302 334460 192358
rect 334516 192302 411180 192358
rect 411236 192302 411252 192358
rect 334444 192286 411252 192302
rect 134412 192178 263860 192194
rect 134412 192122 134428 192178
rect 134484 192122 263788 192178
rect 263844 192122 263860 192178
rect 134412 192106 263860 192122
rect 455404 192178 455492 192646
rect 526636 192358 579812 192374
rect 526636 192302 526652 192358
rect 526708 192302 579812 192358
rect 526636 192286 579812 192302
rect 455404 192122 455420 192178
rect 455476 192122 455492 192178
rect 455404 192106 455492 192122
rect 579724 192178 579812 192286
rect 579724 192122 579740 192178
rect 579796 192122 579812 192178
rect 579724 192106 579812 192122
rect -1916 190350 597980 190446
rect -1916 190294 -1820 190350
rect -1764 190294 -1696 190350
rect -1640 190294 -1572 190350
rect -1516 190294 -1448 190350
rect -1392 190294 9234 190350
rect 9290 190294 9358 190350
rect 9414 190294 9482 190350
rect 9538 190294 9606 190350
rect 9662 190294 39878 190350
rect 39934 190294 40002 190350
rect 40058 190294 70674 190350
rect 70730 190294 70798 190350
rect 70854 190294 70922 190350
rect 70978 190294 71046 190350
rect 71102 190294 101878 190350
rect 101934 190294 102002 190350
rect 102058 190294 132114 190350
rect 132170 190294 132238 190350
rect 132294 190294 132362 190350
rect 132418 190294 132486 190350
rect 132542 190294 163878 190350
rect 163934 190294 164002 190350
rect 164058 190294 193554 190350
rect 193610 190294 193678 190350
rect 193734 190294 193802 190350
rect 193858 190294 193926 190350
rect 193982 190294 224274 190350
rect 224330 190294 224398 190350
rect 224454 190294 224522 190350
rect 224578 190294 224646 190350
rect 224702 190294 225878 190350
rect 225934 190294 226002 190350
rect 226058 190294 254994 190350
rect 255050 190294 255118 190350
rect 255174 190294 255242 190350
rect 255298 190294 255366 190350
rect 255422 190294 287878 190350
rect 287934 190294 288002 190350
rect 288058 190294 318598 190350
rect 318654 190294 318722 190350
rect 318778 190294 347154 190350
rect 347210 190294 347278 190350
rect 347334 190294 347402 190350
rect 347458 190294 347526 190350
rect 347582 190294 371878 190350
rect 371934 190294 372002 190350
rect 372058 190294 377874 190350
rect 377930 190294 377998 190350
rect 378054 190294 378122 190350
rect 378178 190294 378246 190350
rect 378302 190294 408594 190350
rect 408650 190294 408718 190350
rect 408774 190294 408842 190350
rect 408898 190294 408966 190350
rect 409022 190294 433878 190350
rect 433934 190294 434002 190350
rect 434058 190294 439314 190350
rect 439370 190294 439438 190350
rect 439494 190294 439562 190350
rect 439618 190294 439686 190350
rect 439742 190294 470034 190350
rect 470090 190294 470158 190350
rect 470214 190294 470282 190350
rect 470338 190294 470406 190350
rect 470462 190294 495878 190350
rect 495934 190294 496002 190350
rect 496058 190294 500754 190350
rect 500810 190294 500878 190350
rect 500934 190294 501002 190350
rect 501058 190294 501126 190350
rect 501182 190294 531474 190350
rect 531530 190294 531598 190350
rect 531654 190294 531722 190350
rect 531778 190294 531846 190350
rect 531902 190294 557878 190350
rect 557934 190294 558002 190350
rect 558058 190294 562194 190350
rect 562250 190294 562318 190350
rect 562374 190294 562442 190350
rect 562498 190294 562566 190350
rect 562622 190294 592914 190350
rect 592970 190294 593038 190350
rect 593094 190294 593162 190350
rect 593218 190294 593286 190350
rect 593342 190294 597456 190350
rect 597512 190294 597580 190350
rect 597636 190294 597704 190350
rect 597760 190294 597828 190350
rect 597884 190294 597980 190350
rect -1916 190226 597980 190294
rect -1916 190170 -1820 190226
rect -1764 190170 -1696 190226
rect -1640 190170 -1572 190226
rect -1516 190170 -1448 190226
rect -1392 190170 9234 190226
rect 9290 190170 9358 190226
rect 9414 190170 9482 190226
rect 9538 190170 9606 190226
rect 9662 190170 39878 190226
rect 39934 190170 40002 190226
rect 40058 190170 70674 190226
rect 70730 190170 70798 190226
rect 70854 190170 70922 190226
rect 70978 190170 71046 190226
rect 71102 190170 101878 190226
rect 101934 190170 102002 190226
rect 102058 190170 132114 190226
rect 132170 190170 132238 190226
rect 132294 190170 132362 190226
rect 132418 190170 132486 190226
rect 132542 190170 163878 190226
rect 163934 190170 164002 190226
rect 164058 190170 193554 190226
rect 193610 190170 193678 190226
rect 193734 190170 193802 190226
rect 193858 190170 193926 190226
rect 193982 190170 224274 190226
rect 224330 190170 224398 190226
rect 224454 190170 224522 190226
rect 224578 190170 224646 190226
rect 224702 190170 225878 190226
rect 225934 190170 226002 190226
rect 226058 190170 254994 190226
rect 255050 190170 255118 190226
rect 255174 190170 255242 190226
rect 255298 190170 255366 190226
rect 255422 190170 287878 190226
rect 287934 190170 288002 190226
rect 288058 190170 318598 190226
rect 318654 190170 318722 190226
rect 318778 190170 347154 190226
rect 347210 190170 347278 190226
rect 347334 190170 347402 190226
rect 347458 190170 347526 190226
rect 347582 190170 371878 190226
rect 371934 190170 372002 190226
rect 372058 190170 377874 190226
rect 377930 190170 377998 190226
rect 378054 190170 378122 190226
rect 378178 190170 378246 190226
rect 378302 190170 408594 190226
rect 408650 190170 408718 190226
rect 408774 190170 408842 190226
rect 408898 190170 408966 190226
rect 409022 190170 433878 190226
rect 433934 190170 434002 190226
rect 434058 190170 439314 190226
rect 439370 190170 439438 190226
rect 439494 190170 439562 190226
rect 439618 190170 439686 190226
rect 439742 190170 470034 190226
rect 470090 190170 470158 190226
rect 470214 190170 470282 190226
rect 470338 190170 470406 190226
rect 470462 190170 495878 190226
rect 495934 190170 496002 190226
rect 496058 190170 500754 190226
rect 500810 190170 500878 190226
rect 500934 190170 501002 190226
rect 501058 190170 501126 190226
rect 501182 190170 531474 190226
rect 531530 190170 531598 190226
rect 531654 190170 531722 190226
rect 531778 190170 531846 190226
rect 531902 190170 557878 190226
rect 557934 190170 558002 190226
rect 558058 190170 562194 190226
rect 562250 190170 562318 190226
rect 562374 190170 562442 190226
rect 562498 190170 562566 190226
rect 562622 190170 592914 190226
rect 592970 190170 593038 190226
rect 593094 190170 593162 190226
rect 593218 190170 593286 190226
rect 593342 190170 597456 190226
rect 597512 190170 597580 190226
rect 597636 190170 597704 190226
rect 597760 190170 597828 190226
rect 597884 190170 597980 190226
rect -1916 190102 597980 190170
rect -1916 190046 -1820 190102
rect -1764 190046 -1696 190102
rect -1640 190046 -1572 190102
rect -1516 190046 -1448 190102
rect -1392 190046 9234 190102
rect 9290 190046 9358 190102
rect 9414 190046 9482 190102
rect 9538 190046 9606 190102
rect 9662 190046 39878 190102
rect 39934 190046 40002 190102
rect 40058 190046 70674 190102
rect 70730 190046 70798 190102
rect 70854 190046 70922 190102
rect 70978 190046 71046 190102
rect 71102 190046 101878 190102
rect 101934 190046 102002 190102
rect 102058 190046 132114 190102
rect 132170 190046 132238 190102
rect 132294 190046 132362 190102
rect 132418 190046 132486 190102
rect 132542 190046 163878 190102
rect 163934 190046 164002 190102
rect 164058 190046 193554 190102
rect 193610 190046 193678 190102
rect 193734 190046 193802 190102
rect 193858 190046 193926 190102
rect 193982 190046 224274 190102
rect 224330 190046 224398 190102
rect 224454 190046 224522 190102
rect 224578 190046 224646 190102
rect 224702 190046 225878 190102
rect 225934 190046 226002 190102
rect 226058 190046 254994 190102
rect 255050 190046 255118 190102
rect 255174 190046 255242 190102
rect 255298 190046 255366 190102
rect 255422 190046 287878 190102
rect 287934 190046 288002 190102
rect 288058 190046 318598 190102
rect 318654 190046 318722 190102
rect 318778 190046 347154 190102
rect 347210 190046 347278 190102
rect 347334 190046 347402 190102
rect 347458 190046 347526 190102
rect 347582 190046 371878 190102
rect 371934 190046 372002 190102
rect 372058 190046 377874 190102
rect 377930 190046 377998 190102
rect 378054 190046 378122 190102
rect 378178 190046 378246 190102
rect 378302 190046 408594 190102
rect 408650 190046 408718 190102
rect 408774 190046 408842 190102
rect 408898 190046 408966 190102
rect 409022 190046 433878 190102
rect 433934 190046 434002 190102
rect 434058 190046 439314 190102
rect 439370 190046 439438 190102
rect 439494 190046 439562 190102
rect 439618 190046 439686 190102
rect 439742 190046 470034 190102
rect 470090 190046 470158 190102
rect 470214 190046 470282 190102
rect 470338 190046 470406 190102
rect 470462 190046 495878 190102
rect 495934 190046 496002 190102
rect 496058 190046 500754 190102
rect 500810 190046 500878 190102
rect 500934 190046 501002 190102
rect 501058 190046 501126 190102
rect 501182 190046 531474 190102
rect 531530 190046 531598 190102
rect 531654 190046 531722 190102
rect 531778 190046 531846 190102
rect 531902 190046 557878 190102
rect 557934 190046 558002 190102
rect 558058 190046 562194 190102
rect 562250 190046 562318 190102
rect 562374 190046 562442 190102
rect 562498 190046 562566 190102
rect 562622 190046 592914 190102
rect 592970 190046 593038 190102
rect 593094 190046 593162 190102
rect 593218 190046 593286 190102
rect 593342 190046 597456 190102
rect 597512 190046 597580 190102
rect 597636 190046 597704 190102
rect 597760 190046 597828 190102
rect 597884 190046 597980 190102
rect -1916 189978 597980 190046
rect -1916 189922 -1820 189978
rect -1764 189922 -1696 189978
rect -1640 189922 -1572 189978
rect -1516 189922 -1448 189978
rect -1392 189922 9234 189978
rect 9290 189922 9358 189978
rect 9414 189922 9482 189978
rect 9538 189922 9606 189978
rect 9662 189922 39878 189978
rect 39934 189922 40002 189978
rect 40058 189922 70674 189978
rect 70730 189922 70798 189978
rect 70854 189922 70922 189978
rect 70978 189922 71046 189978
rect 71102 189922 101878 189978
rect 101934 189922 102002 189978
rect 102058 189922 132114 189978
rect 132170 189922 132238 189978
rect 132294 189922 132362 189978
rect 132418 189922 132486 189978
rect 132542 189922 163878 189978
rect 163934 189922 164002 189978
rect 164058 189922 193554 189978
rect 193610 189922 193678 189978
rect 193734 189922 193802 189978
rect 193858 189922 193926 189978
rect 193982 189922 224274 189978
rect 224330 189922 224398 189978
rect 224454 189922 224522 189978
rect 224578 189922 224646 189978
rect 224702 189922 225878 189978
rect 225934 189922 226002 189978
rect 226058 189922 254994 189978
rect 255050 189922 255118 189978
rect 255174 189922 255242 189978
rect 255298 189922 255366 189978
rect 255422 189922 287878 189978
rect 287934 189922 288002 189978
rect 288058 189922 318598 189978
rect 318654 189922 318722 189978
rect 318778 189922 347154 189978
rect 347210 189922 347278 189978
rect 347334 189922 347402 189978
rect 347458 189922 347526 189978
rect 347582 189922 371878 189978
rect 371934 189922 372002 189978
rect 372058 189922 377874 189978
rect 377930 189922 377998 189978
rect 378054 189922 378122 189978
rect 378178 189922 378246 189978
rect 378302 189922 408594 189978
rect 408650 189922 408718 189978
rect 408774 189922 408842 189978
rect 408898 189922 408966 189978
rect 409022 189922 433878 189978
rect 433934 189922 434002 189978
rect 434058 189922 439314 189978
rect 439370 189922 439438 189978
rect 439494 189922 439562 189978
rect 439618 189922 439686 189978
rect 439742 189922 470034 189978
rect 470090 189922 470158 189978
rect 470214 189922 470282 189978
rect 470338 189922 470406 189978
rect 470462 189922 495878 189978
rect 495934 189922 496002 189978
rect 496058 189922 500754 189978
rect 500810 189922 500878 189978
rect 500934 189922 501002 189978
rect 501058 189922 501126 189978
rect 501182 189922 531474 189978
rect 531530 189922 531598 189978
rect 531654 189922 531722 189978
rect 531778 189922 531846 189978
rect 531902 189922 557878 189978
rect 557934 189922 558002 189978
rect 558058 189922 562194 189978
rect 562250 189922 562318 189978
rect 562374 189922 562442 189978
rect 562498 189922 562566 189978
rect 562622 189922 592914 189978
rect 592970 189922 593038 189978
rect 593094 189922 593162 189978
rect 593218 189922 593286 189978
rect 593342 189922 597456 189978
rect 597512 189922 597580 189978
rect 597636 189922 597704 189978
rect 597760 189922 597828 189978
rect 597884 189922 597980 189978
rect -1916 189826 597980 189922
rect 169692 189658 263860 189674
rect 169692 189602 169708 189658
rect 169764 189602 263788 189658
rect 263844 189602 263860 189658
rect 169692 189586 263860 189602
rect 403212 189658 472180 189674
rect 403212 189602 403228 189658
rect 403284 189602 472108 189658
rect 472164 189602 472180 189658
rect 403212 189586 472180 189602
rect 188060 189478 263972 189494
rect 188060 189422 188076 189478
rect 188132 189422 263900 189478
rect 263956 189422 263972 189478
rect 188060 189406 263972 189422
rect 335116 188938 394900 188954
rect 335116 188882 335132 188938
rect 335188 188882 394828 188938
rect 394884 188882 394900 188938
rect 335116 188866 394900 188882
rect 341836 188038 472180 188054
rect 341836 187982 341852 188038
rect 341908 187982 472108 188038
rect 472164 187982 472180 188038
rect 341836 187966 472180 187982
rect 187276 187498 263972 187514
rect 187276 187442 187292 187498
rect 187348 187442 263900 187498
rect 263956 187442 263972 187498
rect 187276 187426 263972 187442
rect 169692 187318 264084 187334
rect 169692 187262 169708 187318
rect 169764 187262 264012 187318
rect 264068 187262 264084 187318
rect 169692 187246 264084 187262
rect 336124 187318 396580 187334
rect 336124 187262 336140 187318
rect 336196 187262 396508 187318
rect 396564 187262 396580 187318
rect 336124 187246 396580 187262
rect 20060 186418 258708 186434
rect 20060 186362 20076 186418
rect 20132 186362 258636 186418
rect 258692 186362 258708 186418
rect 20060 186346 258708 186362
rect 336012 186418 455380 186434
rect 336012 186362 336028 186418
rect 336084 186362 455308 186418
rect 455364 186362 455380 186418
rect 336012 186346 455380 186362
rect 127580 186238 258484 186254
rect 127580 186182 127596 186238
rect 127652 186182 258412 186238
rect 258468 186182 258484 186238
rect 127580 186166 258484 186182
rect 342620 186238 393332 186254
rect 342620 186182 342636 186238
rect 342692 186182 393260 186238
rect 393316 186182 393332 186238
rect 342620 186166 393332 186182
rect 82668 186058 169780 186074
rect 82668 186002 82684 186058
rect 82740 186002 169708 186058
rect 169764 186002 169780 186058
rect 82668 185986 169780 186002
rect 191532 186058 263860 186074
rect 191532 186002 191548 186058
rect 191604 186002 263788 186058
rect 263844 186002 263860 186058
rect 191532 185986 263860 186002
rect -1916 184350 597980 184446
rect -1916 184294 -860 184350
rect -804 184294 -736 184350
rect -680 184294 -612 184350
rect -556 184294 -488 184350
rect -432 184294 5514 184350
rect 5570 184294 5638 184350
rect 5694 184294 5762 184350
rect 5818 184294 5886 184350
rect 5942 184294 24518 184350
rect 24574 184294 24642 184350
rect 24698 184294 36234 184350
rect 36290 184294 36358 184350
rect 36414 184294 36482 184350
rect 36538 184294 36606 184350
rect 36662 184294 55238 184350
rect 55294 184294 55362 184350
rect 55418 184294 66954 184350
rect 67010 184294 67078 184350
rect 67134 184294 67202 184350
rect 67258 184294 67326 184350
rect 67382 184294 86518 184350
rect 86574 184294 86642 184350
rect 86698 184294 97674 184350
rect 97730 184294 97798 184350
rect 97854 184294 97922 184350
rect 97978 184294 98046 184350
rect 98102 184294 117238 184350
rect 117294 184294 117362 184350
rect 117418 184294 128394 184350
rect 128450 184294 128518 184350
rect 128574 184294 128642 184350
rect 128698 184294 128766 184350
rect 128822 184294 148518 184350
rect 148574 184294 148642 184350
rect 148698 184294 159114 184350
rect 159170 184294 159238 184350
rect 159294 184294 159362 184350
rect 159418 184294 159486 184350
rect 159542 184294 179238 184350
rect 179294 184294 179362 184350
rect 179418 184294 189834 184350
rect 189890 184294 189958 184350
rect 190014 184294 190082 184350
rect 190138 184294 190206 184350
rect 190262 184294 210518 184350
rect 210574 184294 210642 184350
rect 210698 184294 220554 184350
rect 220610 184294 220678 184350
rect 220734 184294 220802 184350
rect 220858 184294 220926 184350
rect 220982 184294 241238 184350
rect 241294 184294 241362 184350
rect 241418 184294 251274 184350
rect 251330 184294 251398 184350
rect 251454 184294 251522 184350
rect 251578 184294 251646 184350
rect 251702 184294 272518 184350
rect 272574 184294 272642 184350
rect 272698 184294 303238 184350
rect 303294 184294 303362 184350
rect 303418 184294 343434 184350
rect 343490 184294 343558 184350
rect 343614 184294 343682 184350
rect 343738 184294 343806 184350
rect 343862 184294 356518 184350
rect 356574 184294 356642 184350
rect 356698 184294 374154 184350
rect 374210 184294 374278 184350
rect 374334 184294 374402 184350
rect 374458 184294 374526 184350
rect 374582 184294 387238 184350
rect 387294 184294 387362 184350
rect 387418 184294 404874 184350
rect 404930 184294 404998 184350
rect 405054 184294 405122 184350
rect 405178 184294 405246 184350
rect 405302 184294 418518 184350
rect 418574 184294 418642 184350
rect 418698 184294 435594 184350
rect 435650 184294 435718 184350
rect 435774 184294 435842 184350
rect 435898 184294 435966 184350
rect 436022 184294 449238 184350
rect 449294 184294 449362 184350
rect 449418 184294 466314 184350
rect 466370 184294 466438 184350
rect 466494 184294 466562 184350
rect 466618 184294 466686 184350
rect 466742 184294 480518 184350
rect 480574 184294 480642 184350
rect 480698 184294 497034 184350
rect 497090 184294 497158 184350
rect 497214 184294 497282 184350
rect 497338 184294 497406 184350
rect 497462 184294 511238 184350
rect 511294 184294 511362 184350
rect 511418 184294 527754 184350
rect 527810 184294 527878 184350
rect 527934 184294 528002 184350
rect 528058 184294 528126 184350
rect 528182 184294 542518 184350
rect 542574 184294 542642 184350
rect 542698 184294 558474 184350
rect 558530 184294 558598 184350
rect 558654 184294 558722 184350
rect 558778 184294 558846 184350
rect 558902 184294 573238 184350
rect 573294 184294 573362 184350
rect 573418 184294 589194 184350
rect 589250 184294 589318 184350
rect 589374 184294 589442 184350
rect 589498 184294 589566 184350
rect 589622 184294 596496 184350
rect 596552 184294 596620 184350
rect 596676 184294 596744 184350
rect 596800 184294 596868 184350
rect 596924 184294 597980 184350
rect -1916 184226 597980 184294
rect -1916 184170 -860 184226
rect -804 184170 -736 184226
rect -680 184170 -612 184226
rect -556 184170 -488 184226
rect -432 184170 5514 184226
rect 5570 184170 5638 184226
rect 5694 184170 5762 184226
rect 5818 184170 5886 184226
rect 5942 184170 24518 184226
rect 24574 184170 24642 184226
rect 24698 184170 36234 184226
rect 36290 184170 36358 184226
rect 36414 184170 36482 184226
rect 36538 184170 36606 184226
rect 36662 184170 55238 184226
rect 55294 184170 55362 184226
rect 55418 184170 66954 184226
rect 67010 184170 67078 184226
rect 67134 184170 67202 184226
rect 67258 184170 67326 184226
rect 67382 184170 86518 184226
rect 86574 184170 86642 184226
rect 86698 184170 97674 184226
rect 97730 184170 97798 184226
rect 97854 184170 97922 184226
rect 97978 184170 98046 184226
rect 98102 184170 117238 184226
rect 117294 184170 117362 184226
rect 117418 184170 128394 184226
rect 128450 184170 128518 184226
rect 128574 184170 128642 184226
rect 128698 184170 128766 184226
rect 128822 184170 148518 184226
rect 148574 184170 148642 184226
rect 148698 184170 159114 184226
rect 159170 184170 159238 184226
rect 159294 184170 159362 184226
rect 159418 184170 159486 184226
rect 159542 184170 179238 184226
rect 179294 184170 179362 184226
rect 179418 184170 189834 184226
rect 189890 184170 189958 184226
rect 190014 184170 190082 184226
rect 190138 184170 190206 184226
rect 190262 184170 210518 184226
rect 210574 184170 210642 184226
rect 210698 184170 220554 184226
rect 220610 184170 220678 184226
rect 220734 184170 220802 184226
rect 220858 184170 220926 184226
rect 220982 184170 241238 184226
rect 241294 184170 241362 184226
rect 241418 184170 251274 184226
rect 251330 184170 251398 184226
rect 251454 184170 251522 184226
rect 251578 184170 251646 184226
rect 251702 184170 272518 184226
rect 272574 184170 272642 184226
rect 272698 184170 303238 184226
rect 303294 184170 303362 184226
rect 303418 184170 343434 184226
rect 343490 184170 343558 184226
rect 343614 184170 343682 184226
rect 343738 184170 343806 184226
rect 343862 184170 356518 184226
rect 356574 184170 356642 184226
rect 356698 184170 374154 184226
rect 374210 184170 374278 184226
rect 374334 184170 374402 184226
rect 374458 184170 374526 184226
rect 374582 184170 387238 184226
rect 387294 184170 387362 184226
rect 387418 184170 404874 184226
rect 404930 184170 404998 184226
rect 405054 184170 405122 184226
rect 405178 184170 405246 184226
rect 405302 184170 418518 184226
rect 418574 184170 418642 184226
rect 418698 184170 435594 184226
rect 435650 184170 435718 184226
rect 435774 184170 435842 184226
rect 435898 184170 435966 184226
rect 436022 184170 449238 184226
rect 449294 184170 449362 184226
rect 449418 184170 466314 184226
rect 466370 184170 466438 184226
rect 466494 184170 466562 184226
rect 466618 184170 466686 184226
rect 466742 184170 480518 184226
rect 480574 184170 480642 184226
rect 480698 184170 497034 184226
rect 497090 184170 497158 184226
rect 497214 184170 497282 184226
rect 497338 184170 497406 184226
rect 497462 184170 511238 184226
rect 511294 184170 511362 184226
rect 511418 184170 527754 184226
rect 527810 184170 527878 184226
rect 527934 184170 528002 184226
rect 528058 184170 528126 184226
rect 528182 184170 542518 184226
rect 542574 184170 542642 184226
rect 542698 184170 558474 184226
rect 558530 184170 558598 184226
rect 558654 184170 558722 184226
rect 558778 184170 558846 184226
rect 558902 184170 573238 184226
rect 573294 184170 573362 184226
rect 573418 184170 589194 184226
rect 589250 184170 589318 184226
rect 589374 184170 589442 184226
rect 589498 184170 589566 184226
rect 589622 184170 596496 184226
rect 596552 184170 596620 184226
rect 596676 184170 596744 184226
rect 596800 184170 596868 184226
rect 596924 184170 597980 184226
rect -1916 184102 597980 184170
rect -1916 184046 -860 184102
rect -804 184046 -736 184102
rect -680 184046 -612 184102
rect -556 184046 -488 184102
rect -432 184046 5514 184102
rect 5570 184046 5638 184102
rect 5694 184046 5762 184102
rect 5818 184046 5886 184102
rect 5942 184046 24518 184102
rect 24574 184046 24642 184102
rect 24698 184046 36234 184102
rect 36290 184046 36358 184102
rect 36414 184046 36482 184102
rect 36538 184046 36606 184102
rect 36662 184046 55238 184102
rect 55294 184046 55362 184102
rect 55418 184046 66954 184102
rect 67010 184046 67078 184102
rect 67134 184046 67202 184102
rect 67258 184046 67326 184102
rect 67382 184046 86518 184102
rect 86574 184046 86642 184102
rect 86698 184046 97674 184102
rect 97730 184046 97798 184102
rect 97854 184046 97922 184102
rect 97978 184046 98046 184102
rect 98102 184046 117238 184102
rect 117294 184046 117362 184102
rect 117418 184046 128394 184102
rect 128450 184046 128518 184102
rect 128574 184046 128642 184102
rect 128698 184046 128766 184102
rect 128822 184046 148518 184102
rect 148574 184046 148642 184102
rect 148698 184046 159114 184102
rect 159170 184046 159238 184102
rect 159294 184046 159362 184102
rect 159418 184046 159486 184102
rect 159542 184046 179238 184102
rect 179294 184046 179362 184102
rect 179418 184046 189834 184102
rect 189890 184046 189958 184102
rect 190014 184046 190082 184102
rect 190138 184046 190206 184102
rect 190262 184046 210518 184102
rect 210574 184046 210642 184102
rect 210698 184046 220554 184102
rect 220610 184046 220678 184102
rect 220734 184046 220802 184102
rect 220858 184046 220926 184102
rect 220982 184046 241238 184102
rect 241294 184046 241362 184102
rect 241418 184046 251274 184102
rect 251330 184046 251398 184102
rect 251454 184046 251522 184102
rect 251578 184046 251646 184102
rect 251702 184046 272518 184102
rect 272574 184046 272642 184102
rect 272698 184046 303238 184102
rect 303294 184046 303362 184102
rect 303418 184046 343434 184102
rect 343490 184046 343558 184102
rect 343614 184046 343682 184102
rect 343738 184046 343806 184102
rect 343862 184046 356518 184102
rect 356574 184046 356642 184102
rect 356698 184046 374154 184102
rect 374210 184046 374278 184102
rect 374334 184046 374402 184102
rect 374458 184046 374526 184102
rect 374582 184046 387238 184102
rect 387294 184046 387362 184102
rect 387418 184046 404874 184102
rect 404930 184046 404998 184102
rect 405054 184046 405122 184102
rect 405178 184046 405246 184102
rect 405302 184046 418518 184102
rect 418574 184046 418642 184102
rect 418698 184046 435594 184102
rect 435650 184046 435718 184102
rect 435774 184046 435842 184102
rect 435898 184046 435966 184102
rect 436022 184046 449238 184102
rect 449294 184046 449362 184102
rect 449418 184046 466314 184102
rect 466370 184046 466438 184102
rect 466494 184046 466562 184102
rect 466618 184046 466686 184102
rect 466742 184046 480518 184102
rect 480574 184046 480642 184102
rect 480698 184046 497034 184102
rect 497090 184046 497158 184102
rect 497214 184046 497282 184102
rect 497338 184046 497406 184102
rect 497462 184046 511238 184102
rect 511294 184046 511362 184102
rect 511418 184046 527754 184102
rect 527810 184046 527878 184102
rect 527934 184046 528002 184102
rect 528058 184046 528126 184102
rect 528182 184046 542518 184102
rect 542574 184046 542642 184102
rect 542698 184046 558474 184102
rect 558530 184046 558598 184102
rect 558654 184046 558722 184102
rect 558778 184046 558846 184102
rect 558902 184046 573238 184102
rect 573294 184046 573362 184102
rect 573418 184046 589194 184102
rect 589250 184046 589318 184102
rect 589374 184046 589442 184102
rect 589498 184046 589566 184102
rect 589622 184046 596496 184102
rect 596552 184046 596620 184102
rect 596676 184046 596744 184102
rect 596800 184046 596868 184102
rect 596924 184046 597980 184102
rect -1916 183978 597980 184046
rect -1916 183922 -860 183978
rect -804 183922 -736 183978
rect -680 183922 -612 183978
rect -556 183922 -488 183978
rect -432 183922 5514 183978
rect 5570 183922 5638 183978
rect 5694 183922 5762 183978
rect 5818 183922 5886 183978
rect 5942 183922 24518 183978
rect 24574 183922 24642 183978
rect 24698 183922 36234 183978
rect 36290 183922 36358 183978
rect 36414 183922 36482 183978
rect 36538 183922 36606 183978
rect 36662 183922 55238 183978
rect 55294 183922 55362 183978
rect 55418 183922 66954 183978
rect 67010 183922 67078 183978
rect 67134 183922 67202 183978
rect 67258 183922 67326 183978
rect 67382 183922 86518 183978
rect 86574 183922 86642 183978
rect 86698 183922 97674 183978
rect 97730 183922 97798 183978
rect 97854 183922 97922 183978
rect 97978 183922 98046 183978
rect 98102 183922 117238 183978
rect 117294 183922 117362 183978
rect 117418 183922 128394 183978
rect 128450 183922 128518 183978
rect 128574 183922 128642 183978
rect 128698 183922 128766 183978
rect 128822 183922 148518 183978
rect 148574 183922 148642 183978
rect 148698 183922 159114 183978
rect 159170 183922 159238 183978
rect 159294 183922 159362 183978
rect 159418 183922 159486 183978
rect 159542 183922 179238 183978
rect 179294 183922 179362 183978
rect 179418 183922 189834 183978
rect 189890 183922 189958 183978
rect 190014 183922 190082 183978
rect 190138 183922 190206 183978
rect 190262 183922 210518 183978
rect 210574 183922 210642 183978
rect 210698 183922 220554 183978
rect 220610 183922 220678 183978
rect 220734 183922 220802 183978
rect 220858 183922 220926 183978
rect 220982 183922 241238 183978
rect 241294 183922 241362 183978
rect 241418 183922 251274 183978
rect 251330 183922 251398 183978
rect 251454 183922 251522 183978
rect 251578 183922 251646 183978
rect 251702 183922 272518 183978
rect 272574 183922 272642 183978
rect 272698 183922 303238 183978
rect 303294 183922 303362 183978
rect 303418 183922 343434 183978
rect 343490 183922 343558 183978
rect 343614 183922 343682 183978
rect 343738 183922 343806 183978
rect 343862 183922 356518 183978
rect 356574 183922 356642 183978
rect 356698 183922 374154 183978
rect 374210 183922 374278 183978
rect 374334 183922 374402 183978
rect 374458 183922 374526 183978
rect 374582 183922 387238 183978
rect 387294 183922 387362 183978
rect 387418 183922 404874 183978
rect 404930 183922 404998 183978
rect 405054 183922 405122 183978
rect 405178 183922 405246 183978
rect 405302 183922 418518 183978
rect 418574 183922 418642 183978
rect 418698 183922 435594 183978
rect 435650 183922 435718 183978
rect 435774 183922 435842 183978
rect 435898 183922 435966 183978
rect 436022 183922 449238 183978
rect 449294 183922 449362 183978
rect 449418 183922 466314 183978
rect 466370 183922 466438 183978
rect 466494 183922 466562 183978
rect 466618 183922 466686 183978
rect 466742 183922 480518 183978
rect 480574 183922 480642 183978
rect 480698 183922 497034 183978
rect 497090 183922 497158 183978
rect 497214 183922 497282 183978
rect 497338 183922 497406 183978
rect 497462 183922 511238 183978
rect 511294 183922 511362 183978
rect 511418 183922 527754 183978
rect 527810 183922 527878 183978
rect 527934 183922 528002 183978
rect 528058 183922 528126 183978
rect 528182 183922 542518 183978
rect 542574 183922 542642 183978
rect 542698 183922 558474 183978
rect 558530 183922 558598 183978
rect 558654 183922 558722 183978
rect 558778 183922 558846 183978
rect 558902 183922 573238 183978
rect 573294 183922 573362 183978
rect 573418 183922 589194 183978
rect 589250 183922 589318 183978
rect 589374 183922 589442 183978
rect 589498 183922 589566 183978
rect 589622 183922 596496 183978
rect 596552 183922 596620 183978
rect 596676 183922 596744 183978
rect 596800 183922 596868 183978
rect 596924 183922 597980 183978
rect -1916 183826 597980 183922
rect -1916 172350 597980 172446
rect -1916 172294 -1820 172350
rect -1764 172294 -1696 172350
rect -1640 172294 -1572 172350
rect -1516 172294 -1448 172350
rect -1392 172294 9234 172350
rect 9290 172294 9358 172350
rect 9414 172294 9482 172350
rect 9538 172294 9606 172350
rect 9662 172294 39954 172350
rect 40010 172294 40078 172350
rect 40134 172294 40202 172350
rect 40258 172294 40326 172350
rect 40382 172294 70674 172350
rect 70730 172294 70798 172350
rect 70854 172294 70922 172350
rect 70978 172294 71046 172350
rect 71102 172294 101394 172350
rect 101450 172294 101518 172350
rect 101574 172294 101642 172350
rect 101698 172294 101766 172350
rect 101822 172294 132114 172350
rect 132170 172294 132238 172350
rect 132294 172294 132362 172350
rect 132418 172294 132486 172350
rect 132542 172294 162834 172350
rect 162890 172294 162958 172350
rect 163014 172294 163082 172350
rect 163138 172294 163206 172350
rect 163262 172294 193554 172350
rect 193610 172294 193678 172350
rect 193734 172294 193802 172350
rect 193858 172294 193926 172350
rect 193982 172294 224274 172350
rect 224330 172294 224398 172350
rect 224454 172294 224522 172350
rect 224578 172294 224646 172350
rect 224702 172294 254994 172350
rect 255050 172294 255118 172350
rect 255174 172294 255242 172350
rect 255298 172294 255366 172350
rect 255422 172294 287878 172350
rect 287934 172294 288002 172350
rect 288058 172294 318598 172350
rect 318654 172294 318722 172350
rect 318778 172294 347154 172350
rect 347210 172294 347278 172350
rect 347334 172294 347402 172350
rect 347458 172294 347526 172350
rect 347582 172294 377874 172350
rect 377930 172294 377998 172350
rect 378054 172294 378122 172350
rect 378178 172294 378246 172350
rect 378302 172294 408594 172350
rect 408650 172294 408718 172350
rect 408774 172294 408842 172350
rect 408898 172294 408966 172350
rect 409022 172294 439314 172350
rect 439370 172294 439438 172350
rect 439494 172294 439562 172350
rect 439618 172294 439686 172350
rect 439742 172294 470034 172350
rect 470090 172294 470158 172350
rect 470214 172294 470282 172350
rect 470338 172294 470406 172350
rect 470462 172294 500754 172350
rect 500810 172294 500878 172350
rect 500934 172294 501002 172350
rect 501058 172294 501126 172350
rect 501182 172294 531474 172350
rect 531530 172294 531598 172350
rect 531654 172294 531722 172350
rect 531778 172294 531846 172350
rect 531902 172294 562194 172350
rect 562250 172294 562318 172350
rect 562374 172294 562442 172350
rect 562498 172294 562566 172350
rect 562622 172294 592914 172350
rect 592970 172294 593038 172350
rect 593094 172294 593162 172350
rect 593218 172294 593286 172350
rect 593342 172294 597456 172350
rect 597512 172294 597580 172350
rect 597636 172294 597704 172350
rect 597760 172294 597828 172350
rect 597884 172294 597980 172350
rect -1916 172226 597980 172294
rect -1916 172170 -1820 172226
rect -1764 172170 -1696 172226
rect -1640 172170 -1572 172226
rect -1516 172170 -1448 172226
rect -1392 172170 9234 172226
rect 9290 172170 9358 172226
rect 9414 172170 9482 172226
rect 9538 172170 9606 172226
rect 9662 172170 39954 172226
rect 40010 172170 40078 172226
rect 40134 172170 40202 172226
rect 40258 172170 40326 172226
rect 40382 172170 70674 172226
rect 70730 172170 70798 172226
rect 70854 172170 70922 172226
rect 70978 172170 71046 172226
rect 71102 172170 101394 172226
rect 101450 172170 101518 172226
rect 101574 172170 101642 172226
rect 101698 172170 101766 172226
rect 101822 172170 132114 172226
rect 132170 172170 132238 172226
rect 132294 172170 132362 172226
rect 132418 172170 132486 172226
rect 132542 172170 162834 172226
rect 162890 172170 162958 172226
rect 163014 172170 163082 172226
rect 163138 172170 163206 172226
rect 163262 172170 193554 172226
rect 193610 172170 193678 172226
rect 193734 172170 193802 172226
rect 193858 172170 193926 172226
rect 193982 172170 224274 172226
rect 224330 172170 224398 172226
rect 224454 172170 224522 172226
rect 224578 172170 224646 172226
rect 224702 172170 254994 172226
rect 255050 172170 255118 172226
rect 255174 172170 255242 172226
rect 255298 172170 255366 172226
rect 255422 172170 287878 172226
rect 287934 172170 288002 172226
rect 288058 172170 318598 172226
rect 318654 172170 318722 172226
rect 318778 172170 347154 172226
rect 347210 172170 347278 172226
rect 347334 172170 347402 172226
rect 347458 172170 347526 172226
rect 347582 172170 377874 172226
rect 377930 172170 377998 172226
rect 378054 172170 378122 172226
rect 378178 172170 378246 172226
rect 378302 172170 408594 172226
rect 408650 172170 408718 172226
rect 408774 172170 408842 172226
rect 408898 172170 408966 172226
rect 409022 172170 439314 172226
rect 439370 172170 439438 172226
rect 439494 172170 439562 172226
rect 439618 172170 439686 172226
rect 439742 172170 470034 172226
rect 470090 172170 470158 172226
rect 470214 172170 470282 172226
rect 470338 172170 470406 172226
rect 470462 172170 500754 172226
rect 500810 172170 500878 172226
rect 500934 172170 501002 172226
rect 501058 172170 501126 172226
rect 501182 172170 531474 172226
rect 531530 172170 531598 172226
rect 531654 172170 531722 172226
rect 531778 172170 531846 172226
rect 531902 172170 562194 172226
rect 562250 172170 562318 172226
rect 562374 172170 562442 172226
rect 562498 172170 562566 172226
rect 562622 172170 592914 172226
rect 592970 172170 593038 172226
rect 593094 172170 593162 172226
rect 593218 172170 593286 172226
rect 593342 172170 597456 172226
rect 597512 172170 597580 172226
rect 597636 172170 597704 172226
rect 597760 172170 597828 172226
rect 597884 172170 597980 172226
rect -1916 172102 597980 172170
rect -1916 172046 -1820 172102
rect -1764 172046 -1696 172102
rect -1640 172046 -1572 172102
rect -1516 172046 -1448 172102
rect -1392 172046 9234 172102
rect 9290 172046 9358 172102
rect 9414 172046 9482 172102
rect 9538 172046 9606 172102
rect 9662 172046 39954 172102
rect 40010 172046 40078 172102
rect 40134 172046 40202 172102
rect 40258 172046 40326 172102
rect 40382 172046 70674 172102
rect 70730 172046 70798 172102
rect 70854 172046 70922 172102
rect 70978 172046 71046 172102
rect 71102 172046 101394 172102
rect 101450 172046 101518 172102
rect 101574 172046 101642 172102
rect 101698 172046 101766 172102
rect 101822 172046 132114 172102
rect 132170 172046 132238 172102
rect 132294 172046 132362 172102
rect 132418 172046 132486 172102
rect 132542 172046 162834 172102
rect 162890 172046 162958 172102
rect 163014 172046 163082 172102
rect 163138 172046 163206 172102
rect 163262 172046 193554 172102
rect 193610 172046 193678 172102
rect 193734 172046 193802 172102
rect 193858 172046 193926 172102
rect 193982 172046 224274 172102
rect 224330 172046 224398 172102
rect 224454 172046 224522 172102
rect 224578 172046 224646 172102
rect 224702 172046 254994 172102
rect 255050 172046 255118 172102
rect 255174 172046 255242 172102
rect 255298 172046 255366 172102
rect 255422 172046 287878 172102
rect 287934 172046 288002 172102
rect 288058 172046 318598 172102
rect 318654 172046 318722 172102
rect 318778 172046 347154 172102
rect 347210 172046 347278 172102
rect 347334 172046 347402 172102
rect 347458 172046 347526 172102
rect 347582 172046 377874 172102
rect 377930 172046 377998 172102
rect 378054 172046 378122 172102
rect 378178 172046 378246 172102
rect 378302 172046 408594 172102
rect 408650 172046 408718 172102
rect 408774 172046 408842 172102
rect 408898 172046 408966 172102
rect 409022 172046 439314 172102
rect 439370 172046 439438 172102
rect 439494 172046 439562 172102
rect 439618 172046 439686 172102
rect 439742 172046 470034 172102
rect 470090 172046 470158 172102
rect 470214 172046 470282 172102
rect 470338 172046 470406 172102
rect 470462 172046 500754 172102
rect 500810 172046 500878 172102
rect 500934 172046 501002 172102
rect 501058 172046 501126 172102
rect 501182 172046 531474 172102
rect 531530 172046 531598 172102
rect 531654 172046 531722 172102
rect 531778 172046 531846 172102
rect 531902 172046 562194 172102
rect 562250 172046 562318 172102
rect 562374 172046 562442 172102
rect 562498 172046 562566 172102
rect 562622 172046 592914 172102
rect 592970 172046 593038 172102
rect 593094 172046 593162 172102
rect 593218 172046 593286 172102
rect 593342 172046 597456 172102
rect 597512 172046 597580 172102
rect 597636 172046 597704 172102
rect 597760 172046 597828 172102
rect 597884 172046 597980 172102
rect -1916 171978 597980 172046
rect -1916 171922 -1820 171978
rect -1764 171922 -1696 171978
rect -1640 171922 -1572 171978
rect -1516 171922 -1448 171978
rect -1392 171922 9234 171978
rect 9290 171922 9358 171978
rect 9414 171922 9482 171978
rect 9538 171922 9606 171978
rect 9662 171922 39954 171978
rect 40010 171922 40078 171978
rect 40134 171922 40202 171978
rect 40258 171922 40326 171978
rect 40382 171922 70674 171978
rect 70730 171922 70798 171978
rect 70854 171922 70922 171978
rect 70978 171922 71046 171978
rect 71102 171922 101394 171978
rect 101450 171922 101518 171978
rect 101574 171922 101642 171978
rect 101698 171922 101766 171978
rect 101822 171922 132114 171978
rect 132170 171922 132238 171978
rect 132294 171922 132362 171978
rect 132418 171922 132486 171978
rect 132542 171922 162834 171978
rect 162890 171922 162958 171978
rect 163014 171922 163082 171978
rect 163138 171922 163206 171978
rect 163262 171922 193554 171978
rect 193610 171922 193678 171978
rect 193734 171922 193802 171978
rect 193858 171922 193926 171978
rect 193982 171922 224274 171978
rect 224330 171922 224398 171978
rect 224454 171922 224522 171978
rect 224578 171922 224646 171978
rect 224702 171922 254994 171978
rect 255050 171922 255118 171978
rect 255174 171922 255242 171978
rect 255298 171922 255366 171978
rect 255422 171922 287878 171978
rect 287934 171922 288002 171978
rect 288058 171922 318598 171978
rect 318654 171922 318722 171978
rect 318778 171922 347154 171978
rect 347210 171922 347278 171978
rect 347334 171922 347402 171978
rect 347458 171922 347526 171978
rect 347582 171922 377874 171978
rect 377930 171922 377998 171978
rect 378054 171922 378122 171978
rect 378178 171922 378246 171978
rect 378302 171922 408594 171978
rect 408650 171922 408718 171978
rect 408774 171922 408842 171978
rect 408898 171922 408966 171978
rect 409022 171922 439314 171978
rect 439370 171922 439438 171978
rect 439494 171922 439562 171978
rect 439618 171922 439686 171978
rect 439742 171922 470034 171978
rect 470090 171922 470158 171978
rect 470214 171922 470282 171978
rect 470338 171922 470406 171978
rect 470462 171922 500754 171978
rect 500810 171922 500878 171978
rect 500934 171922 501002 171978
rect 501058 171922 501126 171978
rect 501182 171922 531474 171978
rect 531530 171922 531598 171978
rect 531654 171922 531722 171978
rect 531778 171922 531846 171978
rect 531902 171922 562194 171978
rect 562250 171922 562318 171978
rect 562374 171922 562442 171978
rect 562498 171922 562566 171978
rect 562622 171922 592914 171978
rect 592970 171922 593038 171978
rect 593094 171922 593162 171978
rect 593218 171922 593286 171978
rect 593342 171922 597456 171978
rect 597512 171922 597580 171978
rect 597636 171922 597704 171978
rect 597760 171922 597828 171978
rect 597884 171922 597980 171978
rect -1916 171826 597980 171922
rect -1916 166350 597980 166446
rect -1916 166294 -860 166350
rect -804 166294 -736 166350
rect -680 166294 -612 166350
rect -556 166294 -488 166350
rect -432 166294 5514 166350
rect 5570 166294 5638 166350
rect 5694 166294 5762 166350
rect 5818 166294 5886 166350
rect 5942 166294 36234 166350
rect 36290 166294 36358 166350
rect 36414 166294 36482 166350
rect 36538 166294 36606 166350
rect 36662 166294 66954 166350
rect 67010 166294 67078 166350
rect 67134 166294 67202 166350
rect 67258 166294 67326 166350
rect 67382 166294 97674 166350
rect 97730 166294 97798 166350
rect 97854 166294 97922 166350
rect 97978 166294 98046 166350
rect 98102 166294 128394 166350
rect 128450 166294 128518 166350
rect 128574 166294 128642 166350
rect 128698 166294 128766 166350
rect 128822 166294 159114 166350
rect 159170 166294 159238 166350
rect 159294 166294 159362 166350
rect 159418 166294 159486 166350
rect 159542 166294 189834 166350
rect 189890 166294 189958 166350
rect 190014 166294 190082 166350
rect 190138 166294 190206 166350
rect 190262 166294 220554 166350
rect 220610 166294 220678 166350
rect 220734 166294 220802 166350
rect 220858 166294 220926 166350
rect 220982 166294 251274 166350
rect 251330 166294 251398 166350
rect 251454 166294 251522 166350
rect 251578 166294 251646 166350
rect 251702 166294 272518 166350
rect 272574 166294 272642 166350
rect 272698 166294 303238 166350
rect 303294 166294 303362 166350
rect 303418 166294 343434 166350
rect 343490 166294 343558 166350
rect 343614 166294 343682 166350
rect 343738 166294 343806 166350
rect 343862 166294 374154 166350
rect 374210 166294 374278 166350
rect 374334 166294 374402 166350
rect 374458 166294 374526 166350
rect 374582 166294 404874 166350
rect 404930 166294 404998 166350
rect 405054 166294 405122 166350
rect 405178 166294 405246 166350
rect 405302 166294 435594 166350
rect 435650 166294 435718 166350
rect 435774 166294 435842 166350
rect 435898 166294 435966 166350
rect 436022 166294 466314 166350
rect 466370 166294 466438 166350
rect 466494 166294 466562 166350
rect 466618 166294 466686 166350
rect 466742 166294 497034 166350
rect 497090 166294 497158 166350
rect 497214 166294 497282 166350
rect 497338 166294 497406 166350
rect 497462 166294 527754 166350
rect 527810 166294 527878 166350
rect 527934 166294 528002 166350
rect 528058 166294 528126 166350
rect 528182 166294 558474 166350
rect 558530 166294 558598 166350
rect 558654 166294 558722 166350
rect 558778 166294 558846 166350
rect 558902 166294 589194 166350
rect 589250 166294 589318 166350
rect 589374 166294 589442 166350
rect 589498 166294 589566 166350
rect 589622 166294 596496 166350
rect 596552 166294 596620 166350
rect 596676 166294 596744 166350
rect 596800 166294 596868 166350
rect 596924 166294 597980 166350
rect -1916 166226 597980 166294
rect -1916 166170 -860 166226
rect -804 166170 -736 166226
rect -680 166170 -612 166226
rect -556 166170 -488 166226
rect -432 166170 5514 166226
rect 5570 166170 5638 166226
rect 5694 166170 5762 166226
rect 5818 166170 5886 166226
rect 5942 166170 36234 166226
rect 36290 166170 36358 166226
rect 36414 166170 36482 166226
rect 36538 166170 36606 166226
rect 36662 166170 66954 166226
rect 67010 166170 67078 166226
rect 67134 166170 67202 166226
rect 67258 166170 67326 166226
rect 67382 166170 97674 166226
rect 97730 166170 97798 166226
rect 97854 166170 97922 166226
rect 97978 166170 98046 166226
rect 98102 166170 128394 166226
rect 128450 166170 128518 166226
rect 128574 166170 128642 166226
rect 128698 166170 128766 166226
rect 128822 166170 159114 166226
rect 159170 166170 159238 166226
rect 159294 166170 159362 166226
rect 159418 166170 159486 166226
rect 159542 166170 189834 166226
rect 189890 166170 189958 166226
rect 190014 166170 190082 166226
rect 190138 166170 190206 166226
rect 190262 166170 220554 166226
rect 220610 166170 220678 166226
rect 220734 166170 220802 166226
rect 220858 166170 220926 166226
rect 220982 166170 251274 166226
rect 251330 166170 251398 166226
rect 251454 166170 251522 166226
rect 251578 166170 251646 166226
rect 251702 166170 272518 166226
rect 272574 166170 272642 166226
rect 272698 166170 303238 166226
rect 303294 166170 303362 166226
rect 303418 166170 343434 166226
rect 343490 166170 343558 166226
rect 343614 166170 343682 166226
rect 343738 166170 343806 166226
rect 343862 166170 374154 166226
rect 374210 166170 374278 166226
rect 374334 166170 374402 166226
rect 374458 166170 374526 166226
rect 374582 166170 404874 166226
rect 404930 166170 404998 166226
rect 405054 166170 405122 166226
rect 405178 166170 405246 166226
rect 405302 166170 435594 166226
rect 435650 166170 435718 166226
rect 435774 166170 435842 166226
rect 435898 166170 435966 166226
rect 436022 166170 466314 166226
rect 466370 166170 466438 166226
rect 466494 166170 466562 166226
rect 466618 166170 466686 166226
rect 466742 166170 497034 166226
rect 497090 166170 497158 166226
rect 497214 166170 497282 166226
rect 497338 166170 497406 166226
rect 497462 166170 527754 166226
rect 527810 166170 527878 166226
rect 527934 166170 528002 166226
rect 528058 166170 528126 166226
rect 528182 166170 558474 166226
rect 558530 166170 558598 166226
rect 558654 166170 558722 166226
rect 558778 166170 558846 166226
rect 558902 166170 589194 166226
rect 589250 166170 589318 166226
rect 589374 166170 589442 166226
rect 589498 166170 589566 166226
rect 589622 166170 596496 166226
rect 596552 166170 596620 166226
rect 596676 166170 596744 166226
rect 596800 166170 596868 166226
rect 596924 166170 597980 166226
rect -1916 166102 597980 166170
rect -1916 166046 -860 166102
rect -804 166046 -736 166102
rect -680 166046 -612 166102
rect -556 166046 -488 166102
rect -432 166046 5514 166102
rect 5570 166046 5638 166102
rect 5694 166046 5762 166102
rect 5818 166046 5886 166102
rect 5942 166046 36234 166102
rect 36290 166046 36358 166102
rect 36414 166046 36482 166102
rect 36538 166046 36606 166102
rect 36662 166046 66954 166102
rect 67010 166046 67078 166102
rect 67134 166046 67202 166102
rect 67258 166046 67326 166102
rect 67382 166046 97674 166102
rect 97730 166046 97798 166102
rect 97854 166046 97922 166102
rect 97978 166046 98046 166102
rect 98102 166046 128394 166102
rect 128450 166046 128518 166102
rect 128574 166046 128642 166102
rect 128698 166046 128766 166102
rect 128822 166046 159114 166102
rect 159170 166046 159238 166102
rect 159294 166046 159362 166102
rect 159418 166046 159486 166102
rect 159542 166046 189834 166102
rect 189890 166046 189958 166102
rect 190014 166046 190082 166102
rect 190138 166046 190206 166102
rect 190262 166046 220554 166102
rect 220610 166046 220678 166102
rect 220734 166046 220802 166102
rect 220858 166046 220926 166102
rect 220982 166046 251274 166102
rect 251330 166046 251398 166102
rect 251454 166046 251522 166102
rect 251578 166046 251646 166102
rect 251702 166046 272518 166102
rect 272574 166046 272642 166102
rect 272698 166046 303238 166102
rect 303294 166046 303362 166102
rect 303418 166046 343434 166102
rect 343490 166046 343558 166102
rect 343614 166046 343682 166102
rect 343738 166046 343806 166102
rect 343862 166046 374154 166102
rect 374210 166046 374278 166102
rect 374334 166046 374402 166102
rect 374458 166046 374526 166102
rect 374582 166046 404874 166102
rect 404930 166046 404998 166102
rect 405054 166046 405122 166102
rect 405178 166046 405246 166102
rect 405302 166046 435594 166102
rect 435650 166046 435718 166102
rect 435774 166046 435842 166102
rect 435898 166046 435966 166102
rect 436022 166046 466314 166102
rect 466370 166046 466438 166102
rect 466494 166046 466562 166102
rect 466618 166046 466686 166102
rect 466742 166046 497034 166102
rect 497090 166046 497158 166102
rect 497214 166046 497282 166102
rect 497338 166046 497406 166102
rect 497462 166046 527754 166102
rect 527810 166046 527878 166102
rect 527934 166046 528002 166102
rect 528058 166046 528126 166102
rect 528182 166046 558474 166102
rect 558530 166046 558598 166102
rect 558654 166046 558722 166102
rect 558778 166046 558846 166102
rect 558902 166046 589194 166102
rect 589250 166046 589318 166102
rect 589374 166046 589442 166102
rect 589498 166046 589566 166102
rect 589622 166046 596496 166102
rect 596552 166046 596620 166102
rect 596676 166046 596744 166102
rect 596800 166046 596868 166102
rect 596924 166046 597980 166102
rect -1916 165978 597980 166046
rect -1916 165922 -860 165978
rect -804 165922 -736 165978
rect -680 165922 -612 165978
rect -556 165922 -488 165978
rect -432 165922 5514 165978
rect 5570 165922 5638 165978
rect 5694 165922 5762 165978
rect 5818 165922 5886 165978
rect 5942 165922 36234 165978
rect 36290 165922 36358 165978
rect 36414 165922 36482 165978
rect 36538 165922 36606 165978
rect 36662 165922 66954 165978
rect 67010 165922 67078 165978
rect 67134 165922 67202 165978
rect 67258 165922 67326 165978
rect 67382 165922 97674 165978
rect 97730 165922 97798 165978
rect 97854 165922 97922 165978
rect 97978 165922 98046 165978
rect 98102 165922 128394 165978
rect 128450 165922 128518 165978
rect 128574 165922 128642 165978
rect 128698 165922 128766 165978
rect 128822 165922 159114 165978
rect 159170 165922 159238 165978
rect 159294 165922 159362 165978
rect 159418 165922 159486 165978
rect 159542 165922 189834 165978
rect 189890 165922 189958 165978
rect 190014 165922 190082 165978
rect 190138 165922 190206 165978
rect 190262 165922 220554 165978
rect 220610 165922 220678 165978
rect 220734 165922 220802 165978
rect 220858 165922 220926 165978
rect 220982 165922 251274 165978
rect 251330 165922 251398 165978
rect 251454 165922 251522 165978
rect 251578 165922 251646 165978
rect 251702 165922 272518 165978
rect 272574 165922 272642 165978
rect 272698 165922 303238 165978
rect 303294 165922 303362 165978
rect 303418 165922 343434 165978
rect 343490 165922 343558 165978
rect 343614 165922 343682 165978
rect 343738 165922 343806 165978
rect 343862 165922 374154 165978
rect 374210 165922 374278 165978
rect 374334 165922 374402 165978
rect 374458 165922 374526 165978
rect 374582 165922 404874 165978
rect 404930 165922 404998 165978
rect 405054 165922 405122 165978
rect 405178 165922 405246 165978
rect 405302 165922 435594 165978
rect 435650 165922 435718 165978
rect 435774 165922 435842 165978
rect 435898 165922 435966 165978
rect 436022 165922 466314 165978
rect 466370 165922 466438 165978
rect 466494 165922 466562 165978
rect 466618 165922 466686 165978
rect 466742 165922 497034 165978
rect 497090 165922 497158 165978
rect 497214 165922 497282 165978
rect 497338 165922 497406 165978
rect 497462 165922 527754 165978
rect 527810 165922 527878 165978
rect 527934 165922 528002 165978
rect 528058 165922 528126 165978
rect 528182 165922 558474 165978
rect 558530 165922 558598 165978
rect 558654 165922 558722 165978
rect 558778 165922 558846 165978
rect 558902 165922 589194 165978
rect 589250 165922 589318 165978
rect 589374 165922 589442 165978
rect 589498 165922 589566 165978
rect 589622 165922 596496 165978
rect 596552 165922 596620 165978
rect 596676 165922 596744 165978
rect 596800 165922 596868 165978
rect 596924 165922 597980 165978
rect -1916 165826 597980 165922
rect -1916 154350 597980 154446
rect -1916 154294 -1820 154350
rect -1764 154294 -1696 154350
rect -1640 154294 -1572 154350
rect -1516 154294 -1448 154350
rect -1392 154294 9234 154350
rect 9290 154294 9358 154350
rect 9414 154294 9482 154350
rect 9538 154294 9606 154350
rect 9662 154294 39954 154350
rect 40010 154294 40078 154350
rect 40134 154294 40202 154350
rect 40258 154294 40326 154350
rect 40382 154294 70674 154350
rect 70730 154294 70798 154350
rect 70854 154294 70922 154350
rect 70978 154294 71046 154350
rect 71102 154294 101394 154350
rect 101450 154294 101518 154350
rect 101574 154294 101642 154350
rect 101698 154294 101766 154350
rect 101822 154294 132114 154350
rect 132170 154294 132238 154350
rect 132294 154294 132362 154350
rect 132418 154294 132486 154350
rect 132542 154294 162834 154350
rect 162890 154294 162958 154350
rect 163014 154294 163082 154350
rect 163138 154294 163206 154350
rect 163262 154294 193554 154350
rect 193610 154294 193678 154350
rect 193734 154294 193802 154350
rect 193858 154294 193926 154350
rect 193982 154294 224274 154350
rect 224330 154294 224398 154350
rect 224454 154294 224522 154350
rect 224578 154294 224646 154350
rect 224702 154294 254994 154350
rect 255050 154294 255118 154350
rect 255174 154294 255242 154350
rect 255298 154294 255366 154350
rect 255422 154294 287878 154350
rect 287934 154294 288002 154350
rect 288058 154294 318598 154350
rect 318654 154294 318722 154350
rect 318778 154294 347154 154350
rect 347210 154294 347278 154350
rect 347334 154294 347402 154350
rect 347458 154294 347526 154350
rect 347582 154294 377874 154350
rect 377930 154294 377998 154350
rect 378054 154294 378122 154350
rect 378178 154294 378246 154350
rect 378302 154294 408594 154350
rect 408650 154294 408718 154350
rect 408774 154294 408842 154350
rect 408898 154294 408966 154350
rect 409022 154294 439314 154350
rect 439370 154294 439438 154350
rect 439494 154294 439562 154350
rect 439618 154294 439686 154350
rect 439742 154294 470034 154350
rect 470090 154294 470158 154350
rect 470214 154294 470282 154350
rect 470338 154294 470406 154350
rect 470462 154294 500754 154350
rect 500810 154294 500878 154350
rect 500934 154294 501002 154350
rect 501058 154294 501126 154350
rect 501182 154294 531474 154350
rect 531530 154294 531598 154350
rect 531654 154294 531722 154350
rect 531778 154294 531846 154350
rect 531902 154294 562194 154350
rect 562250 154294 562318 154350
rect 562374 154294 562442 154350
rect 562498 154294 562566 154350
rect 562622 154294 592914 154350
rect 592970 154294 593038 154350
rect 593094 154294 593162 154350
rect 593218 154294 593286 154350
rect 593342 154294 597456 154350
rect 597512 154294 597580 154350
rect 597636 154294 597704 154350
rect 597760 154294 597828 154350
rect 597884 154294 597980 154350
rect -1916 154226 597980 154294
rect -1916 154170 -1820 154226
rect -1764 154170 -1696 154226
rect -1640 154170 -1572 154226
rect -1516 154170 -1448 154226
rect -1392 154170 9234 154226
rect 9290 154170 9358 154226
rect 9414 154170 9482 154226
rect 9538 154170 9606 154226
rect 9662 154170 39954 154226
rect 40010 154170 40078 154226
rect 40134 154170 40202 154226
rect 40258 154170 40326 154226
rect 40382 154170 70674 154226
rect 70730 154170 70798 154226
rect 70854 154170 70922 154226
rect 70978 154170 71046 154226
rect 71102 154170 101394 154226
rect 101450 154170 101518 154226
rect 101574 154170 101642 154226
rect 101698 154170 101766 154226
rect 101822 154170 132114 154226
rect 132170 154170 132238 154226
rect 132294 154170 132362 154226
rect 132418 154170 132486 154226
rect 132542 154170 162834 154226
rect 162890 154170 162958 154226
rect 163014 154170 163082 154226
rect 163138 154170 163206 154226
rect 163262 154170 193554 154226
rect 193610 154170 193678 154226
rect 193734 154170 193802 154226
rect 193858 154170 193926 154226
rect 193982 154170 224274 154226
rect 224330 154170 224398 154226
rect 224454 154170 224522 154226
rect 224578 154170 224646 154226
rect 224702 154170 254994 154226
rect 255050 154170 255118 154226
rect 255174 154170 255242 154226
rect 255298 154170 255366 154226
rect 255422 154170 287878 154226
rect 287934 154170 288002 154226
rect 288058 154170 318598 154226
rect 318654 154170 318722 154226
rect 318778 154170 347154 154226
rect 347210 154170 347278 154226
rect 347334 154170 347402 154226
rect 347458 154170 347526 154226
rect 347582 154170 377874 154226
rect 377930 154170 377998 154226
rect 378054 154170 378122 154226
rect 378178 154170 378246 154226
rect 378302 154170 408594 154226
rect 408650 154170 408718 154226
rect 408774 154170 408842 154226
rect 408898 154170 408966 154226
rect 409022 154170 439314 154226
rect 439370 154170 439438 154226
rect 439494 154170 439562 154226
rect 439618 154170 439686 154226
rect 439742 154170 470034 154226
rect 470090 154170 470158 154226
rect 470214 154170 470282 154226
rect 470338 154170 470406 154226
rect 470462 154170 500754 154226
rect 500810 154170 500878 154226
rect 500934 154170 501002 154226
rect 501058 154170 501126 154226
rect 501182 154170 531474 154226
rect 531530 154170 531598 154226
rect 531654 154170 531722 154226
rect 531778 154170 531846 154226
rect 531902 154170 562194 154226
rect 562250 154170 562318 154226
rect 562374 154170 562442 154226
rect 562498 154170 562566 154226
rect 562622 154170 592914 154226
rect 592970 154170 593038 154226
rect 593094 154170 593162 154226
rect 593218 154170 593286 154226
rect 593342 154170 597456 154226
rect 597512 154170 597580 154226
rect 597636 154170 597704 154226
rect 597760 154170 597828 154226
rect 597884 154170 597980 154226
rect -1916 154102 597980 154170
rect -1916 154046 -1820 154102
rect -1764 154046 -1696 154102
rect -1640 154046 -1572 154102
rect -1516 154046 -1448 154102
rect -1392 154046 9234 154102
rect 9290 154046 9358 154102
rect 9414 154046 9482 154102
rect 9538 154046 9606 154102
rect 9662 154046 39954 154102
rect 40010 154046 40078 154102
rect 40134 154046 40202 154102
rect 40258 154046 40326 154102
rect 40382 154046 70674 154102
rect 70730 154046 70798 154102
rect 70854 154046 70922 154102
rect 70978 154046 71046 154102
rect 71102 154046 101394 154102
rect 101450 154046 101518 154102
rect 101574 154046 101642 154102
rect 101698 154046 101766 154102
rect 101822 154046 132114 154102
rect 132170 154046 132238 154102
rect 132294 154046 132362 154102
rect 132418 154046 132486 154102
rect 132542 154046 162834 154102
rect 162890 154046 162958 154102
rect 163014 154046 163082 154102
rect 163138 154046 163206 154102
rect 163262 154046 193554 154102
rect 193610 154046 193678 154102
rect 193734 154046 193802 154102
rect 193858 154046 193926 154102
rect 193982 154046 224274 154102
rect 224330 154046 224398 154102
rect 224454 154046 224522 154102
rect 224578 154046 224646 154102
rect 224702 154046 254994 154102
rect 255050 154046 255118 154102
rect 255174 154046 255242 154102
rect 255298 154046 255366 154102
rect 255422 154046 287878 154102
rect 287934 154046 288002 154102
rect 288058 154046 318598 154102
rect 318654 154046 318722 154102
rect 318778 154046 347154 154102
rect 347210 154046 347278 154102
rect 347334 154046 347402 154102
rect 347458 154046 347526 154102
rect 347582 154046 377874 154102
rect 377930 154046 377998 154102
rect 378054 154046 378122 154102
rect 378178 154046 378246 154102
rect 378302 154046 408594 154102
rect 408650 154046 408718 154102
rect 408774 154046 408842 154102
rect 408898 154046 408966 154102
rect 409022 154046 439314 154102
rect 439370 154046 439438 154102
rect 439494 154046 439562 154102
rect 439618 154046 439686 154102
rect 439742 154046 470034 154102
rect 470090 154046 470158 154102
rect 470214 154046 470282 154102
rect 470338 154046 470406 154102
rect 470462 154046 500754 154102
rect 500810 154046 500878 154102
rect 500934 154046 501002 154102
rect 501058 154046 501126 154102
rect 501182 154046 531474 154102
rect 531530 154046 531598 154102
rect 531654 154046 531722 154102
rect 531778 154046 531846 154102
rect 531902 154046 562194 154102
rect 562250 154046 562318 154102
rect 562374 154046 562442 154102
rect 562498 154046 562566 154102
rect 562622 154046 592914 154102
rect 592970 154046 593038 154102
rect 593094 154046 593162 154102
rect 593218 154046 593286 154102
rect 593342 154046 597456 154102
rect 597512 154046 597580 154102
rect 597636 154046 597704 154102
rect 597760 154046 597828 154102
rect 597884 154046 597980 154102
rect -1916 153978 597980 154046
rect -1916 153922 -1820 153978
rect -1764 153922 -1696 153978
rect -1640 153922 -1572 153978
rect -1516 153922 -1448 153978
rect -1392 153922 9234 153978
rect 9290 153922 9358 153978
rect 9414 153922 9482 153978
rect 9538 153922 9606 153978
rect 9662 153922 39954 153978
rect 40010 153922 40078 153978
rect 40134 153922 40202 153978
rect 40258 153922 40326 153978
rect 40382 153922 70674 153978
rect 70730 153922 70798 153978
rect 70854 153922 70922 153978
rect 70978 153922 71046 153978
rect 71102 153922 101394 153978
rect 101450 153922 101518 153978
rect 101574 153922 101642 153978
rect 101698 153922 101766 153978
rect 101822 153922 132114 153978
rect 132170 153922 132238 153978
rect 132294 153922 132362 153978
rect 132418 153922 132486 153978
rect 132542 153922 162834 153978
rect 162890 153922 162958 153978
rect 163014 153922 163082 153978
rect 163138 153922 163206 153978
rect 163262 153922 193554 153978
rect 193610 153922 193678 153978
rect 193734 153922 193802 153978
rect 193858 153922 193926 153978
rect 193982 153922 224274 153978
rect 224330 153922 224398 153978
rect 224454 153922 224522 153978
rect 224578 153922 224646 153978
rect 224702 153922 254994 153978
rect 255050 153922 255118 153978
rect 255174 153922 255242 153978
rect 255298 153922 255366 153978
rect 255422 153922 287878 153978
rect 287934 153922 288002 153978
rect 288058 153922 318598 153978
rect 318654 153922 318722 153978
rect 318778 153922 347154 153978
rect 347210 153922 347278 153978
rect 347334 153922 347402 153978
rect 347458 153922 347526 153978
rect 347582 153922 377874 153978
rect 377930 153922 377998 153978
rect 378054 153922 378122 153978
rect 378178 153922 378246 153978
rect 378302 153922 408594 153978
rect 408650 153922 408718 153978
rect 408774 153922 408842 153978
rect 408898 153922 408966 153978
rect 409022 153922 439314 153978
rect 439370 153922 439438 153978
rect 439494 153922 439562 153978
rect 439618 153922 439686 153978
rect 439742 153922 470034 153978
rect 470090 153922 470158 153978
rect 470214 153922 470282 153978
rect 470338 153922 470406 153978
rect 470462 153922 500754 153978
rect 500810 153922 500878 153978
rect 500934 153922 501002 153978
rect 501058 153922 501126 153978
rect 501182 153922 531474 153978
rect 531530 153922 531598 153978
rect 531654 153922 531722 153978
rect 531778 153922 531846 153978
rect 531902 153922 562194 153978
rect 562250 153922 562318 153978
rect 562374 153922 562442 153978
rect 562498 153922 562566 153978
rect 562622 153922 592914 153978
rect 592970 153922 593038 153978
rect 593094 153922 593162 153978
rect 593218 153922 593286 153978
rect 593342 153922 597456 153978
rect 597512 153922 597580 153978
rect 597636 153922 597704 153978
rect 597760 153922 597828 153978
rect 597884 153922 597980 153978
rect -1916 153826 597980 153922
rect -1916 148350 597980 148446
rect -1916 148294 -860 148350
rect -804 148294 -736 148350
rect -680 148294 -612 148350
rect -556 148294 -488 148350
rect -432 148294 5514 148350
rect 5570 148294 5638 148350
rect 5694 148294 5762 148350
rect 5818 148294 5886 148350
rect 5942 148294 36234 148350
rect 36290 148294 36358 148350
rect 36414 148294 36482 148350
rect 36538 148294 36606 148350
rect 36662 148294 66954 148350
rect 67010 148294 67078 148350
rect 67134 148294 67202 148350
rect 67258 148294 67326 148350
rect 67382 148294 97674 148350
rect 97730 148294 97798 148350
rect 97854 148294 97922 148350
rect 97978 148294 98046 148350
rect 98102 148294 128394 148350
rect 128450 148294 128518 148350
rect 128574 148294 128642 148350
rect 128698 148294 128766 148350
rect 128822 148294 159114 148350
rect 159170 148294 159238 148350
rect 159294 148294 159362 148350
rect 159418 148294 159486 148350
rect 159542 148294 189834 148350
rect 189890 148294 189958 148350
rect 190014 148294 190082 148350
rect 190138 148294 190206 148350
rect 190262 148294 220554 148350
rect 220610 148294 220678 148350
rect 220734 148294 220802 148350
rect 220858 148294 220926 148350
rect 220982 148294 251274 148350
rect 251330 148294 251398 148350
rect 251454 148294 251522 148350
rect 251578 148294 251646 148350
rect 251702 148294 272518 148350
rect 272574 148294 272642 148350
rect 272698 148294 303238 148350
rect 303294 148294 303362 148350
rect 303418 148294 343434 148350
rect 343490 148294 343558 148350
rect 343614 148294 343682 148350
rect 343738 148294 343806 148350
rect 343862 148294 374154 148350
rect 374210 148294 374278 148350
rect 374334 148294 374402 148350
rect 374458 148294 374526 148350
rect 374582 148294 404874 148350
rect 404930 148294 404998 148350
rect 405054 148294 405122 148350
rect 405178 148294 405246 148350
rect 405302 148294 435594 148350
rect 435650 148294 435718 148350
rect 435774 148294 435842 148350
rect 435898 148294 435966 148350
rect 436022 148294 466314 148350
rect 466370 148294 466438 148350
rect 466494 148294 466562 148350
rect 466618 148294 466686 148350
rect 466742 148294 497034 148350
rect 497090 148294 497158 148350
rect 497214 148294 497282 148350
rect 497338 148294 497406 148350
rect 497462 148294 527754 148350
rect 527810 148294 527878 148350
rect 527934 148294 528002 148350
rect 528058 148294 528126 148350
rect 528182 148294 558474 148350
rect 558530 148294 558598 148350
rect 558654 148294 558722 148350
rect 558778 148294 558846 148350
rect 558902 148294 589194 148350
rect 589250 148294 589318 148350
rect 589374 148294 589442 148350
rect 589498 148294 589566 148350
rect 589622 148294 596496 148350
rect 596552 148294 596620 148350
rect 596676 148294 596744 148350
rect 596800 148294 596868 148350
rect 596924 148294 597980 148350
rect -1916 148226 597980 148294
rect -1916 148170 -860 148226
rect -804 148170 -736 148226
rect -680 148170 -612 148226
rect -556 148170 -488 148226
rect -432 148170 5514 148226
rect 5570 148170 5638 148226
rect 5694 148170 5762 148226
rect 5818 148170 5886 148226
rect 5942 148170 36234 148226
rect 36290 148170 36358 148226
rect 36414 148170 36482 148226
rect 36538 148170 36606 148226
rect 36662 148170 66954 148226
rect 67010 148170 67078 148226
rect 67134 148170 67202 148226
rect 67258 148170 67326 148226
rect 67382 148170 97674 148226
rect 97730 148170 97798 148226
rect 97854 148170 97922 148226
rect 97978 148170 98046 148226
rect 98102 148170 128394 148226
rect 128450 148170 128518 148226
rect 128574 148170 128642 148226
rect 128698 148170 128766 148226
rect 128822 148170 159114 148226
rect 159170 148170 159238 148226
rect 159294 148170 159362 148226
rect 159418 148170 159486 148226
rect 159542 148170 189834 148226
rect 189890 148170 189958 148226
rect 190014 148170 190082 148226
rect 190138 148170 190206 148226
rect 190262 148170 220554 148226
rect 220610 148170 220678 148226
rect 220734 148170 220802 148226
rect 220858 148170 220926 148226
rect 220982 148170 251274 148226
rect 251330 148170 251398 148226
rect 251454 148170 251522 148226
rect 251578 148170 251646 148226
rect 251702 148170 272518 148226
rect 272574 148170 272642 148226
rect 272698 148170 303238 148226
rect 303294 148170 303362 148226
rect 303418 148170 343434 148226
rect 343490 148170 343558 148226
rect 343614 148170 343682 148226
rect 343738 148170 343806 148226
rect 343862 148170 374154 148226
rect 374210 148170 374278 148226
rect 374334 148170 374402 148226
rect 374458 148170 374526 148226
rect 374582 148170 404874 148226
rect 404930 148170 404998 148226
rect 405054 148170 405122 148226
rect 405178 148170 405246 148226
rect 405302 148170 435594 148226
rect 435650 148170 435718 148226
rect 435774 148170 435842 148226
rect 435898 148170 435966 148226
rect 436022 148170 466314 148226
rect 466370 148170 466438 148226
rect 466494 148170 466562 148226
rect 466618 148170 466686 148226
rect 466742 148170 497034 148226
rect 497090 148170 497158 148226
rect 497214 148170 497282 148226
rect 497338 148170 497406 148226
rect 497462 148170 527754 148226
rect 527810 148170 527878 148226
rect 527934 148170 528002 148226
rect 528058 148170 528126 148226
rect 528182 148170 558474 148226
rect 558530 148170 558598 148226
rect 558654 148170 558722 148226
rect 558778 148170 558846 148226
rect 558902 148170 589194 148226
rect 589250 148170 589318 148226
rect 589374 148170 589442 148226
rect 589498 148170 589566 148226
rect 589622 148170 596496 148226
rect 596552 148170 596620 148226
rect 596676 148170 596744 148226
rect 596800 148170 596868 148226
rect 596924 148170 597980 148226
rect -1916 148102 597980 148170
rect -1916 148046 -860 148102
rect -804 148046 -736 148102
rect -680 148046 -612 148102
rect -556 148046 -488 148102
rect -432 148046 5514 148102
rect 5570 148046 5638 148102
rect 5694 148046 5762 148102
rect 5818 148046 5886 148102
rect 5942 148046 36234 148102
rect 36290 148046 36358 148102
rect 36414 148046 36482 148102
rect 36538 148046 36606 148102
rect 36662 148046 66954 148102
rect 67010 148046 67078 148102
rect 67134 148046 67202 148102
rect 67258 148046 67326 148102
rect 67382 148046 97674 148102
rect 97730 148046 97798 148102
rect 97854 148046 97922 148102
rect 97978 148046 98046 148102
rect 98102 148046 128394 148102
rect 128450 148046 128518 148102
rect 128574 148046 128642 148102
rect 128698 148046 128766 148102
rect 128822 148046 159114 148102
rect 159170 148046 159238 148102
rect 159294 148046 159362 148102
rect 159418 148046 159486 148102
rect 159542 148046 189834 148102
rect 189890 148046 189958 148102
rect 190014 148046 190082 148102
rect 190138 148046 190206 148102
rect 190262 148046 220554 148102
rect 220610 148046 220678 148102
rect 220734 148046 220802 148102
rect 220858 148046 220926 148102
rect 220982 148046 251274 148102
rect 251330 148046 251398 148102
rect 251454 148046 251522 148102
rect 251578 148046 251646 148102
rect 251702 148046 272518 148102
rect 272574 148046 272642 148102
rect 272698 148046 303238 148102
rect 303294 148046 303362 148102
rect 303418 148046 343434 148102
rect 343490 148046 343558 148102
rect 343614 148046 343682 148102
rect 343738 148046 343806 148102
rect 343862 148046 374154 148102
rect 374210 148046 374278 148102
rect 374334 148046 374402 148102
rect 374458 148046 374526 148102
rect 374582 148046 404874 148102
rect 404930 148046 404998 148102
rect 405054 148046 405122 148102
rect 405178 148046 405246 148102
rect 405302 148046 435594 148102
rect 435650 148046 435718 148102
rect 435774 148046 435842 148102
rect 435898 148046 435966 148102
rect 436022 148046 466314 148102
rect 466370 148046 466438 148102
rect 466494 148046 466562 148102
rect 466618 148046 466686 148102
rect 466742 148046 497034 148102
rect 497090 148046 497158 148102
rect 497214 148046 497282 148102
rect 497338 148046 497406 148102
rect 497462 148046 527754 148102
rect 527810 148046 527878 148102
rect 527934 148046 528002 148102
rect 528058 148046 528126 148102
rect 528182 148046 558474 148102
rect 558530 148046 558598 148102
rect 558654 148046 558722 148102
rect 558778 148046 558846 148102
rect 558902 148046 589194 148102
rect 589250 148046 589318 148102
rect 589374 148046 589442 148102
rect 589498 148046 589566 148102
rect 589622 148046 596496 148102
rect 596552 148046 596620 148102
rect 596676 148046 596744 148102
rect 596800 148046 596868 148102
rect 596924 148046 597980 148102
rect -1916 147978 597980 148046
rect -1916 147922 -860 147978
rect -804 147922 -736 147978
rect -680 147922 -612 147978
rect -556 147922 -488 147978
rect -432 147922 5514 147978
rect 5570 147922 5638 147978
rect 5694 147922 5762 147978
rect 5818 147922 5886 147978
rect 5942 147922 36234 147978
rect 36290 147922 36358 147978
rect 36414 147922 36482 147978
rect 36538 147922 36606 147978
rect 36662 147922 66954 147978
rect 67010 147922 67078 147978
rect 67134 147922 67202 147978
rect 67258 147922 67326 147978
rect 67382 147922 97674 147978
rect 97730 147922 97798 147978
rect 97854 147922 97922 147978
rect 97978 147922 98046 147978
rect 98102 147922 128394 147978
rect 128450 147922 128518 147978
rect 128574 147922 128642 147978
rect 128698 147922 128766 147978
rect 128822 147922 159114 147978
rect 159170 147922 159238 147978
rect 159294 147922 159362 147978
rect 159418 147922 159486 147978
rect 159542 147922 189834 147978
rect 189890 147922 189958 147978
rect 190014 147922 190082 147978
rect 190138 147922 190206 147978
rect 190262 147922 220554 147978
rect 220610 147922 220678 147978
rect 220734 147922 220802 147978
rect 220858 147922 220926 147978
rect 220982 147922 251274 147978
rect 251330 147922 251398 147978
rect 251454 147922 251522 147978
rect 251578 147922 251646 147978
rect 251702 147922 272518 147978
rect 272574 147922 272642 147978
rect 272698 147922 303238 147978
rect 303294 147922 303362 147978
rect 303418 147922 343434 147978
rect 343490 147922 343558 147978
rect 343614 147922 343682 147978
rect 343738 147922 343806 147978
rect 343862 147922 374154 147978
rect 374210 147922 374278 147978
rect 374334 147922 374402 147978
rect 374458 147922 374526 147978
rect 374582 147922 404874 147978
rect 404930 147922 404998 147978
rect 405054 147922 405122 147978
rect 405178 147922 405246 147978
rect 405302 147922 435594 147978
rect 435650 147922 435718 147978
rect 435774 147922 435842 147978
rect 435898 147922 435966 147978
rect 436022 147922 466314 147978
rect 466370 147922 466438 147978
rect 466494 147922 466562 147978
rect 466618 147922 466686 147978
rect 466742 147922 497034 147978
rect 497090 147922 497158 147978
rect 497214 147922 497282 147978
rect 497338 147922 497406 147978
rect 497462 147922 527754 147978
rect 527810 147922 527878 147978
rect 527934 147922 528002 147978
rect 528058 147922 528126 147978
rect 528182 147922 558474 147978
rect 558530 147922 558598 147978
rect 558654 147922 558722 147978
rect 558778 147922 558846 147978
rect 558902 147922 589194 147978
rect 589250 147922 589318 147978
rect 589374 147922 589442 147978
rect 589498 147922 589566 147978
rect 589622 147922 596496 147978
rect 596552 147922 596620 147978
rect 596676 147922 596744 147978
rect 596800 147922 596868 147978
rect 596924 147922 597980 147978
rect -1916 147826 597980 147922
rect 141916 137818 263860 137834
rect 141916 137762 141932 137818
rect 141988 137762 263788 137818
rect 263844 137762 263860 137818
rect 141916 137746 263860 137762
rect -1916 136350 597980 136446
rect -1916 136294 -1820 136350
rect -1764 136294 -1696 136350
rect -1640 136294 -1572 136350
rect -1516 136294 -1448 136350
rect -1392 136294 9234 136350
rect 9290 136294 9358 136350
rect 9414 136294 9482 136350
rect 9538 136294 9606 136350
rect 9662 136294 39878 136350
rect 39934 136294 40002 136350
rect 40058 136294 70674 136350
rect 70730 136294 70798 136350
rect 70854 136294 70922 136350
rect 70978 136294 71046 136350
rect 71102 136294 101878 136350
rect 101934 136294 102002 136350
rect 102058 136294 132114 136350
rect 132170 136294 132238 136350
rect 132294 136294 132362 136350
rect 132418 136294 132486 136350
rect 132542 136294 162834 136350
rect 162890 136294 162958 136350
rect 163014 136294 163082 136350
rect 163138 136294 163206 136350
rect 163262 136294 163878 136350
rect 163934 136294 164002 136350
rect 164058 136294 193554 136350
rect 193610 136294 193678 136350
rect 193734 136294 193802 136350
rect 193858 136294 193926 136350
rect 193982 136294 224274 136350
rect 224330 136294 224398 136350
rect 224454 136294 224522 136350
rect 224578 136294 224646 136350
rect 224702 136294 225878 136350
rect 225934 136294 226002 136350
rect 226058 136294 254994 136350
rect 255050 136294 255118 136350
rect 255174 136294 255242 136350
rect 255298 136294 255366 136350
rect 255422 136294 287878 136350
rect 287934 136294 288002 136350
rect 288058 136294 318598 136350
rect 318654 136294 318722 136350
rect 318778 136294 347154 136350
rect 347210 136294 347278 136350
rect 347334 136294 347402 136350
rect 347458 136294 347526 136350
rect 347582 136294 371878 136350
rect 371934 136294 372002 136350
rect 372058 136294 377874 136350
rect 377930 136294 377998 136350
rect 378054 136294 378122 136350
rect 378178 136294 378246 136350
rect 378302 136294 408594 136350
rect 408650 136294 408718 136350
rect 408774 136294 408842 136350
rect 408898 136294 408966 136350
rect 409022 136294 433878 136350
rect 433934 136294 434002 136350
rect 434058 136294 439314 136350
rect 439370 136294 439438 136350
rect 439494 136294 439562 136350
rect 439618 136294 439686 136350
rect 439742 136294 470034 136350
rect 470090 136294 470158 136350
rect 470214 136294 470282 136350
rect 470338 136294 470406 136350
rect 470462 136294 495878 136350
rect 495934 136294 496002 136350
rect 496058 136294 500754 136350
rect 500810 136294 500878 136350
rect 500934 136294 501002 136350
rect 501058 136294 501126 136350
rect 501182 136294 531474 136350
rect 531530 136294 531598 136350
rect 531654 136294 531722 136350
rect 531778 136294 531846 136350
rect 531902 136294 557878 136350
rect 557934 136294 558002 136350
rect 558058 136294 562194 136350
rect 562250 136294 562318 136350
rect 562374 136294 562442 136350
rect 562498 136294 562566 136350
rect 562622 136294 592914 136350
rect 592970 136294 593038 136350
rect 593094 136294 593162 136350
rect 593218 136294 593286 136350
rect 593342 136294 597456 136350
rect 597512 136294 597580 136350
rect 597636 136294 597704 136350
rect 597760 136294 597828 136350
rect 597884 136294 597980 136350
rect -1916 136226 597980 136294
rect -1916 136170 -1820 136226
rect -1764 136170 -1696 136226
rect -1640 136170 -1572 136226
rect -1516 136170 -1448 136226
rect -1392 136170 9234 136226
rect 9290 136170 9358 136226
rect 9414 136170 9482 136226
rect 9538 136170 9606 136226
rect 9662 136170 39878 136226
rect 39934 136170 40002 136226
rect 40058 136170 70674 136226
rect 70730 136170 70798 136226
rect 70854 136170 70922 136226
rect 70978 136170 71046 136226
rect 71102 136170 101878 136226
rect 101934 136170 102002 136226
rect 102058 136170 132114 136226
rect 132170 136170 132238 136226
rect 132294 136170 132362 136226
rect 132418 136170 132486 136226
rect 132542 136170 162834 136226
rect 162890 136170 162958 136226
rect 163014 136170 163082 136226
rect 163138 136170 163206 136226
rect 163262 136170 163878 136226
rect 163934 136170 164002 136226
rect 164058 136170 193554 136226
rect 193610 136170 193678 136226
rect 193734 136170 193802 136226
rect 193858 136170 193926 136226
rect 193982 136170 224274 136226
rect 224330 136170 224398 136226
rect 224454 136170 224522 136226
rect 224578 136170 224646 136226
rect 224702 136170 225878 136226
rect 225934 136170 226002 136226
rect 226058 136170 254994 136226
rect 255050 136170 255118 136226
rect 255174 136170 255242 136226
rect 255298 136170 255366 136226
rect 255422 136170 287878 136226
rect 287934 136170 288002 136226
rect 288058 136170 318598 136226
rect 318654 136170 318722 136226
rect 318778 136170 347154 136226
rect 347210 136170 347278 136226
rect 347334 136170 347402 136226
rect 347458 136170 347526 136226
rect 347582 136170 371878 136226
rect 371934 136170 372002 136226
rect 372058 136170 377874 136226
rect 377930 136170 377998 136226
rect 378054 136170 378122 136226
rect 378178 136170 378246 136226
rect 378302 136170 408594 136226
rect 408650 136170 408718 136226
rect 408774 136170 408842 136226
rect 408898 136170 408966 136226
rect 409022 136170 433878 136226
rect 433934 136170 434002 136226
rect 434058 136170 439314 136226
rect 439370 136170 439438 136226
rect 439494 136170 439562 136226
rect 439618 136170 439686 136226
rect 439742 136170 470034 136226
rect 470090 136170 470158 136226
rect 470214 136170 470282 136226
rect 470338 136170 470406 136226
rect 470462 136170 495878 136226
rect 495934 136170 496002 136226
rect 496058 136170 500754 136226
rect 500810 136170 500878 136226
rect 500934 136170 501002 136226
rect 501058 136170 501126 136226
rect 501182 136170 531474 136226
rect 531530 136170 531598 136226
rect 531654 136170 531722 136226
rect 531778 136170 531846 136226
rect 531902 136170 557878 136226
rect 557934 136170 558002 136226
rect 558058 136170 562194 136226
rect 562250 136170 562318 136226
rect 562374 136170 562442 136226
rect 562498 136170 562566 136226
rect 562622 136170 592914 136226
rect 592970 136170 593038 136226
rect 593094 136170 593162 136226
rect 593218 136170 593286 136226
rect 593342 136170 597456 136226
rect 597512 136170 597580 136226
rect 597636 136170 597704 136226
rect 597760 136170 597828 136226
rect 597884 136170 597980 136226
rect -1916 136102 597980 136170
rect -1916 136046 -1820 136102
rect -1764 136046 -1696 136102
rect -1640 136046 -1572 136102
rect -1516 136046 -1448 136102
rect -1392 136046 9234 136102
rect 9290 136046 9358 136102
rect 9414 136046 9482 136102
rect 9538 136046 9606 136102
rect 9662 136046 39878 136102
rect 39934 136046 40002 136102
rect 40058 136046 70674 136102
rect 70730 136046 70798 136102
rect 70854 136046 70922 136102
rect 70978 136046 71046 136102
rect 71102 136046 101878 136102
rect 101934 136046 102002 136102
rect 102058 136046 132114 136102
rect 132170 136046 132238 136102
rect 132294 136046 132362 136102
rect 132418 136046 132486 136102
rect 132542 136046 162834 136102
rect 162890 136046 162958 136102
rect 163014 136046 163082 136102
rect 163138 136046 163206 136102
rect 163262 136046 163878 136102
rect 163934 136046 164002 136102
rect 164058 136046 193554 136102
rect 193610 136046 193678 136102
rect 193734 136046 193802 136102
rect 193858 136046 193926 136102
rect 193982 136046 224274 136102
rect 224330 136046 224398 136102
rect 224454 136046 224522 136102
rect 224578 136046 224646 136102
rect 224702 136046 225878 136102
rect 225934 136046 226002 136102
rect 226058 136046 254994 136102
rect 255050 136046 255118 136102
rect 255174 136046 255242 136102
rect 255298 136046 255366 136102
rect 255422 136046 287878 136102
rect 287934 136046 288002 136102
rect 288058 136046 318598 136102
rect 318654 136046 318722 136102
rect 318778 136046 347154 136102
rect 347210 136046 347278 136102
rect 347334 136046 347402 136102
rect 347458 136046 347526 136102
rect 347582 136046 371878 136102
rect 371934 136046 372002 136102
rect 372058 136046 377874 136102
rect 377930 136046 377998 136102
rect 378054 136046 378122 136102
rect 378178 136046 378246 136102
rect 378302 136046 408594 136102
rect 408650 136046 408718 136102
rect 408774 136046 408842 136102
rect 408898 136046 408966 136102
rect 409022 136046 433878 136102
rect 433934 136046 434002 136102
rect 434058 136046 439314 136102
rect 439370 136046 439438 136102
rect 439494 136046 439562 136102
rect 439618 136046 439686 136102
rect 439742 136046 470034 136102
rect 470090 136046 470158 136102
rect 470214 136046 470282 136102
rect 470338 136046 470406 136102
rect 470462 136046 495878 136102
rect 495934 136046 496002 136102
rect 496058 136046 500754 136102
rect 500810 136046 500878 136102
rect 500934 136046 501002 136102
rect 501058 136046 501126 136102
rect 501182 136046 531474 136102
rect 531530 136046 531598 136102
rect 531654 136046 531722 136102
rect 531778 136046 531846 136102
rect 531902 136046 557878 136102
rect 557934 136046 558002 136102
rect 558058 136046 562194 136102
rect 562250 136046 562318 136102
rect 562374 136046 562442 136102
rect 562498 136046 562566 136102
rect 562622 136046 592914 136102
rect 592970 136046 593038 136102
rect 593094 136046 593162 136102
rect 593218 136046 593286 136102
rect 593342 136046 597456 136102
rect 597512 136046 597580 136102
rect 597636 136046 597704 136102
rect 597760 136046 597828 136102
rect 597884 136046 597980 136102
rect -1916 135978 597980 136046
rect -1916 135922 -1820 135978
rect -1764 135922 -1696 135978
rect -1640 135922 -1572 135978
rect -1516 135922 -1448 135978
rect -1392 135922 9234 135978
rect 9290 135922 9358 135978
rect 9414 135922 9482 135978
rect 9538 135922 9606 135978
rect 9662 135922 39878 135978
rect 39934 135922 40002 135978
rect 40058 135922 70674 135978
rect 70730 135922 70798 135978
rect 70854 135922 70922 135978
rect 70978 135922 71046 135978
rect 71102 135922 101878 135978
rect 101934 135922 102002 135978
rect 102058 135922 132114 135978
rect 132170 135922 132238 135978
rect 132294 135922 132362 135978
rect 132418 135922 132486 135978
rect 132542 135922 162834 135978
rect 162890 135922 162958 135978
rect 163014 135922 163082 135978
rect 163138 135922 163206 135978
rect 163262 135922 163878 135978
rect 163934 135922 164002 135978
rect 164058 135922 193554 135978
rect 193610 135922 193678 135978
rect 193734 135922 193802 135978
rect 193858 135922 193926 135978
rect 193982 135922 224274 135978
rect 224330 135922 224398 135978
rect 224454 135922 224522 135978
rect 224578 135922 224646 135978
rect 224702 135922 225878 135978
rect 225934 135922 226002 135978
rect 226058 135922 254994 135978
rect 255050 135922 255118 135978
rect 255174 135922 255242 135978
rect 255298 135922 255366 135978
rect 255422 135922 287878 135978
rect 287934 135922 288002 135978
rect 288058 135922 318598 135978
rect 318654 135922 318722 135978
rect 318778 135922 347154 135978
rect 347210 135922 347278 135978
rect 347334 135922 347402 135978
rect 347458 135922 347526 135978
rect 347582 135922 371878 135978
rect 371934 135922 372002 135978
rect 372058 135922 377874 135978
rect 377930 135922 377998 135978
rect 378054 135922 378122 135978
rect 378178 135922 378246 135978
rect 378302 135922 408594 135978
rect 408650 135922 408718 135978
rect 408774 135922 408842 135978
rect 408898 135922 408966 135978
rect 409022 135922 433878 135978
rect 433934 135922 434002 135978
rect 434058 135922 439314 135978
rect 439370 135922 439438 135978
rect 439494 135922 439562 135978
rect 439618 135922 439686 135978
rect 439742 135922 470034 135978
rect 470090 135922 470158 135978
rect 470214 135922 470282 135978
rect 470338 135922 470406 135978
rect 470462 135922 495878 135978
rect 495934 135922 496002 135978
rect 496058 135922 500754 135978
rect 500810 135922 500878 135978
rect 500934 135922 501002 135978
rect 501058 135922 501126 135978
rect 501182 135922 531474 135978
rect 531530 135922 531598 135978
rect 531654 135922 531722 135978
rect 531778 135922 531846 135978
rect 531902 135922 557878 135978
rect 557934 135922 558002 135978
rect 558058 135922 562194 135978
rect 562250 135922 562318 135978
rect 562374 135922 562442 135978
rect 562498 135922 562566 135978
rect 562622 135922 592914 135978
rect 592970 135922 593038 135978
rect 593094 135922 593162 135978
rect 593218 135922 593286 135978
rect 593342 135922 597456 135978
rect 597512 135922 597580 135978
rect 597636 135922 597704 135978
rect 597760 135922 597828 135978
rect 597884 135922 597980 135978
rect -1916 135826 597980 135922
rect 334444 133498 457060 133514
rect 334444 133442 334460 133498
rect 334516 133442 456988 133498
rect 457044 133442 457060 133498
rect 334444 133426 457060 133442
rect 138556 132958 263860 132974
rect 138556 132902 138572 132958
rect 138628 132902 263788 132958
rect 263844 132902 263860 132958
rect 138556 132886 263860 132902
rect 80428 132778 263972 132794
rect 80428 132722 80444 132778
rect 80500 132722 263900 132778
rect 263956 132722 263972 132778
rect 80428 132706 263972 132722
rect 20060 131338 263972 131354
rect 20060 131282 20076 131338
rect 20132 131282 263900 131338
rect 263956 131282 263972 131338
rect 20060 131266 263972 131282
rect 334444 131338 400724 131354
rect 334444 131282 334460 131338
rect 334516 131282 400652 131338
rect 400708 131282 400724 131338
rect 334444 131266 400724 131282
rect 18380 131158 264868 131174
rect 18380 131102 18396 131158
rect 18452 131102 264796 131158
rect 264852 131102 264868 131158
rect 18380 131086 264868 131102
rect 334444 131158 404084 131174
rect 334444 131102 334460 131158
rect 334516 131102 404012 131158
rect 404068 131102 404084 131158
rect 334444 131086 404084 131102
rect -1916 130350 597980 130446
rect -1916 130294 -860 130350
rect -804 130294 -736 130350
rect -680 130294 -612 130350
rect -556 130294 -488 130350
rect -432 130294 5514 130350
rect 5570 130294 5638 130350
rect 5694 130294 5762 130350
rect 5818 130294 5886 130350
rect 5942 130294 24518 130350
rect 24574 130294 24642 130350
rect 24698 130294 36234 130350
rect 36290 130294 36358 130350
rect 36414 130294 36482 130350
rect 36538 130294 36606 130350
rect 36662 130294 55238 130350
rect 55294 130294 55362 130350
rect 55418 130294 66954 130350
rect 67010 130294 67078 130350
rect 67134 130294 67202 130350
rect 67258 130294 67326 130350
rect 67382 130294 86518 130350
rect 86574 130294 86642 130350
rect 86698 130294 97674 130350
rect 97730 130294 97798 130350
rect 97854 130294 97922 130350
rect 97978 130294 98046 130350
rect 98102 130294 117238 130350
rect 117294 130294 117362 130350
rect 117418 130294 128394 130350
rect 128450 130294 128518 130350
rect 128574 130294 128642 130350
rect 128698 130294 128766 130350
rect 128822 130294 148518 130350
rect 148574 130294 148642 130350
rect 148698 130294 159114 130350
rect 159170 130294 159238 130350
rect 159294 130294 159362 130350
rect 159418 130294 159486 130350
rect 159542 130294 179238 130350
rect 179294 130294 179362 130350
rect 179418 130294 189834 130350
rect 189890 130294 189958 130350
rect 190014 130294 190082 130350
rect 190138 130294 190206 130350
rect 190262 130294 210518 130350
rect 210574 130294 210642 130350
rect 210698 130294 220554 130350
rect 220610 130294 220678 130350
rect 220734 130294 220802 130350
rect 220858 130294 220926 130350
rect 220982 130294 241238 130350
rect 241294 130294 241362 130350
rect 241418 130294 251274 130350
rect 251330 130294 251398 130350
rect 251454 130294 251522 130350
rect 251578 130294 251646 130350
rect 251702 130294 272518 130350
rect 272574 130294 272642 130350
rect 272698 130294 303238 130350
rect 303294 130294 303362 130350
rect 303418 130294 343434 130350
rect 343490 130294 343558 130350
rect 343614 130294 343682 130350
rect 343738 130294 343806 130350
rect 343862 130294 356518 130350
rect 356574 130294 356642 130350
rect 356698 130294 374154 130350
rect 374210 130294 374278 130350
rect 374334 130294 374402 130350
rect 374458 130294 374526 130350
rect 374582 130294 387238 130350
rect 387294 130294 387362 130350
rect 387418 130294 404874 130350
rect 404930 130294 404998 130350
rect 405054 130294 405122 130350
rect 405178 130294 405246 130350
rect 405302 130294 418518 130350
rect 418574 130294 418642 130350
rect 418698 130294 435594 130350
rect 435650 130294 435718 130350
rect 435774 130294 435842 130350
rect 435898 130294 435966 130350
rect 436022 130294 449238 130350
rect 449294 130294 449362 130350
rect 449418 130294 466314 130350
rect 466370 130294 466438 130350
rect 466494 130294 466562 130350
rect 466618 130294 466686 130350
rect 466742 130294 480518 130350
rect 480574 130294 480642 130350
rect 480698 130294 497034 130350
rect 497090 130294 497158 130350
rect 497214 130294 497282 130350
rect 497338 130294 497406 130350
rect 497462 130294 511238 130350
rect 511294 130294 511362 130350
rect 511418 130294 527754 130350
rect 527810 130294 527878 130350
rect 527934 130294 528002 130350
rect 528058 130294 528126 130350
rect 528182 130294 542518 130350
rect 542574 130294 542642 130350
rect 542698 130294 558474 130350
rect 558530 130294 558598 130350
rect 558654 130294 558722 130350
rect 558778 130294 558846 130350
rect 558902 130294 573238 130350
rect 573294 130294 573362 130350
rect 573418 130294 589194 130350
rect 589250 130294 589318 130350
rect 589374 130294 589442 130350
rect 589498 130294 589566 130350
rect 589622 130294 596496 130350
rect 596552 130294 596620 130350
rect 596676 130294 596744 130350
rect 596800 130294 596868 130350
rect 596924 130294 597980 130350
rect -1916 130226 597980 130294
rect -1916 130170 -860 130226
rect -804 130170 -736 130226
rect -680 130170 -612 130226
rect -556 130170 -488 130226
rect -432 130170 5514 130226
rect 5570 130170 5638 130226
rect 5694 130170 5762 130226
rect 5818 130170 5886 130226
rect 5942 130170 24518 130226
rect 24574 130170 24642 130226
rect 24698 130170 36234 130226
rect 36290 130170 36358 130226
rect 36414 130170 36482 130226
rect 36538 130170 36606 130226
rect 36662 130170 55238 130226
rect 55294 130170 55362 130226
rect 55418 130170 66954 130226
rect 67010 130170 67078 130226
rect 67134 130170 67202 130226
rect 67258 130170 67326 130226
rect 67382 130170 86518 130226
rect 86574 130170 86642 130226
rect 86698 130170 97674 130226
rect 97730 130170 97798 130226
rect 97854 130170 97922 130226
rect 97978 130170 98046 130226
rect 98102 130170 117238 130226
rect 117294 130170 117362 130226
rect 117418 130170 128394 130226
rect 128450 130170 128518 130226
rect 128574 130170 128642 130226
rect 128698 130170 128766 130226
rect 128822 130170 148518 130226
rect 148574 130170 148642 130226
rect 148698 130170 159114 130226
rect 159170 130170 159238 130226
rect 159294 130170 159362 130226
rect 159418 130170 159486 130226
rect 159542 130170 179238 130226
rect 179294 130170 179362 130226
rect 179418 130170 189834 130226
rect 189890 130170 189958 130226
rect 190014 130170 190082 130226
rect 190138 130170 190206 130226
rect 190262 130170 210518 130226
rect 210574 130170 210642 130226
rect 210698 130170 220554 130226
rect 220610 130170 220678 130226
rect 220734 130170 220802 130226
rect 220858 130170 220926 130226
rect 220982 130170 241238 130226
rect 241294 130170 241362 130226
rect 241418 130170 251274 130226
rect 251330 130170 251398 130226
rect 251454 130170 251522 130226
rect 251578 130170 251646 130226
rect 251702 130170 272518 130226
rect 272574 130170 272642 130226
rect 272698 130170 303238 130226
rect 303294 130170 303362 130226
rect 303418 130170 343434 130226
rect 343490 130170 343558 130226
rect 343614 130170 343682 130226
rect 343738 130170 343806 130226
rect 343862 130170 356518 130226
rect 356574 130170 356642 130226
rect 356698 130170 374154 130226
rect 374210 130170 374278 130226
rect 374334 130170 374402 130226
rect 374458 130170 374526 130226
rect 374582 130170 387238 130226
rect 387294 130170 387362 130226
rect 387418 130170 404874 130226
rect 404930 130170 404998 130226
rect 405054 130170 405122 130226
rect 405178 130170 405246 130226
rect 405302 130170 418518 130226
rect 418574 130170 418642 130226
rect 418698 130170 435594 130226
rect 435650 130170 435718 130226
rect 435774 130170 435842 130226
rect 435898 130170 435966 130226
rect 436022 130170 449238 130226
rect 449294 130170 449362 130226
rect 449418 130170 466314 130226
rect 466370 130170 466438 130226
rect 466494 130170 466562 130226
rect 466618 130170 466686 130226
rect 466742 130170 480518 130226
rect 480574 130170 480642 130226
rect 480698 130170 497034 130226
rect 497090 130170 497158 130226
rect 497214 130170 497282 130226
rect 497338 130170 497406 130226
rect 497462 130170 511238 130226
rect 511294 130170 511362 130226
rect 511418 130170 527754 130226
rect 527810 130170 527878 130226
rect 527934 130170 528002 130226
rect 528058 130170 528126 130226
rect 528182 130170 542518 130226
rect 542574 130170 542642 130226
rect 542698 130170 558474 130226
rect 558530 130170 558598 130226
rect 558654 130170 558722 130226
rect 558778 130170 558846 130226
rect 558902 130170 573238 130226
rect 573294 130170 573362 130226
rect 573418 130170 589194 130226
rect 589250 130170 589318 130226
rect 589374 130170 589442 130226
rect 589498 130170 589566 130226
rect 589622 130170 596496 130226
rect 596552 130170 596620 130226
rect 596676 130170 596744 130226
rect 596800 130170 596868 130226
rect 596924 130170 597980 130226
rect -1916 130102 597980 130170
rect -1916 130046 -860 130102
rect -804 130046 -736 130102
rect -680 130046 -612 130102
rect -556 130046 -488 130102
rect -432 130046 5514 130102
rect 5570 130046 5638 130102
rect 5694 130046 5762 130102
rect 5818 130046 5886 130102
rect 5942 130046 24518 130102
rect 24574 130046 24642 130102
rect 24698 130046 36234 130102
rect 36290 130046 36358 130102
rect 36414 130046 36482 130102
rect 36538 130046 36606 130102
rect 36662 130046 55238 130102
rect 55294 130046 55362 130102
rect 55418 130046 66954 130102
rect 67010 130046 67078 130102
rect 67134 130046 67202 130102
rect 67258 130046 67326 130102
rect 67382 130046 86518 130102
rect 86574 130046 86642 130102
rect 86698 130046 97674 130102
rect 97730 130046 97798 130102
rect 97854 130046 97922 130102
rect 97978 130046 98046 130102
rect 98102 130046 117238 130102
rect 117294 130046 117362 130102
rect 117418 130046 128394 130102
rect 128450 130046 128518 130102
rect 128574 130046 128642 130102
rect 128698 130046 128766 130102
rect 128822 130046 148518 130102
rect 148574 130046 148642 130102
rect 148698 130046 159114 130102
rect 159170 130046 159238 130102
rect 159294 130046 159362 130102
rect 159418 130046 159486 130102
rect 159542 130046 179238 130102
rect 179294 130046 179362 130102
rect 179418 130046 189834 130102
rect 189890 130046 189958 130102
rect 190014 130046 190082 130102
rect 190138 130046 190206 130102
rect 190262 130046 210518 130102
rect 210574 130046 210642 130102
rect 210698 130046 220554 130102
rect 220610 130046 220678 130102
rect 220734 130046 220802 130102
rect 220858 130046 220926 130102
rect 220982 130046 241238 130102
rect 241294 130046 241362 130102
rect 241418 130046 251274 130102
rect 251330 130046 251398 130102
rect 251454 130046 251522 130102
rect 251578 130046 251646 130102
rect 251702 130046 272518 130102
rect 272574 130046 272642 130102
rect 272698 130046 303238 130102
rect 303294 130046 303362 130102
rect 303418 130046 343434 130102
rect 343490 130046 343558 130102
rect 343614 130046 343682 130102
rect 343738 130046 343806 130102
rect 343862 130046 356518 130102
rect 356574 130046 356642 130102
rect 356698 130046 374154 130102
rect 374210 130046 374278 130102
rect 374334 130046 374402 130102
rect 374458 130046 374526 130102
rect 374582 130046 387238 130102
rect 387294 130046 387362 130102
rect 387418 130046 404874 130102
rect 404930 130046 404998 130102
rect 405054 130046 405122 130102
rect 405178 130046 405246 130102
rect 405302 130046 418518 130102
rect 418574 130046 418642 130102
rect 418698 130046 435594 130102
rect 435650 130046 435718 130102
rect 435774 130046 435842 130102
rect 435898 130046 435966 130102
rect 436022 130046 449238 130102
rect 449294 130046 449362 130102
rect 449418 130046 466314 130102
rect 466370 130046 466438 130102
rect 466494 130046 466562 130102
rect 466618 130046 466686 130102
rect 466742 130046 480518 130102
rect 480574 130046 480642 130102
rect 480698 130046 497034 130102
rect 497090 130046 497158 130102
rect 497214 130046 497282 130102
rect 497338 130046 497406 130102
rect 497462 130046 511238 130102
rect 511294 130046 511362 130102
rect 511418 130046 527754 130102
rect 527810 130046 527878 130102
rect 527934 130046 528002 130102
rect 528058 130046 528126 130102
rect 528182 130046 542518 130102
rect 542574 130046 542642 130102
rect 542698 130046 558474 130102
rect 558530 130046 558598 130102
rect 558654 130046 558722 130102
rect 558778 130046 558846 130102
rect 558902 130046 573238 130102
rect 573294 130046 573362 130102
rect 573418 130046 589194 130102
rect 589250 130046 589318 130102
rect 589374 130046 589442 130102
rect 589498 130046 589566 130102
rect 589622 130046 596496 130102
rect 596552 130046 596620 130102
rect 596676 130046 596744 130102
rect 596800 130046 596868 130102
rect 596924 130046 597980 130102
rect -1916 129978 597980 130046
rect -1916 129922 -860 129978
rect -804 129922 -736 129978
rect -680 129922 -612 129978
rect -556 129922 -488 129978
rect -432 129922 5514 129978
rect 5570 129922 5638 129978
rect 5694 129922 5762 129978
rect 5818 129922 5886 129978
rect 5942 129922 24518 129978
rect 24574 129922 24642 129978
rect 24698 129922 36234 129978
rect 36290 129922 36358 129978
rect 36414 129922 36482 129978
rect 36538 129922 36606 129978
rect 36662 129922 55238 129978
rect 55294 129922 55362 129978
rect 55418 129922 66954 129978
rect 67010 129922 67078 129978
rect 67134 129922 67202 129978
rect 67258 129922 67326 129978
rect 67382 129922 86518 129978
rect 86574 129922 86642 129978
rect 86698 129922 97674 129978
rect 97730 129922 97798 129978
rect 97854 129922 97922 129978
rect 97978 129922 98046 129978
rect 98102 129922 117238 129978
rect 117294 129922 117362 129978
rect 117418 129922 128394 129978
rect 128450 129922 128518 129978
rect 128574 129922 128642 129978
rect 128698 129922 128766 129978
rect 128822 129922 148518 129978
rect 148574 129922 148642 129978
rect 148698 129922 159114 129978
rect 159170 129922 159238 129978
rect 159294 129922 159362 129978
rect 159418 129922 159486 129978
rect 159542 129922 179238 129978
rect 179294 129922 179362 129978
rect 179418 129922 189834 129978
rect 189890 129922 189958 129978
rect 190014 129922 190082 129978
rect 190138 129922 190206 129978
rect 190262 129922 210518 129978
rect 210574 129922 210642 129978
rect 210698 129922 220554 129978
rect 220610 129922 220678 129978
rect 220734 129922 220802 129978
rect 220858 129922 220926 129978
rect 220982 129922 241238 129978
rect 241294 129922 241362 129978
rect 241418 129922 251274 129978
rect 251330 129922 251398 129978
rect 251454 129922 251522 129978
rect 251578 129922 251646 129978
rect 251702 129922 272518 129978
rect 272574 129922 272642 129978
rect 272698 129922 303238 129978
rect 303294 129922 303362 129978
rect 303418 129922 343434 129978
rect 343490 129922 343558 129978
rect 343614 129922 343682 129978
rect 343738 129922 343806 129978
rect 343862 129922 356518 129978
rect 356574 129922 356642 129978
rect 356698 129922 374154 129978
rect 374210 129922 374278 129978
rect 374334 129922 374402 129978
rect 374458 129922 374526 129978
rect 374582 129922 387238 129978
rect 387294 129922 387362 129978
rect 387418 129922 404874 129978
rect 404930 129922 404998 129978
rect 405054 129922 405122 129978
rect 405178 129922 405246 129978
rect 405302 129922 418518 129978
rect 418574 129922 418642 129978
rect 418698 129922 435594 129978
rect 435650 129922 435718 129978
rect 435774 129922 435842 129978
rect 435898 129922 435966 129978
rect 436022 129922 449238 129978
rect 449294 129922 449362 129978
rect 449418 129922 466314 129978
rect 466370 129922 466438 129978
rect 466494 129922 466562 129978
rect 466618 129922 466686 129978
rect 466742 129922 480518 129978
rect 480574 129922 480642 129978
rect 480698 129922 497034 129978
rect 497090 129922 497158 129978
rect 497214 129922 497282 129978
rect 497338 129922 497406 129978
rect 497462 129922 511238 129978
rect 511294 129922 511362 129978
rect 511418 129922 527754 129978
rect 527810 129922 527878 129978
rect 527934 129922 528002 129978
rect 528058 129922 528126 129978
rect 528182 129922 542518 129978
rect 542574 129922 542642 129978
rect 542698 129922 558474 129978
rect 558530 129922 558598 129978
rect 558654 129922 558722 129978
rect 558778 129922 558846 129978
rect 558902 129922 573238 129978
rect 573294 129922 573362 129978
rect 573418 129922 589194 129978
rect 589250 129922 589318 129978
rect 589374 129922 589442 129978
rect 589498 129922 589566 129978
rect 589622 129922 596496 129978
rect 596552 129922 596620 129978
rect 596676 129922 596744 129978
rect 596800 129922 596868 129978
rect 596924 129922 597980 129978
rect -1916 129826 597980 129922
rect 18268 128638 263860 128654
rect 18268 128582 18284 128638
rect 18340 128582 263788 128638
rect 263844 128582 263860 128638
rect 18268 128566 263860 128582
rect 149476 128458 201700 128474
rect 149476 128402 201628 128458
rect 201684 128402 201700 128458
rect 149476 128386 201700 128402
rect 352700 128458 473748 128474
rect 352700 128402 352716 128458
rect 352772 128402 411516 128458
rect 411572 128402 473676 128458
rect 473732 128402 473748 128458
rect 352700 128386 473748 128402
rect 149476 128114 149564 128386
rect 144044 128098 149564 128114
rect 144044 128042 144060 128098
rect 144116 128042 149564 128098
rect 144044 128026 149564 128042
rect 20060 127918 20204 127934
rect 20060 127862 20076 127918
rect 20132 127862 20204 127918
rect 20060 127846 20204 127862
rect 37756 127918 263972 127934
rect 37756 127862 37772 127918
rect 37828 127862 263900 127918
rect 263956 127862 263972 127918
rect 37756 127846 263972 127862
rect 476012 127918 478844 127934
rect 476012 127862 476028 127918
rect 476084 127862 478844 127918
rect 476012 127846 478844 127862
rect 20116 127754 20204 127846
rect 478756 127754 478844 127846
rect 20116 127738 141108 127754
rect 20116 127682 82684 127738
rect 82740 127682 141036 127738
rect 141092 127682 141108 127738
rect 20116 127666 141108 127682
rect 478756 127738 530868 127754
rect 478756 127682 530796 127738
rect 530852 127682 530868 127738
rect 478756 127666 530868 127682
rect 20620 127558 37844 127574
rect 20620 127502 20636 127558
rect 20692 127502 37772 127558
rect 37828 127502 37844 127558
rect 20620 127486 37844 127502
rect 334444 126838 384764 126854
rect 334444 126782 334460 126838
rect 334516 126782 384764 126838
rect 334444 126766 384764 126782
rect 384676 126674 384764 126766
rect 384676 126658 393332 126674
rect 384676 126602 393260 126658
rect 393316 126602 393332 126658
rect 384676 126586 393332 126602
rect 73820 126118 263860 126134
rect 73820 126062 73836 126118
rect 73892 126062 263788 126118
rect 263844 126062 263860 126118
rect 73820 126046 263860 126062
rect 82444 125938 138644 125954
rect 82444 125882 82460 125938
rect 82516 125882 138572 125938
rect 138628 125882 138644 125938
rect 82444 125866 138644 125882
rect 400636 125938 455492 125954
rect 400636 125882 400652 125938
rect 400708 125882 455492 125938
rect 400636 125866 455492 125882
rect 455404 125758 455492 125866
rect 455404 125702 455420 125758
rect 455476 125702 455492 125758
rect 455404 125686 455492 125702
rect 384676 125398 393444 125414
rect 384676 125342 393372 125398
rect 393428 125342 393444 125398
rect 384676 125326 393444 125342
rect 384676 125234 384764 125326
rect 161236 125218 263972 125234
rect 161236 125162 263900 125218
rect 263956 125162 263972 125218
rect 161236 125146 263972 125162
rect 334444 125218 384764 125234
rect 334444 125162 334460 125218
rect 334516 125162 384764 125218
rect 334444 125146 384764 125162
rect 161236 124334 161324 125146
rect 64188 124318 161324 124334
rect 64188 124262 64204 124318
rect 64260 124262 161324 124318
rect 64188 124246 161324 124262
rect 338476 124318 455324 124334
rect 338476 124262 338492 124318
rect 338548 124262 455324 124318
rect 338476 124246 455324 124262
rect 455236 123974 455324 124246
rect 455236 123958 455380 123974
rect 455236 123902 455308 123958
rect 455364 123902 455380 123958
rect 455236 123886 455380 123902
rect 345196 122518 411252 122534
rect 345196 122462 345212 122518
rect 345268 122462 411180 122518
rect 411236 122462 411252 122518
rect 345196 122446 411252 122462
rect 172996 121798 264084 121814
rect 172996 121742 264012 121798
rect 264068 121742 264084 121798
rect 172996 121726 264084 121742
rect 172996 121094 173084 121726
rect 166220 121006 173084 121094
rect 166220 120914 166308 121006
rect 64188 120898 166308 120914
rect 64188 120842 64204 120898
rect 64260 120842 166308 120898
rect 64188 120826 166308 120842
rect 351916 120898 455324 120914
rect 351916 120842 351932 120898
rect 351988 120842 455324 120898
rect 351916 120826 455324 120842
rect 455236 120554 455324 120826
rect 455236 120538 455380 120554
rect 455236 120482 455308 120538
rect 455364 120482 455380 120538
rect 455236 120466 455380 120482
rect -1916 118350 597980 118446
rect -1916 118294 -1820 118350
rect -1764 118294 -1696 118350
rect -1640 118294 -1572 118350
rect -1516 118294 -1448 118350
rect -1392 118294 9234 118350
rect 9290 118294 9358 118350
rect 9414 118294 9482 118350
rect 9538 118294 9606 118350
rect 9662 118294 39878 118350
rect 39934 118294 40002 118350
rect 40058 118294 70674 118350
rect 70730 118294 70798 118350
rect 70854 118294 70922 118350
rect 70978 118294 71046 118350
rect 71102 118294 101878 118350
rect 101934 118294 102002 118350
rect 102058 118294 132114 118350
rect 132170 118294 132238 118350
rect 132294 118294 132362 118350
rect 132418 118294 132486 118350
rect 132542 118294 162834 118350
rect 162890 118294 162958 118350
rect 163014 118294 163082 118350
rect 163138 118294 163206 118350
rect 163262 118294 163878 118350
rect 163934 118294 164002 118350
rect 164058 118294 193554 118350
rect 193610 118294 193678 118350
rect 193734 118294 193802 118350
rect 193858 118294 193926 118350
rect 193982 118294 224274 118350
rect 224330 118294 224398 118350
rect 224454 118294 224522 118350
rect 224578 118294 224646 118350
rect 224702 118294 225878 118350
rect 225934 118294 226002 118350
rect 226058 118294 254994 118350
rect 255050 118294 255118 118350
rect 255174 118294 255242 118350
rect 255298 118294 255366 118350
rect 255422 118294 287878 118350
rect 287934 118294 288002 118350
rect 288058 118294 318598 118350
rect 318654 118294 318722 118350
rect 318778 118294 347154 118350
rect 347210 118294 347278 118350
rect 347334 118294 347402 118350
rect 347458 118294 347526 118350
rect 347582 118294 371878 118350
rect 371934 118294 372002 118350
rect 372058 118294 377874 118350
rect 377930 118294 377998 118350
rect 378054 118294 378122 118350
rect 378178 118294 378246 118350
rect 378302 118294 408594 118350
rect 408650 118294 408718 118350
rect 408774 118294 408842 118350
rect 408898 118294 408966 118350
rect 409022 118294 433878 118350
rect 433934 118294 434002 118350
rect 434058 118294 439314 118350
rect 439370 118294 439438 118350
rect 439494 118294 439562 118350
rect 439618 118294 439686 118350
rect 439742 118294 470034 118350
rect 470090 118294 470158 118350
rect 470214 118294 470282 118350
rect 470338 118294 470406 118350
rect 470462 118294 495878 118350
rect 495934 118294 496002 118350
rect 496058 118294 500754 118350
rect 500810 118294 500878 118350
rect 500934 118294 501002 118350
rect 501058 118294 501126 118350
rect 501182 118294 531474 118350
rect 531530 118294 531598 118350
rect 531654 118294 531722 118350
rect 531778 118294 531846 118350
rect 531902 118294 557878 118350
rect 557934 118294 558002 118350
rect 558058 118294 562194 118350
rect 562250 118294 562318 118350
rect 562374 118294 562442 118350
rect 562498 118294 562566 118350
rect 562622 118294 592914 118350
rect 592970 118294 593038 118350
rect 593094 118294 593162 118350
rect 593218 118294 593286 118350
rect 593342 118294 597456 118350
rect 597512 118294 597580 118350
rect 597636 118294 597704 118350
rect 597760 118294 597828 118350
rect 597884 118294 597980 118350
rect -1916 118226 597980 118294
rect -1916 118170 -1820 118226
rect -1764 118170 -1696 118226
rect -1640 118170 -1572 118226
rect -1516 118170 -1448 118226
rect -1392 118170 9234 118226
rect 9290 118170 9358 118226
rect 9414 118170 9482 118226
rect 9538 118170 9606 118226
rect 9662 118170 39878 118226
rect 39934 118170 40002 118226
rect 40058 118170 70674 118226
rect 70730 118170 70798 118226
rect 70854 118170 70922 118226
rect 70978 118170 71046 118226
rect 71102 118170 101878 118226
rect 101934 118170 102002 118226
rect 102058 118170 132114 118226
rect 132170 118170 132238 118226
rect 132294 118170 132362 118226
rect 132418 118170 132486 118226
rect 132542 118170 162834 118226
rect 162890 118170 162958 118226
rect 163014 118170 163082 118226
rect 163138 118170 163206 118226
rect 163262 118170 163878 118226
rect 163934 118170 164002 118226
rect 164058 118170 193554 118226
rect 193610 118170 193678 118226
rect 193734 118170 193802 118226
rect 193858 118170 193926 118226
rect 193982 118170 224274 118226
rect 224330 118170 224398 118226
rect 224454 118170 224522 118226
rect 224578 118170 224646 118226
rect 224702 118170 225878 118226
rect 225934 118170 226002 118226
rect 226058 118170 254994 118226
rect 255050 118170 255118 118226
rect 255174 118170 255242 118226
rect 255298 118170 255366 118226
rect 255422 118170 287878 118226
rect 287934 118170 288002 118226
rect 288058 118170 318598 118226
rect 318654 118170 318722 118226
rect 318778 118170 347154 118226
rect 347210 118170 347278 118226
rect 347334 118170 347402 118226
rect 347458 118170 347526 118226
rect 347582 118170 371878 118226
rect 371934 118170 372002 118226
rect 372058 118170 377874 118226
rect 377930 118170 377998 118226
rect 378054 118170 378122 118226
rect 378178 118170 378246 118226
rect 378302 118170 408594 118226
rect 408650 118170 408718 118226
rect 408774 118170 408842 118226
rect 408898 118170 408966 118226
rect 409022 118170 433878 118226
rect 433934 118170 434002 118226
rect 434058 118170 439314 118226
rect 439370 118170 439438 118226
rect 439494 118170 439562 118226
rect 439618 118170 439686 118226
rect 439742 118170 470034 118226
rect 470090 118170 470158 118226
rect 470214 118170 470282 118226
rect 470338 118170 470406 118226
rect 470462 118170 495878 118226
rect 495934 118170 496002 118226
rect 496058 118170 500754 118226
rect 500810 118170 500878 118226
rect 500934 118170 501002 118226
rect 501058 118170 501126 118226
rect 501182 118170 531474 118226
rect 531530 118170 531598 118226
rect 531654 118170 531722 118226
rect 531778 118170 531846 118226
rect 531902 118170 557878 118226
rect 557934 118170 558002 118226
rect 558058 118170 562194 118226
rect 562250 118170 562318 118226
rect 562374 118170 562442 118226
rect 562498 118170 562566 118226
rect 562622 118170 592914 118226
rect 592970 118170 593038 118226
rect 593094 118170 593162 118226
rect 593218 118170 593286 118226
rect 593342 118170 597456 118226
rect 597512 118170 597580 118226
rect 597636 118170 597704 118226
rect 597760 118170 597828 118226
rect 597884 118170 597980 118226
rect -1916 118102 597980 118170
rect -1916 118046 -1820 118102
rect -1764 118046 -1696 118102
rect -1640 118046 -1572 118102
rect -1516 118046 -1448 118102
rect -1392 118046 9234 118102
rect 9290 118046 9358 118102
rect 9414 118046 9482 118102
rect 9538 118046 9606 118102
rect 9662 118046 39878 118102
rect 39934 118046 40002 118102
rect 40058 118046 70674 118102
rect 70730 118046 70798 118102
rect 70854 118046 70922 118102
rect 70978 118046 71046 118102
rect 71102 118046 101878 118102
rect 101934 118046 102002 118102
rect 102058 118046 132114 118102
rect 132170 118046 132238 118102
rect 132294 118046 132362 118102
rect 132418 118046 132486 118102
rect 132542 118046 162834 118102
rect 162890 118046 162958 118102
rect 163014 118046 163082 118102
rect 163138 118046 163206 118102
rect 163262 118046 163878 118102
rect 163934 118046 164002 118102
rect 164058 118046 193554 118102
rect 193610 118046 193678 118102
rect 193734 118046 193802 118102
rect 193858 118046 193926 118102
rect 193982 118046 224274 118102
rect 224330 118046 224398 118102
rect 224454 118046 224522 118102
rect 224578 118046 224646 118102
rect 224702 118046 225878 118102
rect 225934 118046 226002 118102
rect 226058 118046 254994 118102
rect 255050 118046 255118 118102
rect 255174 118046 255242 118102
rect 255298 118046 255366 118102
rect 255422 118046 287878 118102
rect 287934 118046 288002 118102
rect 288058 118046 318598 118102
rect 318654 118046 318722 118102
rect 318778 118046 347154 118102
rect 347210 118046 347278 118102
rect 347334 118046 347402 118102
rect 347458 118046 347526 118102
rect 347582 118046 371878 118102
rect 371934 118046 372002 118102
rect 372058 118046 377874 118102
rect 377930 118046 377998 118102
rect 378054 118046 378122 118102
rect 378178 118046 378246 118102
rect 378302 118046 408594 118102
rect 408650 118046 408718 118102
rect 408774 118046 408842 118102
rect 408898 118046 408966 118102
rect 409022 118046 433878 118102
rect 433934 118046 434002 118102
rect 434058 118046 439314 118102
rect 439370 118046 439438 118102
rect 439494 118046 439562 118102
rect 439618 118046 439686 118102
rect 439742 118046 470034 118102
rect 470090 118046 470158 118102
rect 470214 118046 470282 118102
rect 470338 118046 470406 118102
rect 470462 118046 495878 118102
rect 495934 118046 496002 118102
rect 496058 118046 500754 118102
rect 500810 118046 500878 118102
rect 500934 118046 501002 118102
rect 501058 118046 501126 118102
rect 501182 118046 531474 118102
rect 531530 118046 531598 118102
rect 531654 118046 531722 118102
rect 531778 118046 531846 118102
rect 531902 118046 557878 118102
rect 557934 118046 558002 118102
rect 558058 118046 562194 118102
rect 562250 118046 562318 118102
rect 562374 118046 562442 118102
rect 562498 118046 562566 118102
rect 562622 118046 592914 118102
rect 592970 118046 593038 118102
rect 593094 118046 593162 118102
rect 593218 118046 593286 118102
rect 593342 118046 597456 118102
rect 597512 118046 597580 118102
rect 597636 118046 597704 118102
rect 597760 118046 597828 118102
rect 597884 118046 597980 118102
rect -1916 117978 597980 118046
rect -1916 117922 -1820 117978
rect -1764 117922 -1696 117978
rect -1640 117922 -1572 117978
rect -1516 117922 -1448 117978
rect -1392 117922 9234 117978
rect 9290 117922 9358 117978
rect 9414 117922 9482 117978
rect 9538 117922 9606 117978
rect 9662 117922 39878 117978
rect 39934 117922 40002 117978
rect 40058 117922 70674 117978
rect 70730 117922 70798 117978
rect 70854 117922 70922 117978
rect 70978 117922 71046 117978
rect 71102 117922 101878 117978
rect 101934 117922 102002 117978
rect 102058 117922 132114 117978
rect 132170 117922 132238 117978
rect 132294 117922 132362 117978
rect 132418 117922 132486 117978
rect 132542 117922 162834 117978
rect 162890 117922 162958 117978
rect 163014 117922 163082 117978
rect 163138 117922 163206 117978
rect 163262 117922 163878 117978
rect 163934 117922 164002 117978
rect 164058 117922 193554 117978
rect 193610 117922 193678 117978
rect 193734 117922 193802 117978
rect 193858 117922 193926 117978
rect 193982 117922 224274 117978
rect 224330 117922 224398 117978
rect 224454 117922 224522 117978
rect 224578 117922 224646 117978
rect 224702 117922 225878 117978
rect 225934 117922 226002 117978
rect 226058 117922 254994 117978
rect 255050 117922 255118 117978
rect 255174 117922 255242 117978
rect 255298 117922 255366 117978
rect 255422 117922 287878 117978
rect 287934 117922 288002 117978
rect 288058 117922 318598 117978
rect 318654 117922 318722 117978
rect 318778 117922 347154 117978
rect 347210 117922 347278 117978
rect 347334 117922 347402 117978
rect 347458 117922 347526 117978
rect 347582 117922 371878 117978
rect 371934 117922 372002 117978
rect 372058 117922 377874 117978
rect 377930 117922 377998 117978
rect 378054 117922 378122 117978
rect 378178 117922 378246 117978
rect 378302 117922 408594 117978
rect 408650 117922 408718 117978
rect 408774 117922 408842 117978
rect 408898 117922 408966 117978
rect 409022 117922 433878 117978
rect 433934 117922 434002 117978
rect 434058 117922 439314 117978
rect 439370 117922 439438 117978
rect 439494 117922 439562 117978
rect 439618 117922 439686 117978
rect 439742 117922 470034 117978
rect 470090 117922 470158 117978
rect 470214 117922 470282 117978
rect 470338 117922 470406 117978
rect 470462 117922 495878 117978
rect 495934 117922 496002 117978
rect 496058 117922 500754 117978
rect 500810 117922 500878 117978
rect 500934 117922 501002 117978
rect 501058 117922 501126 117978
rect 501182 117922 531474 117978
rect 531530 117922 531598 117978
rect 531654 117922 531722 117978
rect 531778 117922 531846 117978
rect 531902 117922 557878 117978
rect 557934 117922 558002 117978
rect 558058 117922 562194 117978
rect 562250 117922 562318 117978
rect 562374 117922 562442 117978
rect 562498 117922 562566 117978
rect 562622 117922 592914 117978
rect 592970 117922 593038 117978
rect 593094 117922 593162 117978
rect 593218 117922 593286 117978
rect 593342 117922 597456 117978
rect 597512 117922 597580 117978
rect 597636 117922 597704 117978
rect 597760 117922 597828 117978
rect 597884 117922 597980 117978
rect -1916 117826 597980 117922
rect 64188 117478 260052 117494
rect 64188 117422 64204 117478
rect 64260 117422 259980 117478
rect 260036 117422 260052 117478
rect 64188 117406 260052 117422
rect -1916 112350 597980 112446
rect -1916 112294 -860 112350
rect -804 112294 -736 112350
rect -680 112294 -612 112350
rect -556 112294 -488 112350
rect -432 112294 5514 112350
rect 5570 112294 5638 112350
rect 5694 112294 5762 112350
rect 5818 112294 5886 112350
rect 5942 112294 24518 112350
rect 24574 112294 24642 112350
rect 24698 112294 36234 112350
rect 36290 112294 36358 112350
rect 36414 112294 36482 112350
rect 36538 112294 36606 112350
rect 36662 112294 55238 112350
rect 55294 112294 55362 112350
rect 55418 112294 66954 112350
rect 67010 112294 67078 112350
rect 67134 112294 67202 112350
rect 67258 112294 67326 112350
rect 67382 112294 86518 112350
rect 86574 112294 86642 112350
rect 86698 112294 97674 112350
rect 97730 112294 97798 112350
rect 97854 112294 97922 112350
rect 97978 112294 98046 112350
rect 98102 112294 117238 112350
rect 117294 112294 117362 112350
rect 117418 112294 128394 112350
rect 128450 112294 128518 112350
rect 128574 112294 128642 112350
rect 128698 112294 128766 112350
rect 128822 112294 148518 112350
rect 148574 112294 148642 112350
rect 148698 112294 159114 112350
rect 159170 112294 159238 112350
rect 159294 112294 159362 112350
rect 159418 112294 159486 112350
rect 159542 112294 179238 112350
rect 179294 112294 179362 112350
rect 179418 112294 189834 112350
rect 189890 112294 189958 112350
rect 190014 112294 190082 112350
rect 190138 112294 190206 112350
rect 190262 112294 210518 112350
rect 210574 112294 210642 112350
rect 210698 112294 220554 112350
rect 220610 112294 220678 112350
rect 220734 112294 220802 112350
rect 220858 112294 220926 112350
rect 220982 112294 241238 112350
rect 241294 112294 241362 112350
rect 241418 112294 251274 112350
rect 251330 112294 251398 112350
rect 251454 112294 251522 112350
rect 251578 112294 251646 112350
rect 251702 112294 272518 112350
rect 272574 112294 272642 112350
rect 272698 112294 303238 112350
rect 303294 112294 303362 112350
rect 303418 112294 343434 112350
rect 343490 112294 343558 112350
rect 343614 112294 343682 112350
rect 343738 112294 343806 112350
rect 343862 112294 356518 112350
rect 356574 112294 356642 112350
rect 356698 112294 374154 112350
rect 374210 112294 374278 112350
rect 374334 112294 374402 112350
rect 374458 112294 374526 112350
rect 374582 112294 387238 112350
rect 387294 112294 387362 112350
rect 387418 112294 404874 112350
rect 404930 112294 404998 112350
rect 405054 112294 405122 112350
rect 405178 112294 405246 112350
rect 405302 112294 418518 112350
rect 418574 112294 418642 112350
rect 418698 112294 435594 112350
rect 435650 112294 435718 112350
rect 435774 112294 435842 112350
rect 435898 112294 435966 112350
rect 436022 112294 449238 112350
rect 449294 112294 449362 112350
rect 449418 112294 466314 112350
rect 466370 112294 466438 112350
rect 466494 112294 466562 112350
rect 466618 112294 466686 112350
rect 466742 112294 480518 112350
rect 480574 112294 480642 112350
rect 480698 112294 497034 112350
rect 497090 112294 497158 112350
rect 497214 112294 497282 112350
rect 497338 112294 497406 112350
rect 497462 112294 511238 112350
rect 511294 112294 511362 112350
rect 511418 112294 527754 112350
rect 527810 112294 527878 112350
rect 527934 112294 528002 112350
rect 528058 112294 528126 112350
rect 528182 112294 542518 112350
rect 542574 112294 542642 112350
rect 542698 112294 558474 112350
rect 558530 112294 558598 112350
rect 558654 112294 558722 112350
rect 558778 112294 558846 112350
rect 558902 112294 573238 112350
rect 573294 112294 573362 112350
rect 573418 112294 589194 112350
rect 589250 112294 589318 112350
rect 589374 112294 589442 112350
rect 589498 112294 589566 112350
rect 589622 112294 596496 112350
rect 596552 112294 596620 112350
rect 596676 112294 596744 112350
rect 596800 112294 596868 112350
rect 596924 112294 597980 112350
rect -1916 112226 597980 112294
rect -1916 112170 -860 112226
rect -804 112170 -736 112226
rect -680 112170 -612 112226
rect -556 112170 -488 112226
rect -432 112170 5514 112226
rect 5570 112170 5638 112226
rect 5694 112170 5762 112226
rect 5818 112170 5886 112226
rect 5942 112170 24518 112226
rect 24574 112170 24642 112226
rect 24698 112170 36234 112226
rect 36290 112170 36358 112226
rect 36414 112170 36482 112226
rect 36538 112170 36606 112226
rect 36662 112170 55238 112226
rect 55294 112170 55362 112226
rect 55418 112170 66954 112226
rect 67010 112170 67078 112226
rect 67134 112170 67202 112226
rect 67258 112170 67326 112226
rect 67382 112170 86518 112226
rect 86574 112170 86642 112226
rect 86698 112170 97674 112226
rect 97730 112170 97798 112226
rect 97854 112170 97922 112226
rect 97978 112170 98046 112226
rect 98102 112170 117238 112226
rect 117294 112170 117362 112226
rect 117418 112170 128394 112226
rect 128450 112170 128518 112226
rect 128574 112170 128642 112226
rect 128698 112170 128766 112226
rect 128822 112170 148518 112226
rect 148574 112170 148642 112226
rect 148698 112170 159114 112226
rect 159170 112170 159238 112226
rect 159294 112170 159362 112226
rect 159418 112170 159486 112226
rect 159542 112170 179238 112226
rect 179294 112170 179362 112226
rect 179418 112170 189834 112226
rect 189890 112170 189958 112226
rect 190014 112170 190082 112226
rect 190138 112170 190206 112226
rect 190262 112170 210518 112226
rect 210574 112170 210642 112226
rect 210698 112170 220554 112226
rect 220610 112170 220678 112226
rect 220734 112170 220802 112226
rect 220858 112170 220926 112226
rect 220982 112170 241238 112226
rect 241294 112170 241362 112226
rect 241418 112170 251274 112226
rect 251330 112170 251398 112226
rect 251454 112170 251522 112226
rect 251578 112170 251646 112226
rect 251702 112170 272518 112226
rect 272574 112170 272642 112226
rect 272698 112170 303238 112226
rect 303294 112170 303362 112226
rect 303418 112170 343434 112226
rect 343490 112170 343558 112226
rect 343614 112170 343682 112226
rect 343738 112170 343806 112226
rect 343862 112170 356518 112226
rect 356574 112170 356642 112226
rect 356698 112170 374154 112226
rect 374210 112170 374278 112226
rect 374334 112170 374402 112226
rect 374458 112170 374526 112226
rect 374582 112170 387238 112226
rect 387294 112170 387362 112226
rect 387418 112170 404874 112226
rect 404930 112170 404998 112226
rect 405054 112170 405122 112226
rect 405178 112170 405246 112226
rect 405302 112170 418518 112226
rect 418574 112170 418642 112226
rect 418698 112170 435594 112226
rect 435650 112170 435718 112226
rect 435774 112170 435842 112226
rect 435898 112170 435966 112226
rect 436022 112170 449238 112226
rect 449294 112170 449362 112226
rect 449418 112170 466314 112226
rect 466370 112170 466438 112226
rect 466494 112170 466562 112226
rect 466618 112170 466686 112226
rect 466742 112170 480518 112226
rect 480574 112170 480642 112226
rect 480698 112170 497034 112226
rect 497090 112170 497158 112226
rect 497214 112170 497282 112226
rect 497338 112170 497406 112226
rect 497462 112170 511238 112226
rect 511294 112170 511362 112226
rect 511418 112170 527754 112226
rect 527810 112170 527878 112226
rect 527934 112170 528002 112226
rect 528058 112170 528126 112226
rect 528182 112170 542518 112226
rect 542574 112170 542642 112226
rect 542698 112170 558474 112226
rect 558530 112170 558598 112226
rect 558654 112170 558722 112226
rect 558778 112170 558846 112226
rect 558902 112170 573238 112226
rect 573294 112170 573362 112226
rect 573418 112170 589194 112226
rect 589250 112170 589318 112226
rect 589374 112170 589442 112226
rect 589498 112170 589566 112226
rect 589622 112170 596496 112226
rect 596552 112170 596620 112226
rect 596676 112170 596744 112226
rect 596800 112170 596868 112226
rect 596924 112170 597980 112226
rect -1916 112102 597980 112170
rect -1916 112046 -860 112102
rect -804 112046 -736 112102
rect -680 112046 -612 112102
rect -556 112046 -488 112102
rect -432 112046 5514 112102
rect 5570 112046 5638 112102
rect 5694 112046 5762 112102
rect 5818 112046 5886 112102
rect 5942 112046 24518 112102
rect 24574 112046 24642 112102
rect 24698 112046 36234 112102
rect 36290 112046 36358 112102
rect 36414 112046 36482 112102
rect 36538 112046 36606 112102
rect 36662 112046 55238 112102
rect 55294 112046 55362 112102
rect 55418 112046 66954 112102
rect 67010 112046 67078 112102
rect 67134 112046 67202 112102
rect 67258 112046 67326 112102
rect 67382 112046 86518 112102
rect 86574 112046 86642 112102
rect 86698 112046 97674 112102
rect 97730 112046 97798 112102
rect 97854 112046 97922 112102
rect 97978 112046 98046 112102
rect 98102 112046 117238 112102
rect 117294 112046 117362 112102
rect 117418 112046 128394 112102
rect 128450 112046 128518 112102
rect 128574 112046 128642 112102
rect 128698 112046 128766 112102
rect 128822 112046 148518 112102
rect 148574 112046 148642 112102
rect 148698 112046 159114 112102
rect 159170 112046 159238 112102
rect 159294 112046 159362 112102
rect 159418 112046 159486 112102
rect 159542 112046 179238 112102
rect 179294 112046 179362 112102
rect 179418 112046 189834 112102
rect 189890 112046 189958 112102
rect 190014 112046 190082 112102
rect 190138 112046 190206 112102
rect 190262 112046 210518 112102
rect 210574 112046 210642 112102
rect 210698 112046 220554 112102
rect 220610 112046 220678 112102
rect 220734 112046 220802 112102
rect 220858 112046 220926 112102
rect 220982 112046 241238 112102
rect 241294 112046 241362 112102
rect 241418 112046 251274 112102
rect 251330 112046 251398 112102
rect 251454 112046 251522 112102
rect 251578 112046 251646 112102
rect 251702 112046 272518 112102
rect 272574 112046 272642 112102
rect 272698 112046 303238 112102
rect 303294 112046 303362 112102
rect 303418 112046 343434 112102
rect 343490 112046 343558 112102
rect 343614 112046 343682 112102
rect 343738 112046 343806 112102
rect 343862 112046 356518 112102
rect 356574 112046 356642 112102
rect 356698 112046 374154 112102
rect 374210 112046 374278 112102
rect 374334 112046 374402 112102
rect 374458 112046 374526 112102
rect 374582 112046 387238 112102
rect 387294 112046 387362 112102
rect 387418 112046 404874 112102
rect 404930 112046 404998 112102
rect 405054 112046 405122 112102
rect 405178 112046 405246 112102
rect 405302 112046 418518 112102
rect 418574 112046 418642 112102
rect 418698 112046 435594 112102
rect 435650 112046 435718 112102
rect 435774 112046 435842 112102
rect 435898 112046 435966 112102
rect 436022 112046 449238 112102
rect 449294 112046 449362 112102
rect 449418 112046 466314 112102
rect 466370 112046 466438 112102
rect 466494 112046 466562 112102
rect 466618 112046 466686 112102
rect 466742 112046 480518 112102
rect 480574 112046 480642 112102
rect 480698 112046 497034 112102
rect 497090 112046 497158 112102
rect 497214 112046 497282 112102
rect 497338 112046 497406 112102
rect 497462 112046 511238 112102
rect 511294 112046 511362 112102
rect 511418 112046 527754 112102
rect 527810 112046 527878 112102
rect 527934 112046 528002 112102
rect 528058 112046 528126 112102
rect 528182 112046 542518 112102
rect 542574 112046 542642 112102
rect 542698 112046 558474 112102
rect 558530 112046 558598 112102
rect 558654 112046 558722 112102
rect 558778 112046 558846 112102
rect 558902 112046 573238 112102
rect 573294 112046 573362 112102
rect 573418 112046 589194 112102
rect 589250 112046 589318 112102
rect 589374 112046 589442 112102
rect 589498 112046 589566 112102
rect 589622 112046 596496 112102
rect 596552 112046 596620 112102
rect 596676 112046 596744 112102
rect 596800 112046 596868 112102
rect 596924 112046 597980 112102
rect -1916 111978 597980 112046
rect -1916 111922 -860 111978
rect -804 111922 -736 111978
rect -680 111922 -612 111978
rect -556 111922 -488 111978
rect -432 111922 5514 111978
rect 5570 111922 5638 111978
rect 5694 111922 5762 111978
rect 5818 111922 5886 111978
rect 5942 111922 24518 111978
rect 24574 111922 24642 111978
rect 24698 111922 36234 111978
rect 36290 111922 36358 111978
rect 36414 111922 36482 111978
rect 36538 111922 36606 111978
rect 36662 111922 55238 111978
rect 55294 111922 55362 111978
rect 55418 111922 66954 111978
rect 67010 111922 67078 111978
rect 67134 111922 67202 111978
rect 67258 111922 67326 111978
rect 67382 111922 86518 111978
rect 86574 111922 86642 111978
rect 86698 111922 97674 111978
rect 97730 111922 97798 111978
rect 97854 111922 97922 111978
rect 97978 111922 98046 111978
rect 98102 111922 117238 111978
rect 117294 111922 117362 111978
rect 117418 111922 128394 111978
rect 128450 111922 128518 111978
rect 128574 111922 128642 111978
rect 128698 111922 128766 111978
rect 128822 111922 148518 111978
rect 148574 111922 148642 111978
rect 148698 111922 159114 111978
rect 159170 111922 159238 111978
rect 159294 111922 159362 111978
rect 159418 111922 159486 111978
rect 159542 111922 179238 111978
rect 179294 111922 179362 111978
rect 179418 111922 189834 111978
rect 189890 111922 189958 111978
rect 190014 111922 190082 111978
rect 190138 111922 190206 111978
rect 190262 111922 210518 111978
rect 210574 111922 210642 111978
rect 210698 111922 220554 111978
rect 220610 111922 220678 111978
rect 220734 111922 220802 111978
rect 220858 111922 220926 111978
rect 220982 111922 241238 111978
rect 241294 111922 241362 111978
rect 241418 111922 251274 111978
rect 251330 111922 251398 111978
rect 251454 111922 251522 111978
rect 251578 111922 251646 111978
rect 251702 111922 272518 111978
rect 272574 111922 272642 111978
rect 272698 111922 303238 111978
rect 303294 111922 303362 111978
rect 303418 111922 343434 111978
rect 343490 111922 343558 111978
rect 343614 111922 343682 111978
rect 343738 111922 343806 111978
rect 343862 111922 356518 111978
rect 356574 111922 356642 111978
rect 356698 111922 374154 111978
rect 374210 111922 374278 111978
rect 374334 111922 374402 111978
rect 374458 111922 374526 111978
rect 374582 111922 387238 111978
rect 387294 111922 387362 111978
rect 387418 111922 404874 111978
rect 404930 111922 404998 111978
rect 405054 111922 405122 111978
rect 405178 111922 405246 111978
rect 405302 111922 418518 111978
rect 418574 111922 418642 111978
rect 418698 111922 435594 111978
rect 435650 111922 435718 111978
rect 435774 111922 435842 111978
rect 435898 111922 435966 111978
rect 436022 111922 449238 111978
rect 449294 111922 449362 111978
rect 449418 111922 466314 111978
rect 466370 111922 466438 111978
rect 466494 111922 466562 111978
rect 466618 111922 466686 111978
rect 466742 111922 480518 111978
rect 480574 111922 480642 111978
rect 480698 111922 497034 111978
rect 497090 111922 497158 111978
rect 497214 111922 497282 111978
rect 497338 111922 497406 111978
rect 497462 111922 511238 111978
rect 511294 111922 511362 111978
rect 511418 111922 527754 111978
rect 527810 111922 527878 111978
rect 527934 111922 528002 111978
rect 528058 111922 528126 111978
rect 528182 111922 542518 111978
rect 542574 111922 542642 111978
rect 542698 111922 558474 111978
rect 558530 111922 558598 111978
rect 558654 111922 558722 111978
rect 558778 111922 558846 111978
rect 558902 111922 573238 111978
rect 573294 111922 573362 111978
rect 573418 111922 589194 111978
rect 589250 111922 589318 111978
rect 589374 111922 589442 111978
rect 589498 111922 589566 111978
rect 589622 111922 596496 111978
rect 596552 111922 596620 111978
rect 596676 111922 596744 111978
rect 596800 111922 596868 111978
rect 596924 111922 597980 111978
rect -1916 111826 597980 111922
rect -1916 100350 597980 100446
rect -1916 100294 -1820 100350
rect -1764 100294 -1696 100350
rect -1640 100294 -1572 100350
rect -1516 100294 -1448 100350
rect -1392 100294 9234 100350
rect 9290 100294 9358 100350
rect 9414 100294 9482 100350
rect 9538 100294 9606 100350
rect 9662 100294 39954 100350
rect 40010 100294 40078 100350
rect 40134 100294 40202 100350
rect 40258 100294 40326 100350
rect 40382 100294 70674 100350
rect 70730 100294 70798 100350
rect 70854 100294 70922 100350
rect 70978 100294 71046 100350
rect 71102 100294 101394 100350
rect 101450 100294 101518 100350
rect 101574 100294 101642 100350
rect 101698 100294 101766 100350
rect 101822 100294 132114 100350
rect 132170 100294 132238 100350
rect 132294 100294 132362 100350
rect 132418 100294 132486 100350
rect 132542 100294 162834 100350
rect 162890 100294 162958 100350
rect 163014 100294 163082 100350
rect 163138 100294 163206 100350
rect 163262 100294 193554 100350
rect 193610 100294 193678 100350
rect 193734 100294 193802 100350
rect 193858 100294 193926 100350
rect 193982 100294 224274 100350
rect 224330 100294 224398 100350
rect 224454 100294 224522 100350
rect 224578 100294 224646 100350
rect 224702 100294 254994 100350
rect 255050 100294 255118 100350
rect 255174 100294 255242 100350
rect 255298 100294 255366 100350
rect 255422 100294 287878 100350
rect 287934 100294 288002 100350
rect 288058 100294 318598 100350
rect 318654 100294 318722 100350
rect 318778 100294 347154 100350
rect 347210 100294 347278 100350
rect 347334 100294 347402 100350
rect 347458 100294 347526 100350
rect 347582 100294 377874 100350
rect 377930 100294 377998 100350
rect 378054 100294 378122 100350
rect 378178 100294 378246 100350
rect 378302 100294 408594 100350
rect 408650 100294 408718 100350
rect 408774 100294 408842 100350
rect 408898 100294 408966 100350
rect 409022 100294 439314 100350
rect 439370 100294 439438 100350
rect 439494 100294 439562 100350
rect 439618 100294 439686 100350
rect 439742 100294 470034 100350
rect 470090 100294 470158 100350
rect 470214 100294 470282 100350
rect 470338 100294 470406 100350
rect 470462 100294 500754 100350
rect 500810 100294 500878 100350
rect 500934 100294 501002 100350
rect 501058 100294 501126 100350
rect 501182 100294 531474 100350
rect 531530 100294 531598 100350
rect 531654 100294 531722 100350
rect 531778 100294 531846 100350
rect 531902 100294 562194 100350
rect 562250 100294 562318 100350
rect 562374 100294 562442 100350
rect 562498 100294 562566 100350
rect 562622 100294 592914 100350
rect 592970 100294 593038 100350
rect 593094 100294 593162 100350
rect 593218 100294 593286 100350
rect 593342 100294 597456 100350
rect 597512 100294 597580 100350
rect 597636 100294 597704 100350
rect 597760 100294 597828 100350
rect 597884 100294 597980 100350
rect -1916 100226 597980 100294
rect -1916 100170 -1820 100226
rect -1764 100170 -1696 100226
rect -1640 100170 -1572 100226
rect -1516 100170 -1448 100226
rect -1392 100170 9234 100226
rect 9290 100170 9358 100226
rect 9414 100170 9482 100226
rect 9538 100170 9606 100226
rect 9662 100170 39954 100226
rect 40010 100170 40078 100226
rect 40134 100170 40202 100226
rect 40258 100170 40326 100226
rect 40382 100170 70674 100226
rect 70730 100170 70798 100226
rect 70854 100170 70922 100226
rect 70978 100170 71046 100226
rect 71102 100170 101394 100226
rect 101450 100170 101518 100226
rect 101574 100170 101642 100226
rect 101698 100170 101766 100226
rect 101822 100170 132114 100226
rect 132170 100170 132238 100226
rect 132294 100170 132362 100226
rect 132418 100170 132486 100226
rect 132542 100170 162834 100226
rect 162890 100170 162958 100226
rect 163014 100170 163082 100226
rect 163138 100170 163206 100226
rect 163262 100170 193554 100226
rect 193610 100170 193678 100226
rect 193734 100170 193802 100226
rect 193858 100170 193926 100226
rect 193982 100170 224274 100226
rect 224330 100170 224398 100226
rect 224454 100170 224522 100226
rect 224578 100170 224646 100226
rect 224702 100170 254994 100226
rect 255050 100170 255118 100226
rect 255174 100170 255242 100226
rect 255298 100170 255366 100226
rect 255422 100170 287878 100226
rect 287934 100170 288002 100226
rect 288058 100170 318598 100226
rect 318654 100170 318722 100226
rect 318778 100170 347154 100226
rect 347210 100170 347278 100226
rect 347334 100170 347402 100226
rect 347458 100170 347526 100226
rect 347582 100170 377874 100226
rect 377930 100170 377998 100226
rect 378054 100170 378122 100226
rect 378178 100170 378246 100226
rect 378302 100170 408594 100226
rect 408650 100170 408718 100226
rect 408774 100170 408842 100226
rect 408898 100170 408966 100226
rect 409022 100170 439314 100226
rect 439370 100170 439438 100226
rect 439494 100170 439562 100226
rect 439618 100170 439686 100226
rect 439742 100170 470034 100226
rect 470090 100170 470158 100226
rect 470214 100170 470282 100226
rect 470338 100170 470406 100226
rect 470462 100170 500754 100226
rect 500810 100170 500878 100226
rect 500934 100170 501002 100226
rect 501058 100170 501126 100226
rect 501182 100170 531474 100226
rect 531530 100170 531598 100226
rect 531654 100170 531722 100226
rect 531778 100170 531846 100226
rect 531902 100170 562194 100226
rect 562250 100170 562318 100226
rect 562374 100170 562442 100226
rect 562498 100170 562566 100226
rect 562622 100170 592914 100226
rect 592970 100170 593038 100226
rect 593094 100170 593162 100226
rect 593218 100170 593286 100226
rect 593342 100170 597456 100226
rect 597512 100170 597580 100226
rect 597636 100170 597704 100226
rect 597760 100170 597828 100226
rect 597884 100170 597980 100226
rect -1916 100102 597980 100170
rect -1916 100046 -1820 100102
rect -1764 100046 -1696 100102
rect -1640 100046 -1572 100102
rect -1516 100046 -1448 100102
rect -1392 100046 9234 100102
rect 9290 100046 9358 100102
rect 9414 100046 9482 100102
rect 9538 100046 9606 100102
rect 9662 100046 39954 100102
rect 40010 100046 40078 100102
rect 40134 100046 40202 100102
rect 40258 100046 40326 100102
rect 40382 100046 70674 100102
rect 70730 100046 70798 100102
rect 70854 100046 70922 100102
rect 70978 100046 71046 100102
rect 71102 100046 101394 100102
rect 101450 100046 101518 100102
rect 101574 100046 101642 100102
rect 101698 100046 101766 100102
rect 101822 100046 132114 100102
rect 132170 100046 132238 100102
rect 132294 100046 132362 100102
rect 132418 100046 132486 100102
rect 132542 100046 162834 100102
rect 162890 100046 162958 100102
rect 163014 100046 163082 100102
rect 163138 100046 163206 100102
rect 163262 100046 193554 100102
rect 193610 100046 193678 100102
rect 193734 100046 193802 100102
rect 193858 100046 193926 100102
rect 193982 100046 224274 100102
rect 224330 100046 224398 100102
rect 224454 100046 224522 100102
rect 224578 100046 224646 100102
rect 224702 100046 254994 100102
rect 255050 100046 255118 100102
rect 255174 100046 255242 100102
rect 255298 100046 255366 100102
rect 255422 100046 287878 100102
rect 287934 100046 288002 100102
rect 288058 100046 318598 100102
rect 318654 100046 318722 100102
rect 318778 100046 347154 100102
rect 347210 100046 347278 100102
rect 347334 100046 347402 100102
rect 347458 100046 347526 100102
rect 347582 100046 377874 100102
rect 377930 100046 377998 100102
rect 378054 100046 378122 100102
rect 378178 100046 378246 100102
rect 378302 100046 408594 100102
rect 408650 100046 408718 100102
rect 408774 100046 408842 100102
rect 408898 100046 408966 100102
rect 409022 100046 439314 100102
rect 439370 100046 439438 100102
rect 439494 100046 439562 100102
rect 439618 100046 439686 100102
rect 439742 100046 470034 100102
rect 470090 100046 470158 100102
rect 470214 100046 470282 100102
rect 470338 100046 470406 100102
rect 470462 100046 500754 100102
rect 500810 100046 500878 100102
rect 500934 100046 501002 100102
rect 501058 100046 501126 100102
rect 501182 100046 531474 100102
rect 531530 100046 531598 100102
rect 531654 100046 531722 100102
rect 531778 100046 531846 100102
rect 531902 100046 562194 100102
rect 562250 100046 562318 100102
rect 562374 100046 562442 100102
rect 562498 100046 562566 100102
rect 562622 100046 592914 100102
rect 592970 100046 593038 100102
rect 593094 100046 593162 100102
rect 593218 100046 593286 100102
rect 593342 100046 597456 100102
rect 597512 100046 597580 100102
rect 597636 100046 597704 100102
rect 597760 100046 597828 100102
rect 597884 100046 597980 100102
rect -1916 99978 597980 100046
rect -1916 99922 -1820 99978
rect -1764 99922 -1696 99978
rect -1640 99922 -1572 99978
rect -1516 99922 -1448 99978
rect -1392 99922 9234 99978
rect 9290 99922 9358 99978
rect 9414 99922 9482 99978
rect 9538 99922 9606 99978
rect 9662 99922 39954 99978
rect 40010 99922 40078 99978
rect 40134 99922 40202 99978
rect 40258 99922 40326 99978
rect 40382 99922 70674 99978
rect 70730 99922 70798 99978
rect 70854 99922 70922 99978
rect 70978 99922 71046 99978
rect 71102 99922 101394 99978
rect 101450 99922 101518 99978
rect 101574 99922 101642 99978
rect 101698 99922 101766 99978
rect 101822 99922 132114 99978
rect 132170 99922 132238 99978
rect 132294 99922 132362 99978
rect 132418 99922 132486 99978
rect 132542 99922 162834 99978
rect 162890 99922 162958 99978
rect 163014 99922 163082 99978
rect 163138 99922 163206 99978
rect 163262 99922 193554 99978
rect 193610 99922 193678 99978
rect 193734 99922 193802 99978
rect 193858 99922 193926 99978
rect 193982 99922 224274 99978
rect 224330 99922 224398 99978
rect 224454 99922 224522 99978
rect 224578 99922 224646 99978
rect 224702 99922 254994 99978
rect 255050 99922 255118 99978
rect 255174 99922 255242 99978
rect 255298 99922 255366 99978
rect 255422 99922 287878 99978
rect 287934 99922 288002 99978
rect 288058 99922 318598 99978
rect 318654 99922 318722 99978
rect 318778 99922 347154 99978
rect 347210 99922 347278 99978
rect 347334 99922 347402 99978
rect 347458 99922 347526 99978
rect 347582 99922 377874 99978
rect 377930 99922 377998 99978
rect 378054 99922 378122 99978
rect 378178 99922 378246 99978
rect 378302 99922 408594 99978
rect 408650 99922 408718 99978
rect 408774 99922 408842 99978
rect 408898 99922 408966 99978
rect 409022 99922 439314 99978
rect 439370 99922 439438 99978
rect 439494 99922 439562 99978
rect 439618 99922 439686 99978
rect 439742 99922 470034 99978
rect 470090 99922 470158 99978
rect 470214 99922 470282 99978
rect 470338 99922 470406 99978
rect 470462 99922 500754 99978
rect 500810 99922 500878 99978
rect 500934 99922 501002 99978
rect 501058 99922 501126 99978
rect 501182 99922 531474 99978
rect 531530 99922 531598 99978
rect 531654 99922 531722 99978
rect 531778 99922 531846 99978
rect 531902 99922 562194 99978
rect 562250 99922 562318 99978
rect 562374 99922 562442 99978
rect 562498 99922 562566 99978
rect 562622 99922 592914 99978
rect 592970 99922 593038 99978
rect 593094 99922 593162 99978
rect 593218 99922 593286 99978
rect 593342 99922 597456 99978
rect 597512 99922 597580 99978
rect 597636 99922 597704 99978
rect 597760 99922 597828 99978
rect 597884 99922 597980 99978
rect -1916 99826 597980 99922
rect -1916 94350 597980 94446
rect -1916 94294 -860 94350
rect -804 94294 -736 94350
rect -680 94294 -612 94350
rect -556 94294 -488 94350
rect -432 94294 5514 94350
rect 5570 94294 5638 94350
rect 5694 94294 5762 94350
rect 5818 94294 5886 94350
rect 5942 94294 36234 94350
rect 36290 94294 36358 94350
rect 36414 94294 36482 94350
rect 36538 94294 36606 94350
rect 36662 94294 66954 94350
rect 67010 94294 67078 94350
rect 67134 94294 67202 94350
rect 67258 94294 67326 94350
rect 67382 94294 97674 94350
rect 97730 94294 97798 94350
rect 97854 94294 97922 94350
rect 97978 94294 98046 94350
rect 98102 94294 128394 94350
rect 128450 94294 128518 94350
rect 128574 94294 128642 94350
rect 128698 94294 128766 94350
rect 128822 94294 159114 94350
rect 159170 94294 159238 94350
rect 159294 94294 159362 94350
rect 159418 94294 159486 94350
rect 159542 94294 189834 94350
rect 189890 94294 189958 94350
rect 190014 94294 190082 94350
rect 190138 94294 190206 94350
rect 190262 94294 220554 94350
rect 220610 94294 220678 94350
rect 220734 94294 220802 94350
rect 220858 94294 220926 94350
rect 220982 94294 251274 94350
rect 251330 94294 251398 94350
rect 251454 94294 251522 94350
rect 251578 94294 251646 94350
rect 251702 94294 272518 94350
rect 272574 94294 272642 94350
rect 272698 94294 303238 94350
rect 303294 94294 303362 94350
rect 303418 94294 343434 94350
rect 343490 94294 343558 94350
rect 343614 94294 343682 94350
rect 343738 94294 343806 94350
rect 343862 94294 374154 94350
rect 374210 94294 374278 94350
rect 374334 94294 374402 94350
rect 374458 94294 374526 94350
rect 374582 94294 404874 94350
rect 404930 94294 404998 94350
rect 405054 94294 405122 94350
rect 405178 94294 405246 94350
rect 405302 94294 435594 94350
rect 435650 94294 435718 94350
rect 435774 94294 435842 94350
rect 435898 94294 435966 94350
rect 436022 94294 466314 94350
rect 466370 94294 466438 94350
rect 466494 94294 466562 94350
rect 466618 94294 466686 94350
rect 466742 94294 497034 94350
rect 497090 94294 497158 94350
rect 497214 94294 497282 94350
rect 497338 94294 497406 94350
rect 497462 94294 527754 94350
rect 527810 94294 527878 94350
rect 527934 94294 528002 94350
rect 528058 94294 528126 94350
rect 528182 94294 558474 94350
rect 558530 94294 558598 94350
rect 558654 94294 558722 94350
rect 558778 94294 558846 94350
rect 558902 94294 589194 94350
rect 589250 94294 589318 94350
rect 589374 94294 589442 94350
rect 589498 94294 589566 94350
rect 589622 94294 596496 94350
rect 596552 94294 596620 94350
rect 596676 94294 596744 94350
rect 596800 94294 596868 94350
rect 596924 94294 597980 94350
rect -1916 94226 597980 94294
rect -1916 94170 -860 94226
rect -804 94170 -736 94226
rect -680 94170 -612 94226
rect -556 94170 -488 94226
rect -432 94170 5514 94226
rect 5570 94170 5638 94226
rect 5694 94170 5762 94226
rect 5818 94170 5886 94226
rect 5942 94170 36234 94226
rect 36290 94170 36358 94226
rect 36414 94170 36482 94226
rect 36538 94170 36606 94226
rect 36662 94170 66954 94226
rect 67010 94170 67078 94226
rect 67134 94170 67202 94226
rect 67258 94170 67326 94226
rect 67382 94170 97674 94226
rect 97730 94170 97798 94226
rect 97854 94170 97922 94226
rect 97978 94170 98046 94226
rect 98102 94170 128394 94226
rect 128450 94170 128518 94226
rect 128574 94170 128642 94226
rect 128698 94170 128766 94226
rect 128822 94170 159114 94226
rect 159170 94170 159238 94226
rect 159294 94170 159362 94226
rect 159418 94170 159486 94226
rect 159542 94170 189834 94226
rect 189890 94170 189958 94226
rect 190014 94170 190082 94226
rect 190138 94170 190206 94226
rect 190262 94170 220554 94226
rect 220610 94170 220678 94226
rect 220734 94170 220802 94226
rect 220858 94170 220926 94226
rect 220982 94170 251274 94226
rect 251330 94170 251398 94226
rect 251454 94170 251522 94226
rect 251578 94170 251646 94226
rect 251702 94170 272518 94226
rect 272574 94170 272642 94226
rect 272698 94170 303238 94226
rect 303294 94170 303362 94226
rect 303418 94170 343434 94226
rect 343490 94170 343558 94226
rect 343614 94170 343682 94226
rect 343738 94170 343806 94226
rect 343862 94170 374154 94226
rect 374210 94170 374278 94226
rect 374334 94170 374402 94226
rect 374458 94170 374526 94226
rect 374582 94170 404874 94226
rect 404930 94170 404998 94226
rect 405054 94170 405122 94226
rect 405178 94170 405246 94226
rect 405302 94170 435594 94226
rect 435650 94170 435718 94226
rect 435774 94170 435842 94226
rect 435898 94170 435966 94226
rect 436022 94170 466314 94226
rect 466370 94170 466438 94226
rect 466494 94170 466562 94226
rect 466618 94170 466686 94226
rect 466742 94170 497034 94226
rect 497090 94170 497158 94226
rect 497214 94170 497282 94226
rect 497338 94170 497406 94226
rect 497462 94170 527754 94226
rect 527810 94170 527878 94226
rect 527934 94170 528002 94226
rect 528058 94170 528126 94226
rect 528182 94170 558474 94226
rect 558530 94170 558598 94226
rect 558654 94170 558722 94226
rect 558778 94170 558846 94226
rect 558902 94170 589194 94226
rect 589250 94170 589318 94226
rect 589374 94170 589442 94226
rect 589498 94170 589566 94226
rect 589622 94170 596496 94226
rect 596552 94170 596620 94226
rect 596676 94170 596744 94226
rect 596800 94170 596868 94226
rect 596924 94170 597980 94226
rect -1916 94102 597980 94170
rect -1916 94046 -860 94102
rect -804 94046 -736 94102
rect -680 94046 -612 94102
rect -556 94046 -488 94102
rect -432 94046 5514 94102
rect 5570 94046 5638 94102
rect 5694 94046 5762 94102
rect 5818 94046 5886 94102
rect 5942 94046 36234 94102
rect 36290 94046 36358 94102
rect 36414 94046 36482 94102
rect 36538 94046 36606 94102
rect 36662 94046 66954 94102
rect 67010 94046 67078 94102
rect 67134 94046 67202 94102
rect 67258 94046 67326 94102
rect 67382 94046 97674 94102
rect 97730 94046 97798 94102
rect 97854 94046 97922 94102
rect 97978 94046 98046 94102
rect 98102 94046 128394 94102
rect 128450 94046 128518 94102
rect 128574 94046 128642 94102
rect 128698 94046 128766 94102
rect 128822 94046 159114 94102
rect 159170 94046 159238 94102
rect 159294 94046 159362 94102
rect 159418 94046 159486 94102
rect 159542 94046 189834 94102
rect 189890 94046 189958 94102
rect 190014 94046 190082 94102
rect 190138 94046 190206 94102
rect 190262 94046 220554 94102
rect 220610 94046 220678 94102
rect 220734 94046 220802 94102
rect 220858 94046 220926 94102
rect 220982 94046 251274 94102
rect 251330 94046 251398 94102
rect 251454 94046 251522 94102
rect 251578 94046 251646 94102
rect 251702 94046 272518 94102
rect 272574 94046 272642 94102
rect 272698 94046 303238 94102
rect 303294 94046 303362 94102
rect 303418 94046 343434 94102
rect 343490 94046 343558 94102
rect 343614 94046 343682 94102
rect 343738 94046 343806 94102
rect 343862 94046 374154 94102
rect 374210 94046 374278 94102
rect 374334 94046 374402 94102
rect 374458 94046 374526 94102
rect 374582 94046 404874 94102
rect 404930 94046 404998 94102
rect 405054 94046 405122 94102
rect 405178 94046 405246 94102
rect 405302 94046 435594 94102
rect 435650 94046 435718 94102
rect 435774 94046 435842 94102
rect 435898 94046 435966 94102
rect 436022 94046 466314 94102
rect 466370 94046 466438 94102
rect 466494 94046 466562 94102
rect 466618 94046 466686 94102
rect 466742 94046 497034 94102
rect 497090 94046 497158 94102
rect 497214 94046 497282 94102
rect 497338 94046 497406 94102
rect 497462 94046 527754 94102
rect 527810 94046 527878 94102
rect 527934 94046 528002 94102
rect 528058 94046 528126 94102
rect 528182 94046 558474 94102
rect 558530 94046 558598 94102
rect 558654 94046 558722 94102
rect 558778 94046 558846 94102
rect 558902 94046 589194 94102
rect 589250 94046 589318 94102
rect 589374 94046 589442 94102
rect 589498 94046 589566 94102
rect 589622 94046 596496 94102
rect 596552 94046 596620 94102
rect 596676 94046 596744 94102
rect 596800 94046 596868 94102
rect 596924 94046 597980 94102
rect -1916 93978 597980 94046
rect -1916 93922 -860 93978
rect -804 93922 -736 93978
rect -680 93922 -612 93978
rect -556 93922 -488 93978
rect -432 93922 5514 93978
rect 5570 93922 5638 93978
rect 5694 93922 5762 93978
rect 5818 93922 5886 93978
rect 5942 93922 36234 93978
rect 36290 93922 36358 93978
rect 36414 93922 36482 93978
rect 36538 93922 36606 93978
rect 36662 93922 66954 93978
rect 67010 93922 67078 93978
rect 67134 93922 67202 93978
rect 67258 93922 67326 93978
rect 67382 93922 97674 93978
rect 97730 93922 97798 93978
rect 97854 93922 97922 93978
rect 97978 93922 98046 93978
rect 98102 93922 128394 93978
rect 128450 93922 128518 93978
rect 128574 93922 128642 93978
rect 128698 93922 128766 93978
rect 128822 93922 159114 93978
rect 159170 93922 159238 93978
rect 159294 93922 159362 93978
rect 159418 93922 159486 93978
rect 159542 93922 189834 93978
rect 189890 93922 189958 93978
rect 190014 93922 190082 93978
rect 190138 93922 190206 93978
rect 190262 93922 220554 93978
rect 220610 93922 220678 93978
rect 220734 93922 220802 93978
rect 220858 93922 220926 93978
rect 220982 93922 251274 93978
rect 251330 93922 251398 93978
rect 251454 93922 251522 93978
rect 251578 93922 251646 93978
rect 251702 93922 272518 93978
rect 272574 93922 272642 93978
rect 272698 93922 303238 93978
rect 303294 93922 303362 93978
rect 303418 93922 343434 93978
rect 343490 93922 343558 93978
rect 343614 93922 343682 93978
rect 343738 93922 343806 93978
rect 343862 93922 374154 93978
rect 374210 93922 374278 93978
rect 374334 93922 374402 93978
rect 374458 93922 374526 93978
rect 374582 93922 404874 93978
rect 404930 93922 404998 93978
rect 405054 93922 405122 93978
rect 405178 93922 405246 93978
rect 405302 93922 435594 93978
rect 435650 93922 435718 93978
rect 435774 93922 435842 93978
rect 435898 93922 435966 93978
rect 436022 93922 466314 93978
rect 466370 93922 466438 93978
rect 466494 93922 466562 93978
rect 466618 93922 466686 93978
rect 466742 93922 497034 93978
rect 497090 93922 497158 93978
rect 497214 93922 497282 93978
rect 497338 93922 497406 93978
rect 497462 93922 527754 93978
rect 527810 93922 527878 93978
rect 527934 93922 528002 93978
rect 528058 93922 528126 93978
rect 528182 93922 558474 93978
rect 558530 93922 558598 93978
rect 558654 93922 558722 93978
rect 558778 93922 558846 93978
rect 558902 93922 589194 93978
rect 589250 93922 589318 93978
rect 589374 93922 589442 93978
rect 589498 93922 589566 93978
rect 589622 93922 596496 93978
rect 596552 93922 596620 93978
rect 596676 93922 596744 93978
rect 596800 93922 596868 93978
rect 596924 93922 597980 93978
rect -1916 93826 597980 93922
rect -1916 82350 597980 82446
rect -1916 82294 -1820 82350
rect -1764 82294 -1696 82350
rect -1640 82294 -1572 82350
rect -1516 82294 -1448 82350
rect -1392 82294 9234 82350
rect 9290 82294 9358 82350
rect 9414 82294 9482 82350
rect 9538 82294 9606 82350
rect 9662 82294 39954 82350
rect 40010 82294 40078 82350
rect 40134 82294 40202 82350
rect 40258 82294 40326 82350
rect 40382 82294 70674 82350
rect 70730 82294 70798 82350
rect 70854 82294 70922 82350
rect 70978 82294 71046 82350
rect 71102 82294 101394 82350
rect 101450 82294 101518 82350
rect 101574 82294 101642 82350
rect 101698 82294 101766 82350
rect 101822 82294 132114 82350
rect 132170 82294 132238 82350
rect 132294 82294 132362 82350
rect 132418 82294 132486 82350
rect 132542 82294 162834 82350
rect 162890 82294 162958 82350
rect 163014 82294 163082 82350
rect 163138 82294 163206 82350
rect 163262 82294 193554 82350
rect 193610 82294 193678 82350
rect 193734 82294 193802 82350
rect 193858 82294 193926 82350
rect 193982 82294 224274 82350
rect 224330 82294 224398 82350
rect 224454 82294 224522 82350
rect 224578 82294 224646 82350
rect 224702 82294 254994 82350
rect 255050 82294 255118 82350
rect 255174 82294 255242 82350
rect 255298 82294 255366 82350
rect 255422 82294 287878 82350
rect 287934 82294 288002 82350
rect 288058 82294 318598 82350
rect 318654 82294 318722 82350
rect 318778 82294 347154 82350
rect 347210 82294 347278 82350
rect 347334 82294 347402 82350
rect 347458 82294 347526 82350
rect 347582 82294 377874 82350
rect 377930 82294 377998 82350
rect 378054 82294 378122 82350
rect 378178 82294 378246 82350
rect 378302 82294 408594 82350
rect 408650 82294 408718 82350
rect 408774 82294 408842 82350
rect 408898 82294 408966 82350
rect 409022 82294 439314 82350
rect 439370 82294 439438 82350
rect 439494 82294 439562 82350
rect 439618 82294 439686 82350
rect 439742 82294 470034 82350
rect 470090 82294 470158 82350
rect 470214 82294 470282 82350
rect 470338 82294 470406 82350
rect 470462 82294 500754 82350
rect 500810 82294 500878 82350
rect 500934 82294 501002 82350
rect 501058 82294 501126 82350
rect 501182 82294 531474 82350
rect 531530 82294 531598 82350
rect 531654 82294 531722 82350
rect 531778 82294 531846 82350
rect 531902 82294 562194 82350
rect 562250 82294 562318 82350
rect 562374 82294 562442 82350
rect 562498 82294 562566 82350
rect 562622 82294 592914 82350
rect 592970 82294 593038 82350
rect 593094 82294 593162 82350
rect 593218 82294 593286 82350
rect 593342 82294 597456 82350
rect 597512 82294 597580 82350
rect 597636 82294 597704 82350
rect 597760 82294 597828 82350
rect 597884 82294 597980 82350
rect -1916 82226 597980 82294
rect -1916 82170 -1820 82226
rect -1764 82170 -1696 82226
rect -1640 82170 -1572 82226
rect -1516 82170 -1448 82226
rect -1392 82170 9234 82226
rect 9290 82170 9358 82226
rect 9414 82170 9482 82226
rect 9538 82170 9606 82226
rect 9662 82170 39954 82226
rect 40010 82170 40078 82226
rect 40134 82170 40202 82226
rect 40258 82170 40326 82226
rect 40382 82170 70674 82226
rect 70730 82170 70798 82226
rect 70854 82170 70922 82226
rect 70978 82170 71046 82226
rect 71102 82170 101394 82226
rect 101450 82170 101518 82226
rect 101574 82170 101642 82226
rect 101698 82170 101766 82226
rect 101822 82170 132114 82226
rect 132170 82170 132238 82226
rect 132294 82170 132362 82226
rect 132418 82170 132486 82226
rect 132542 82170 162834 82226
rect 162890 82170 162958 82226
rect 163014 82170 163082 82226
rect 163138 82170 163206 82226
rect 163262 82170 193554 82226
rect 193610 82170 193678 82226
rect 193734 82170 193802 82226
rect 193858 82170 193926 82226
rect 193982 82170 224274 82226
rect 224330 82170 224398 82226
rect 224454 82170 224522 82226
rect 224578 82170 224646 82226
rect 224702 82170 254994 82226
rect 255050 82170 255118 82226
rect 255174 82170 255242 82226
rect 255298 82170 255366 82226
rect 255422 82170 287878 82226
rect 287934 82170 288002 82226
rect 288058 82170 318598 82226
rect 318654 82170 318722 82226
rect 318778 82170 347154 82226
rect 347210 82170 347278 82226
rect 347334 82170 347402 82226
rect 347458 82170 347526 82226
rect 347582 82170 377874 82226
rect 377930 82170 377998 82226
rect 378054 82170 378122 82226
rect 378178 82170 378246 82226
rect 378302 82170 408594 82226
rect 408650 82170 408718 82226
rect 408774 82170 408842 82226
rect 408898 82170 408966 82226
rect 409022 82170 439314 82226
rect 439370 82170 439438 82226
rect 439494 82170 439562 82226
rect 439618 82170 439686 82226
rect 439742 82170 470034 82226
rect 470090 82170 470158 82226
rect 470214 82170 470282 82226
rect 470338 82170 470406 82226
rect 470462 82170 500754 82226
rect 500810 82170 500878 82226
rect 500934 82170 501002 82226
rect 501058 82170 501126 82226
rect 501182 82170 531474 82226
rect 531530 82170 531598 82226
rect 531654 82170 531722 82226
rect 531778 82170 531846 82226
rect 531902 82170 562194 82226
rect 562250 82170 562318 82226
rect 562374 82170 562442 82226
rect 562498 82170 562566 82226
rect 562622 82170 592914 82226
rect 592970 82170 593038 82226
rect 593094 82170 593162 82226
rect 593218 82170 593286 82226
rect 593342 82170 597456 82226
rect 597512 82170 597580 82226
rect 597636 82170 597704 82226
rect 597760 82170 597828 82226
rect 597884 82170 597980 82226
rect -1916 82102 597980 82170
rect -1916 82046 -1820 82102
rect -1764 82046 -1696 82102
rect -1640 82046 -1572 82102
rect -1516 82046 -1448 82102
rect -1392 82046 9234 82102
rect 9290 82046 9358 82102
rect 9414 82046 9482 82102
rect 9538 82046 9606 82102
rect 9662 82046 39954 82102
rect 40010 82046 40078 82102
rect 40134 82046 40202 82102
rect 40258 82046 40326 82102
rect 40382 82046 70674 82102
rect 70730 82046 70798 82102
rect 70854 82046 70922 82102
rect 70978 82046 71046 82102
rect 71102 82046 101394 82102
rect 101450 82046 101518 82102
rect 101574 82046 101642 82102
rect 101698 82046 101766 82102
rect 101822 82046 132114 82102
rect 132170 82046 132238 82102
rect 132294 82046 132362 82102
rect 132418 82046 132486 82102
rect 132542 82046 162834 82102
rect 162890 82046 162958 82102
rect 163014 82046 163082 82102
rect 163138 82046 163206 82102
rect 163262 82046 193554 82102
rect 193610 82046 193678 82102
rect 193734 82046 193802 82102
rect 193858 82046 193926 82102
rect 193982 82046 224274 82102
rect 224330 82046 224398 82102
rect 224454 82046 224522 82102
rect 224578 82046 224646 82102
rect 224702 82046 254994 82102
rect 255050 82046 255118 82102
rect 255174 82046 255242 82102
rect 255298 82046 255366 82102
rect 255422 82046 287878 82102
rect 287934 82046 288002 82102
rect 288058 82046 318598 82102
rect 318654 82046 318722 82102
rect 318778 82046 347154 82102
rect 347210 82046 347278 82102
rect 347334 82046 347402 82102
rect 347458 82046 347526 82102
rect 347582 82046 377874 82102
rect 377930 82046 377998 82102
rect 378054 82046 378122 82102
rect 378178 82046 378246 82102
rect 378302 82046 408594 82102
rect 408650 82046 408718 82102
rect 408774 82046 408842 82102
rect 408898 82046 408966 82102
rect 409022 82046 439314 82102
rect 439370 82046 439438 82102
rect 439494 82046 439562 82102
rect 439618 82046 439686 82102
rect 439742 82046 470034 82102
rect 470090 82046 470158 82102
rect 470214 82046 470282 82102
rect 470338 82046 470406 82102
rect 470462 82046 500754 82102
rect 500810 82046 500878 82102
rect 500934 82046 501002 82102
rect 501058 82046 501126 82102
rect 501182 82046 531474 82102
rect 531530 82046 531598 82102
rect 531654 82046 531722 82102
rect 531778 82046 531846 82102
rect 531902 82046 562194 82102
rect 562250 82046 562318 82102
rect 562374 82046 562442 82102
rect 562498 82046 562566 82102
rect 562622 82046 592914 82102
rect 592970 82046 593038 82102
rect 593094 82046 593162 82102
rect 593218 82046 593286 82102
rect 593342 82046 597456 82102
rect 597512 82046 597580 82102
rect 597636 82046 597704 82102
rect 597760 82046 597828 82102
rect 597884 82046 597980 82102
rect -1916 81978 597980 82046
rect -1916 81922 -1820 81978
rect -1764 81922 -1696 81978
rect -1640 81922 -1572 81978
rect -1516 81922 -1448 81978
rect -1392 81922 9234 81978
rect 9290 81922 9358 81978
rect 9414 81922 9482 81978
rect 9538 81922 9606 81978
rect 9662 81922 39954 81978
rect 40010 81922 40078 81978
rect 40134 81922 40202 81978
rect 40258 81922 40326 81978
rect 40382 81922 70674 81978
rect 70730 81922 70798 81978
rect 70854 81922 70922 81978
rect 70978 81922 71046 81978
rect 71102 81922 101394 81978
rect 101450 81922 101518 81978
rect 101574 81922 101642 81978
rect 101698 81922 101766 81978
rect 101822 81922 132114 81978
rect 132170 81922 132238 81978
rect 132294 81922 132362 81978
rect 132418 81922 132486 81978
rect 132542 81922 162834 81978
rect 162890 81922 162958 81978
rect 163014 81922 163082 81978
rect 163138 81922 163206 81978
rect 163262 81922 193554 81978
rect 193610 81922 193678 81978
rect 193734 81922 193802 81978
rect 193858 81922 193926 81978
rect 193982 81922 224274 81978
rect 224330 81922 224398 81978
rect 224454 81922 224522 81978
rect 224578 81922 224646 81978
rect 224702 81922 254994 81978
rect 255050 81922 255118 81978
rect 255174 81922 255242 81978
rect 255298 81922 255366 81978
rect 255422 81922 287878 81978
rect 287934 81922 288002 81978
rect 288058 81922 318598 81978
rect 318654 81922 318722 81978
rect 318778 81922 347154 81978
rect 347210 81922 347278 81978
rect 347334 81922 347402 81978
rect 347458 81922 347526 81978
rect 347582 81922 377874 81978
rect 377930 81922 377998 81978
rect 378054 81922 378122 81978
rect 378178 81922 378246 81978
rect 378302 81922 408594 81978
rect 408650 81922 408718 81978
rect 408774 81922 408842 81978
rect 408898 81922 408966 81978
rect 409022 81922 439314 81978
rect 439370 81922 439438 81978
rect 439494 81922 439562 81978
rect 439618 81922 439686 81978
rect 439742 81922 470034 81978
rect 470090 81922 470158 81978
rect 470214 81922 470282 81978
rect 470338 81922 470406 81978
rect 470462 81922 500754 81978
rect 500810 81922 500878 81978
rect 500934 81922 501002 81978
rect 501058 81922 501126 81978
rect 501182 81922 531474 81978
rect 531530 81922 531598 81978
rect 531654 81922 531722 81978
rect 531778 81922 531846 81978
rect 531902 81922 562194 81978
rect 562250 81922 562318 81978
rect 562374 81922 562442 81978
rect 562498 81922 562566 81978
rect 562622 81922 592914 81978
rect 592970 81922 593038 81978
rect 593094 81922 593162 81978
rect 593218 81922 593286 81978
rect 593342 81922 597456 81978
rect 597512 81922 597580 81978
rect 597636 81922 597704 81978
rect 597760 81922 597828 81978
rect 597884 81922 597980 81978
rect -1916 81826 597980 81922
rect -1916 76350 597980 76446
rect -1916 76294 -860 76350
rect -804 76294 -736 76350
rect -680 76294 -612 76350
rect -556 76294 -488 76350
rect -432 76294 5514 76350
rect 5570 76294 5638 76350
rect 5694 76294 5762 76350
rect 5818 76294 5886 76350
rect 5942 76294 36234 76350
rect 36290 76294 36358 76350
rect 36414 76294 36482 76350
rect 36538 76294 36606 76350
rect 36662 76294 66954 76350
rect 67010 76294 67078 76350
rect 67134 76294 67202 76350
rect 67258 76294 67326 76350
rect 67382 76294 97674 76350
rect 97730 76294 97798 76350
rect 97854 76294 97922 76350
rect 97978 76294 98046 76350
rect 98102 76294 128394 76350
rect 128450 76294 128518 76350
rect 128574 76294 128642 76350
rect 128698 76294 128766 76350
rect 128822 76294 159114 76350
rect 159170 76294 159238 76350
rect 159294 76294 159362 76350
rect 159418 76294 159486 76350
rect 159542 76294 189834 76350
rect 189890 76294 189958 76350
rect 190014 76294 190082 76350
rect 190138 76294 190206 76350
rect 190262 76294 220554 76350
rect 220610 76294 220678 76350
rect 220734 76294 220802 76350
rect 220858 76294 220926 76350
rect 220982 76294 251274 76350
rect 251330 76294 251398 76350
rect 251454 76294 251522 76350
rect 251578 76294 251646 76350
rect 251702 76294 272518 76350
rect 272574 76294 272642 76350
rect 272698 76294 303238 76350
rect 303294 76294 303362 76350
rect 303418 76294 343434 76350
rect 343490 76294 343558 76350
rect 343614 76294 343682 76350
rect 343738 76294 343806 76350
rect 343862 76294 374154 76350
rect 374210 76294 374278 76350
rect 374334 76294 374402 76350
rect 374458 76294 374526 76350
rect 374582 76294 404874 76350
rect 404930 76294 404998 76350
rect 405054 76294 405122 76350
rect 405178 76294 405246 76350
rect 405302 76294 435594 76350
rect 435650 76294 435718 76350
rect 435774 76294 435842 76350
rect 435898 76294 435966 76350
rect 436022 76294 466314 76350
rect 466370 76294 466438 76350
rect 466494 76294 466562 76350
rect 466618 76294 466686 76350
rect 466742 76294 497034 76350
rect 497090 76294 497158 76350
rect 497214 76294 497282 76350
rect 497338 76294 497406 76350
rect 497462 76294 527754 76350
rect 527810 76294 527878 76350
rect 527934 76294 528002 76350
rect 528058 76294 528126 76350
rect 528182 76294 558474 76350
rect 558530 76294 558598 76350
rect 558654 76294 558722 76350
rect 558778 76294 558846 76350
rect 558902 76294 589194 76350
rect 589250 76294 589318 76350
rect 589374 76294 589442 76350
rect 589498 76294 589566 76350
rect 589622 76294 596496 76350
rect 596552 76294 596620 76350
rect 596676 76294 596744 76350
rect 596800 76294 596868 76350
rect 596924 76294 597980 76350
rect -1916 76226 597980 76294
rect -1916 76170 -860 76226
rect -804 76170 -736 76226
rect -680 76170 -612 76226
rect -556 76170 -488 76226
rect -432 76170 5514 76226
rect 5570 76170 5638 76226
rect 5694 76170 5762 76226
rect 5818 76170 5886 76226
rect 5942 76170 36234 76226
rect 36290 76170 36358 76226
rect 36414 76170 36482 76226
rect 36538 76170 36606 76226
rect 36662 76170 66954 76226
rect 67010 76170 67078 76226
rect 67134 76170 67202 76226
rect 67258 76170 67326 76226
rect 67382 76170 97674 76226
rect 97730 76170 97798 76226
rect 97854 76170 97922 76226
rect 97978 76170 98046 76226
rect 98102 76170 128394 76226
rect 128450 76170 128518 76226
rect 128574 76170 128642 76226
rect 128698 76170 128766 76226
rect 128822 76170 159114 76226
rect 159170 76170 159238 76226
rect 159294 76170 159362 76226
rect 159418 76170 159486 76226
rect 159542 76170 189834 76226
rect 189890 76170 189958 76226
rect 190014 76170 190082 76226
rect 190138 76170 190206 76226
rect 190262 76170 220554 76226
rect 220610 76170 220678 76226
rect 220734 76170 220802 76226
rect 220858 76170 220926 76226
rect 220982 76170 251274 76226
rect 251330 76170 251398 76226
rect 251454 76170 251522 76226
rect 251578 76170 251646 76226
rect 251702 76170 272518 76226
rect 272574 76170 272642 76226
rect 272698 76170 303238 76226
rect 303294 76170 303362 76226
rect 303418 76170 343434 76226
rect 343490 76170 343558 76226
rect 343614 76170 343682 76226
rect 343738 76170 343806 76226
rect 343862 76170 374154 76226
rect 374210 76170 374278 76226
rect 374334 76170 374402 76226
rect 374458 76170 374526 76226
rect 374582 76170 404874 76226
rect 404930 76170 404998 76226
rect 405054 76170 405122 76226
rect 405178 76170 405246 76226
rect 405302 76170 435594 76226
rect 435650 76170 435718 76226
rect 435774 76170 435842 76226
rect 435898 76170 435966 76226
rect 436022 76170 466314 76226
rect 466370 76170 466438 76226
rect 466494 76170 466562 76226
rect 466618 76170 466686 76226
rect 466742 76170 497034 76226
rect 497090 76170 497158 76226
rect 497214 76170 497282 76226
rect 497338 76170 497406 76226
rect 497462 76170 527754 76226
rect 527810 76170 527878 76226
rect 527934 76170 528002 76226
rect 528058 76170 528126 76226
rect 528182 76170 558474 76226
rect 558530 76170 558598 76226
rect 558654 76170 558722 76226
rect 558778 76170 558846 76226
rect 558902 76170 589194 76226
rect 589250 76170 589318 76226
rect 589374 76170 589442 76226
rect 589498 76170 589566 76226
rect 589622 76170 596496 76226
rect 596552 76170 596620 76226
rect 596676 76170 596744 76226
rect 596800 76170 596868 76226
rect 596924 76170 597980 76226
rect -1916 76102 597980 76170
rect -1916 76046 -860 76102
rect -804 76046 -736 76102
rect -680 76046 -612 76102
rect -556 76046 -488 76102
rect -432 76046 5514 76102
rect 5570 76046 5638 76102
rect 5694 76046 5762 76102
rect 5818 76046 5886 76102
rect 5942 76046 36234 76102
rect 36290 76046 36358 76102
rect 36414 76046 36482 76102
rect 36538 76046 36606 76102
rect 36662 76046 66954 76102
rect 67010 76046 67078 76102
rect 67134 76046 67202 76102
rect 67258 76046 67326 76102
rect 67382 76046 97674 76102
rect 97730 76046 97798 76102
rect 97854 76046 97922 76102
rect 97978 76046 98046 76102
rect 98102 76046 128394 76102
rect 128450 76046 128518 76102
rect 128574 76046 128642 76102
rect 128698 76046 128766 76102
rect 128822 76046 159114 76102
rect 159170 76046 159238 76102
rect 159294 76046 159362 76102
rect 159418 76046 159486 76102
rect 159542 76046 189834 76102
rect 189890 76046 189958 76102
rect 190014 76046 190082 76102
rect 190138 76046 190206 76102
rect 190262 76046 220554 76102
rect 220610 76046 220678 76102
rect 220734 76046 220802 76102
rect 220858 76046 220926 76102
rect 220982 76046 251274 76102
rect 251330 76046 251398 76102
rect 251454 76046 251522 76102
rect 251578 76046 251646 76102
rect 251702 76046 272518 76102
rect 272574 76046 272642 76102
rect 272698 76046 303238 76102
rect 303294 76046 303362 76102
rect 303418 76046 343434 76102
rect 343490 76046 343558 76102
rect 343614 76046 343682 76102
rect 343738 76046 343806 76102
rect 343862 76046 374154 76102
rect 374210 76046 374278 76102
rect 374334 76046 374402 76102
rect 374458 76046 374526 76102
rect 374582 76046 404874 76102
rect 404930 76046 404998 76102
rect 405054 76046 405122 76102
rect 405178 76046 405246 76102
rect 405302 76046 435594 76102
rect 435650 76046 435718 76102
rect 435774 76046 435842 76102
rect 435898 76046 435966 76102
rect 436022 76046 466314 76102
rect 466370 76046 466438 76102
rect 466494 76046 466562 76102
rect 466618 76046 466686 76102
rect 466742 76046 497034 76102
rect 497090 76046 497158 76102
rect 497214 76046 497282 76102
rect 497338 76046 497406 76102
rect 497462 76046 527754 76102
rect 527810 76046 527878 76102
rect 527934 76046 528002 76102
rect 528058 76046 528126 76102
rect 528182 76046 558474 76102
rect 558530 76046 558598 76102
rect 558654 76046 558722 76102
rect 558778 76046 558846 76102
rect 558902 76046 589194 76102
rect 589250 76046 589318 76102
rect 589374 76046 589442 76102
rect 589498 76046 589566 76102
rect 589622 76046 596496 76102
rect 596552 76046 596620 76102
rect 596676 76046 596744 76102
rect 596800 76046 596868 76102
rect 596924 76046 597980 76102
rect -1916 75978 597980 76046
rect -1916 75922 -860 75978
rect -804 75922 -736 75978
rect -680 75922 -612 75978
rect -556 75922 -488 75978
rect -432 75922 5514 75978
rect 5570 75922 5638 75978
rect 5694 75922 5762 75978
rect 5818 75922 5886 75978
rect 5942 75922 36234 75978
rect 36290 75922 36358 75978
rect 36414 75922 36482 75978
rect 36538 75922 36606 75978
rect 36662 75922 66954 75978
rect 67010 75922 67078 75978
rect 67134 75922 67202 75978
rect 67258 75922 67326 75978
rect 67382 75922 97674 75978
rect 97730 75922 97798 75978
rect 97854 75922 97922 75978
rect 97978 75922 98046 75978
rect 98102 75922 128394 75978
rect 128450 75922 128518 75978
rect 128574 75922 128642 75978
rect 128698 75922 128766 75978
rect 128822 75922 159114 75978
rect 159170 75922 159238 75978
rect 159294 75922 159362 75978
rect 159418 75922 159486 75978
rect 159542 75922 189834 75978
rect 189890 75922 189958 75978
rect 190014 75922 190082 75978
rect 190138 75922 190206 75978
rect 190262 75922 220554 75978
rect 220610 75922 220678 75978
rect 220734 75922 220802 75978
rect 220858 75922 220926 75978
rect 220982 75922 251274 75978
rect 251330 75922 251398 75978
rect 251454 75922 251522 75978
rect 251578 75922 251646 75978
rect 251702 75922 272518 75978
rect 272574 75922 272642 75978
rect 272698 75922 303238 75978
rect 303294 75922 303362 75978
rect 303418 75922 343434 75978
rect 343490 75922 343558 75978
rect 343614 75922 343682 75978
rect 343738 75922 343806 75978
rect 343862 75922 374154 75978
rect 374210 75922 374278 75978
rect 374334 75922 374402 75978
rect 374458 75922 374526 75978
rect 374582 75922 404874 75978
rect 404930 75922 404998 75978
rect 405054 75922 405122 75978
rect 405178 75922 405246 75978
rect 405302 75922 435594 75978
rect 435650 75922 435718 75978
rect 435774 75922 435842 75978
rect 435898 75922 435966 75978
rect 436022 75922 466314 75978
rect 466370 75922 466438 75978
rect 466494 75922 466562 75978
rect 466618 75922 466686 75978
rect 466742 75922 497034 75978
rect 497090 75922 497158 75978
rect 497214 75922 497282 75978
rect 497338 75922 497406 75978
rect 497462 75922 527754 75978
rect 527810 75922 527878 75978
rect 527934 75922 528002 75978
rect 528058 75922 528126 75978
rect 528182 75922 558474 75978
rect 558530 75922 558598 75978
rect 558654 75922 558722 75978
rect 558778 75922 558846 75978
rect 558902 75922 589194 75978
rect 589250 75922 589318 75978
rect 589374 75922 589442 75978
rect 589498 75922 589566 75978
rect 589622 75922 596496 75978
rect 596552 75922 596620 75978
rect 596676 75922 596744 75978
rect 596800 75922 596868 75978
rect 596924 75922 597980 75978
rect -1916 75826 597980 75922
rect -1916 64350 597980 64446
rect -1916 64294 -1820 64350
rect -1764 64294 -1696 64350
rect -1640 64294 -1572 64350
rect -1516 64294 -1448 64350
rect -1392 64294 9234 64350
rect 9290 64294 9358 64350
rect 9414 64294 9482 64350
rect 9538 64294 9606 64350
rect 9662 64294 39878 64350
rect 39934 64294 40002 64350
rect 40058 64294 70674 64350
rect 70730 64294 70798 64350
rect 70854 64294 70922 64350
rect 70978 64294 71046 64350
rect 71102 64294 101878 64350
rect 101934 64294 102002 64350
rect 102058 64294 132114 64350
rect 132170 64294 132238 64350
rect 132294 64294 132362 64350
rect 132418 64294 132486 64350
rect 132542 64294 162834 64350
rect 162890 64294 162958 64350
rect 163014 64294 163082 64350
rect 163138 64294 163206 64350
rect 163262 64294 163878 64350
rect 163934 64294 164002 64350
rect 164058 64294 193554 64350
rect 193610 64294 193678 64350
rect 193734 64294 193802 64350
rect 193858 64294 193926 64350
rect 193982 64294 224274 64350
rect 224330 64294 224398 64350
rect 224454 64294 224522 64350
rect 224578 64294 224646 64350
rect 224702 64294 225878 64350
rect 225934 64294 226002 64350
rect 226058 64294 254994 64350
rect 255050 64294 255118 64350
rect 255174 64294 255242 64350
rect 255298 64294 255366 64350
rect 255422 64294 285714 64350
rect 285770 64294 285838 64350
rect 285894 64294 285962 64350
rect 286018 64294 286086 64350
rect 286142 64294 287878 64350
rect 287934 64294 288002 64350
rect 288058 64294 316434 64350
rect 316490 64294 316558 64350
rect 316614 64294 316682 64350
rect 316738 64294 316806 64350
rect 316862 64294 318598 64350
rect 318654 64294 318722 64350
rect 318778 64294 347154 64350
rect 347210 64294 347278 64350
rect 347334 64294 347402 64350
rect 347458 64294 347526 64350
rect 347582 64294 371878 64350
rect 371934 64294 372002 64350
rect 372058 64294 377874 64350
rect 377930 64294 377998 64350
rect 378054 64294 378122 64350
rect 378178 64294 378246 64350
rect 378302 64294 408594 64350
rect 408650 64294 408718 64350
rect 408774 64294 408842 64350
rect 408898 64294 408966 64350
rect 409022 64294 433878 64350
rect 433934 64294 434002 64350
rect 434058 64294 439314 64350
rect 439370 64294 439438 64350
rect 439494 64294 439562 64350
rect 439618 64294 439686 64350
rect 439742 64294 470034 64350
rect 470090 64294 470158 64350
rect 470214 64294 470282 64350
rect 470338 64294 470406 64350
rect 470462 64294 495878 64350
rect 495934 64294 496002 64350
rect 496058 64294 500754 64350
rect 500810 64294 500878 64350
rect 500934 64294 501002 64350
rect 501058 64294 501126 64350
rect 501182 64294 531474 64350
rect 531530 64294 531598 64350
rect 531654 64294 531722 64350
rect 531778 64294 531846 64350
rect 531902 64294 557878 64350
rect 557934 64294 558002 64350
rect 558058 64294 562194 64350
rect 562250 64294 562318 64350
rect 562374 64294 562442 64350
rect 562498 64294 562566 64350
rect 562622 64294 592914 64350
rect 592970 64294 593038 64350
rect 593094 64294 593162 64350
rect 593218 64294 593286 64350
rect 593342 64294 597456 64350
rect 597512 64294 597580 64350
rect 597636 64294 597704 64350
rect 597760 64294 597828 64350
rect 597884 64294 597980 64350
rect -1916 64226 597980 64294
rect -1916 64170 -1820 64226
rect -1764 64170 -1696 64226
rect -1640 64170 -1572 64226
rect -1516 64170 -1448 64226
rect -1392 64170 9234 64226
rect 9290 64170 9358 64226
rect 9414 64170 9482 64226
rect 9538 64170 9606 64226
rect 9662 64170 39878 64226
rect 39934 64170 40002 64226
rect 40058 64170 70674 64226
rect 70730 64170 70798 64226
rect 70854 64170 70922 64226
rect 70978 64170 71046 64226
rect 71102 64170 101878 64226
rect 101934 64170 102002 64226
rect 102058 64170 132114 64226
rect 132170 64170 132238 64226
rect 132294 64170 132362 64226
rect 132418 64170 132486 64226
rect 132542 64170 162834 64226
rect 162890 64170 162958 64226
rect 163014 64170 163082 64226
rect 163138 64170 163206 64226
rect 163262 64170 163878 64226
rect 163934 64170 164002 64226
rect 164058 64170 193554 64226
rect 193610 64170 193678 64226
rect 193734 64170 193802 64226
rect 193858 64170 193926 64226
rect 193982 64170 224274 64226
rect 224330 64170 224398 64226
rect 224454 64170 224522 64226
rect 224578 64170 224646 64226
rect 224702 64170 225878 64226
rect 225934 64170 226002 64226
rect 226058 64170 254994 64226
rect 255050 64170 255118 64226
rect 255174 64170 255242 64226
rect 255298 64170 255366 64226
rect 255422 64170 285714 64226
rect 285770 64170 285838 64226
rect 285894 64170 285962 64226
rect 286018 64170 286086 64226
rect 286142 64170 287878 64226
rect 287934 64170 288002 64226
rect 288058 64170 316434 64226
rect 316490 64170 316558 64226
rect 316614 64170 316682 64226
rect 316738 64170 316806 64226
rect 316862 64170 318598 64226
rect 318654 64170 318722 64226
rect 318778 64170 347154 64226
rect 347210 64170 347278 64226
rect 347334 64170 347402 64226
rect 347458 64170 347526 64226
rect 347582 64170 371878 64226
rect 371934 64170 372002 64226
rect 372058 64170 377874 64226
rect 377930 64170 377998 64226
rect 378054 64170 378122 64226
rect 378178 64170 378246 64226
rect 378302 64170 408594 64226
rect 408650 64170 408718 64226
rect 408774 64170 408842 64226
rect 408898 64170 408966 64226
rect 409022 64170 433878 64226
rect 433934 64170 434002 64226
rect 434058 64170 439314 64226
rect 439370 64170 439438 64226
rect 439494 64170 439562 64226
rect 439618 64170 439686 64226
rect 439742 64170 470034 64226
rect 470090 64170 470158 64226
rect 470214 64170 470282 64226
rect 470338 64170 470406 64226
rect 470462 64170 495878 64226
rect 495934 64170 496002 64226
rect 496058 64170 500754 64226
rect 500810 64170 500878 64226
rect 500934 64170 501002 64226
rect 501058 64170 501126 64226
rect 501182 64170 531474 64226
rect 531530 64170 531598 64226
rect 531654 64170 531722 64226
rect 531778 64170 531846 64226
rect 531902 64170 557878 64226
rect 557934 64170 558002 64226
rect 558058 64170 562194 64226
rect 562250 64170 562318 64226
rect 562374 64170 562442 64226
rect 562498 64170 562566 64226
rect 562622 64170 592914 64226
rect 592970 64170 593038 64226
rect 593094 64170 593162 64226
rect 593218 64170 593286 64226
rect 593342 64170 597456 64226
rect 597512 64170 597580 64226
rect 597636 64170 597704 64226
rect 597760 64170 597828 64226
rect 597884 64170 597980 64226
rect -1916 64102 597980 64170
rect -1916 64046 -1820 64102
rect -1764 64046 -1696 64102
rect -1640 64046 -1572 64102
rect -1516 64046 -1448 64102
rect -1392 64046 9234 64102
rect 9290 64046 9358 64102
rect 9414 64046 9482 64102
rect 9538 64046 9606 64102
rect 9662 64046 39878 64102
rect 39934 64046 40002 64102
rect 40058 64046 70674 64102
rect 70730 64046 70798 64102
rect 70854 64046 70922 64102
rect 70978 64046 71046 64102
rect 71102 64046 101878 64102
rect 101934 64046 102002 64102
rect 102058 64046 132114 64102
rect 132170 64046 132238 64102
rect 132294 64046 132362 64102
rect 132418 64046 132486 64102
rect 132542 64046 162834 64102
rect 162890 64046 162958 64102
rect 163014 64046 163082 64102
rect 163138 64046 163206 64102
rect 163262 64046 163878 64102
rect 163934 64046 164002 64102
rect 164058 64046 193554 64102
rect 193610 64046 193678 64102
rect 193734 64046 193802 64102
rect 193858 64046 193926 64102
rect 193982 64046 224274 64102
rect 224330 64046 224398 64102
rect 224454 64046 224522 64102
rect 224578 64046 224646 64102
rect 224702 64046 225878 64102
rect 225934 64046 226002 64102
rect 226058 64046 254994 64102
rect 255050 64046 255118 64102
rect 255174 64046 255242 64102
rect 255298 64046 255366 64102
rect 255422 64046 285714 64102
rect 285770 64046 285838 64102
rect 285894 64046 285962 64102
rect 286018 64046 286086 64102
rect 286142 64046 287878 64102
rect 287934 64046 288002 64102
rect 288058 64046 316434 64102
rect 316490 64046 316558 64102
rect 316614 64046 316682 64102
rect 316738 64046 316806 64102
rect 316862 64046 318598 64102
rect 318654 64046 318722 64102
rect 318778 64046 347154 64102
rect 347210 64046 347278 64102
rect 347334 64046 347402 64102
rect 347458 64046 347526 64102
rect 347582 64046 371878 64102
rect 371934 64046 372002 64102
rect 372058 64046 377874 64102
rect 377930 64046 377998 64102
rect 378054 64046 378122 64102
rect 378178 64046 378246 64102
rect 378302 64046 408594 64102
rect 408650 64046 408718 64102
rect 408774 64046 408842 64102
rect 408898 64046 408966 64102
rect 409022 64046 433878 64102
rect 433934 64046 434002 64102
rect 434058 64046 439314 64102
rect 439370 64046 439438 64102
rect 439494 64046 439562 64102
rect 439618 64046 439686 64102
rect 439742 64046 470034 64102
rect 470090 64046 470158 64102
rect 470214 64046 470282 64102
rect 470338 64046 470406 64102
rect 470462 64046 495878 64102
rect 495934 64046 496002 64102
rect 496058 64046 500754 64102
rect 500810 64046 500878 64102
rect 500934 64046 501002 64102
rect 501058 64046 501126 64102
rect 501182 64046 531474 64102
rect 531530 64046 531598 64102
rect 531654 64046 531722 64102
rect 531778 64046 531846 64102
rect 531902 64046 557878 64102
rect 557934 64046 558002 64102
rect 558058 64046 562194 64102
rect 562250 64046 562318 64102
rect 562374 64046 562442 64102
rect 562498 64046 562566 64102
rect 562622 64046 592914 64102
rect 592970 64046 593038 64102
rect 593094 64046 593162 64102
rect 593218 64046 593286 64102
rect 593342 64046 597456 64102
rect 597512 64046 597580 64102
rect 597636 64046 597704 64102
rect 597760 64046 597828 64102
rect 597884 64046 597980 64102
rect -1916 63978 597980 64046
rect -1916 63922 -1820 63978
rect -1764 63922 -1696 63978
rect -1640 63922 -1572 63978
rect -1516 63922 -1448 63978
rect -1392 63922 9234 63978
rect 9290 63922 9358 63978
rect 9414 63922 9482 63978
rect 9538 63922 9606 63978
rect 9662 63922 39878 63978
rect 39934 63922 40002 63978
rect 40058 63922 70674 63978
rect 70730 63922 70798 63978
rect 70854 63922 70922 63978
rect 70978 63922 71046 63978
rect 71102 63922 101878 63978
rect 101934 63922 102002 63978
rect 102058 63922 132114 63978
rect 132170 63922 132238 63978
rect 132294 63922 132362 63978
rect 132418 63922 132486 63978
rect 132542 63922 162834 63978
rect 162890 63922 162958 63978
rect 163014 63922 163082 63978
rect 163138 63922 163206 63978
rect 163262 63922 163878 63978
rect 163934 63922 164002 63978
rect 164058 63922 193554 63978
rect 193610 63922 193678 63978
rect 193734 63922 193802 63978
rect 193858 63922 193926 63978
rect 193982 63922 224274 63978
rect 224330 63922 224398 63978
rect 224454 63922 224522 63978
rect 224578 63922 224646 63978
rect 224702 63922 225878 63978
rect 225934 63922 226002 63978
rect 226058 63922 254994 63978
rect 255050 63922 255118 63978
rect 255174 63922 255242 63978
rect 255298 63922 255366 63978
rect 255422 63922 285714 63978
rect 285770 63922 285838 63978
rect 285894 63922 285962 63978
rect 286018 63922 286086 63978
rect 286142 63922 287878 63978
rect 287934 63922 288002 63978
rect 288058 63922 316434 63978
rect 316490 63922 316558 63978
rect 316614 63922 316682 63978
rect 316738 63922 316806 63978
rect 316862 63922 318598 63978
rect 318654 63922 318722 63978
rect 318778 63922 347154 63978
rect 347210 63922 347278 63978
rect 347334 63922 347402 63978
rect 347458 63922 347526 63978
rect 347582 63922 371878 63978
rect 371934 63922 372002 63978
rect 372058 63922 377874 63978
rect 377930 63922 377998 63978
rect 378054 63922 378122 63978
rect 378178 63922 378246 63978
rect 378302 63922 408594 63978
rect 408650 63922 408718 63978
rect 408774 63922 408842 63978
rect 408898 63922 408966 63978
rect 409022 63922 433878 63978
rect 433934 63922 434002 63978
rect 434058 63922 439314 63978
rect 439370 63922 439438 63978
rect 439494 63922 439562 63978
rect 439618 63922 439686 63978
rect 439742 63922 470034 63978
rect 470090 63922 470158 63978
rect 470214 63922 470282 63978
rect 470338 63922 470406 63978
rect 470462 63922 495878 63978
rect 495934 63922 496002 63978
rect 496058 63922 500754 63978
rect 500810 63922 500878 63978
rect 500934 63922 501002 63978
rect 501058 63922 501126 63978
rect 501182 63922 531474 63978
rect 531530 63922 531598 63978
rect 531654 63922 531722 63978
rect 531778 63922 531846 63978
rect 531902 63922 557878 63978
rect 557934 63922 558002 63978
rect 558058 63922 562194 63978
rect 562250 63922 562318 63978
rect 562374 63922 562442 63978
rect 562498 63922 562566 63978
rect 562622 63922 592914 63978
rect 592970 63922 593038 63978
rect 593094 63922 593162 63978
rect 593218 63922 593286 63978
rect 593342 63922 597456 63978
rect 597512 63922 597580 63978
rect 597636 63922 597704 63978
rect 597760 63922 597828 63978
rect 597884 63922 597980 63978
rect -1916 63826 597980 63922
rect -1916 58350 597980 58446
rect -1916 58294 -860 58350
rect -804 58294 -736 58350
rect -680 58294 -612 58350
rect -556 58294 -488 58350
rect -432 58294 5514 58350
rect 5570 58294 5638 58350
rect 5694 58294 5762 58350
rect 5818 58294 5886 58350
rect 5942 58294 24518 58350
rect 24574 58294 24642 58350
rect 24698 58294 36234 58350
rect 36290 58294 36358 58350
rect 36414 58294 36482 58350
rect 36538 58294 36606 58350
rect 36662 58294 55238 58350
rect 55294 58294 55362 58350
rect 55418 58294 66954 58350
rect 67010 58294 67078 58350
rect 67134 58294 67202 58350
rect 67258 58294 67326 58350
rect 67382 58294 86518 58350
rect 86574 58294 86642 58350
rect 86698 58294 97674 58350
rect 97730 58294 97798 58350
rect 97854 58294 97922 58350
rect 97978 58294 98046 58350
rect 98102 58294 117238 58350
rect 117294 58294 117362 58350
rect 117418 58294 128394 58350
rect 128450 58294 128518 58350
rect 128574 58294 128642 58350
rect 128698 58294 128766 58350
rect 128822 58294 148518 58350
rect 148574 58294 148642 58350
rect 148698 58294 159114 58350
rect 159170 58294 159238 58350
rect 159294 58294 159362 58350
rect 159418 58294 159486 58350
rect 159542 58294 179238 58350
rect 179294 58294 179362 58350
rect 179418 58294 189834 58350
rect 189890 58294 189958 58350
rect 190014 58294 190082 58350
rect 190138 58294 190206 58350
rect 190262 58294 210518 58350
rect 210574 58294 210642 58350
rect 210698 58294 220554 58350
rect 220610 58294 220678 58350
rect 220734 58294 220802 58350
rect 220858 58294 220926 58350
rect 220982 58294 241238 58350
rect 241294 58294 241362 58350
rect 241418 58294 251274 58350
rect 251330 58294 251398 58350
rect 251454 58294 251522 58350
rect 251578 58294 251646 58350
rect 251702 58294 272518 58350
rect 272574 58294 272642 58350
rect 272698 58294 281994 58350
rect 282050 58294 282118 58350
rect 282174 58294 282242 58350
rect 282298 58294 282366 58350
rect 282422 58294 303238 58350
rect 303294 58294 303362 58350
rect 303418 58294 312714 58350
rect 312770 58294 312838 58350
rect 312894 58294 312962 58350
rect 313018 58294 313086 58350
rect 313142 58294 343434 58350
rect 343490 58294 343558 58350
rect 343614 58294 343682 58350
rect 343738 58294 343806 58350
rect 343862 58294 356518 58350
rect 356574 58294 356642 58350
rect 356698 58294 374154 58350
rect 374210 58294 374278 58350
rect 374334 58294 374402 58350
rect 374458 58294 374526 58350
rect 374582 58294 387238 58350
rect 387294 58294 387362 58350
rect 387418 58294 404874 58350
rect 404930 58294 404998 58350
rect 405054 58294 405122 58350
rect 405178 58294 405246 58350
rect 405302 58294 418518 58350
rect 418574 58294 418642 58350
rect 418698 58294 435594 58350
rect 435650 58294 435718 58350
rect 435774 58294 435842 58350
rect 435898 58294 435966 58350
rect 436022 58294 449238 58350
rect 449294 58294 449362 58350
rect 449418 58294 466314 58350
rect 466370 58294 466438 58350
rect 466494 58294 466562 58350
rect 466618 58294 466686 58350
rect 466742 58294 480518 58350
rect 480574 58294 480642 58350
rect 480698 58294 497034 58350
rect 497090 58294 497158 58350
rect 497214 58294 497282 58350
rect 497338 58294 497406 58350
rect 497462 58294 511238 58350
rect 511294 58294 511362 58350
rect 511418 58294 527754 58350
rect 527810 58294 527878 58350
rect 527934 58294 528002 58350
rect 528058 58294 528126 58350
rect 528182 58294 542518 58350
rect 542574 58294 542642 58350
rect 542698 58294 558474 58350
rect 558530 58294 558598 58350
rect 558654 58294 558722 58350
rect 558778 58294 558846 58350
rect 558902 58294 573238 58350
rect 573294 58294 573362 58350
rect 573418 58294 589194 58350
rect 589250 58294 589318 58350
rect 589374 58294 589442 58350
rect 589498 58294 589566 58350
rect 589622 58294 596496 58350
rect 596552 58294 596620 58350
rect 596676 58294 596744 58350
rect 596800 58294 596868 58350
rect 596924 58294 597980 58350
rect -1916 58226 597980 58294
rect -1916 58170 -860 58226
rect -804 58170 -736 58226
rect -680 58170 -612 58226
rect -556 58170 -488 58226
rect -432 58170 5514 58226
rect 5570 58170 5638 58226
rect 5694 58170 5762 58226
rect 5818 58170 5886 58226
rect 5942 58170 24518 58226
rect 24574 58170 24642 58226
rect 24698 58170 36234 58226
rect 36290 58170 36358 58226
rect 36414 58170 36482 58226
rect 36538 58170 36606 58226
rect 36662 58170 55238 58226
rect 55294 58170 55362 58226
rect 55418 58170 66954 58226
rect 67010 58170 67078 58226
rect 67134 58170 67202 58226
rect 67258 58170 67326 58226
rect 67382 58170 86518 58226
rect 86574 58170 86642 58226
rect 86698 58170 97674 58226
rect 97730 58170 97798 58226
rect 97854 58170 97922 58226
rect 97978 58170 98046 58226
rect 98102 58170 117238 58226
rect 117294 58170 117362 58226
rect 117418 58170 128394 58226
rect 128450 58170 128518 58226
rect 128574 58170 128642 58226
rect 128698 58170 128766 58226
rect 128822 58170 148518 58226
rect 148574 58170 148642 58226
rect 148698 58170 159114 58226
rect 159170 58170 159238 58226
rect 159294 58170 159362 58226
rect 159418 58170 159486 58226
rect 159542 58170 179238 58226
rect 179294 58170 179362 58226
rect 179418 58170 189834 58226
rect 189890 58170 189958 58226
rect 190014 58170 190082 58226
rect 190138 58170 190206 58226
rect 190262 58170 210518 58226
rect 210574 58170 210642 58226
rect 210698 58170 220554 58226
rect 220610 58170 220678 58226
rect 220734 58170 220802 58226
rect 220858 58170 220926 58226
rect 220982 58170 241238 58226
rect 241294 58170 241362 58226
rect 241418 58170 251274 58226
rect 251330 58170 251398 58226
rect 251454 58170 251522 58226
rect 251578 58170 251646 58226
rect 251702 58170 272518 58226
rect 272574 58170 272642 58226
rect 272698 58170 281994 58226
rect 282050 58170 282118 58226
rect 282174 58170 282242 58226
rect 282298 58170 282366 58226
rect 282422 58170 303238 58226
rect 303294 58170 303362 58226
rect 303418 58170 312714 58226
rect 312770 58170 312838 58226
rect 312894 58170 312962 58226
rect 313018 58170 313086 58226
rect 313142 58170 343434 58226
rect 343490 58170 343558 58226
rect 343614 58170 343682 58226
rect 343738 58170 343806 58226
rect 343862 58170 356518 58226
rect 356574 58170 356642 58226
rect 356698 58170 374154 58226
rect 374210 58170 374278 58226
rect 374334 58170 374402 58226
rect 374458 58170 374526 58226
rect 374582 58170 387238 58226
rect 387294 58170 387362 58226
rect 387418 58170 404874 58226
rect 404930 58170 404998 58226
rect 405054 58170 405122 58226
rect 405178 58170 405246 58226
rect 405302 58170 418518 58226
rect 418574 58170 418642 58226
rect 418698 58170 435594 58226
rect 435650 58170 435718 58226
rect 435774 58170 435842 58226
rect 435898 58170 435966 58226
rect 436022 58170 449238 58226
rect 449294 58170 449362 58226
rect 449418 58170 466314 58226
rect 466370 58170 466438 58226
rect 466494 58170 466562 58226
rect 466618 58170 466686 58226
rect 466742 58170 480518 58226
rect 480574 58170 480642 58226
rect 480698 58170 497034 58226
rect 497090 58170 497158 58226
rect 497214 58170 497282 58226
rect 497338 58170 497406 58226
rect 497462 58170 511238 58226
rect 511294 58170 511362 58226
rect 511418 58170 527754 58226
rect 527810 58170 527878 58226
rect 527934 58170 528002 58226
rect 528058 58170 528126 58226
rect 528182 58170 542518 58226
rect 542574 58170 542642 58226
rect 542698 58170 558474 58226
rect 558530 58170 558598 58226
rect 558654 58170 558722 58226
rect 558778 58170 558846 58226
rect 558902 58170 573238 58226
rect 573294 58170 573362 58226
rect 573418 58170 589194 58226
rect 589250 58170 589318 58226
rect 589374 58170 589442 58226
rect 589498 58170 589566 58226
rect 589622 58170 596496 58226
rect 596552 58170 596620 58226
rect 596676 58170 596744 58226
rect 596800 58170 596868 58226
rect 596924 58170 597980 58226
rect -1916 58102 597980 58170
rect -1916 58046 -860 58102
rect -804 58046 -736 58102
rect -680 58046 -612 58102
rect -556 58046 -488 58102
rect -432 58046 5514 58102
rect 5570 58046 5638 58102
rect 5694 58046 5762 58102
rect 5818 58046 5886 58102
rect 5942 58046 24518 58102
rect 24574 58046 24642 58102
rect 24698 58046 36234 58102
rect 36290 58046 36358 58102
rect 36414 58046 36482 58102
rect 36538 58046 36606 58102
rect 36662 58046 55238 58102
rect 55294 58046 55362 58102
rect 55418 58046 66954 58102
rect 67010 58046 67078 58102
rect 67134 58046 67202 58102
rect 67258 58046 67326 58102
rect 67382 58046 86518 58102
rect 86574 58046 86642 58102
rect 86698 58046 97674 58102
rect 97730 58046 97798 58102
rect 97854 58046 97922 58102
rect 97978 58046 98046 58102
rect 98102 58046 117238 58102
rect 117294 58046 117362 58102
rect 117418 58046 128394 58102
rect 128450 58046 128518 58102
rect 128574 58046 128642 58102
rect 128698 58046 128766 58102
rect 128822 58046 148518 58102
rect 148574 58046 148642 58102
rect 148698 58046 159114 58102
rect 159170 58046 159238 58102
rect 159294 58046 159362 58102
rect 159418 58046 159486 58102
rect 159542 58046 179238 58102
rect 179294 58046 179362 58102
rect 179418 58046 189834 58102
rect 189890 58046 189958 58102
rect 190014 58046 190082 58102
rect 190138 58046 190206 58102
rect 190262 58046 210518 58102
rect 210574 58046 210642 58102
rect 210698 58046 220554 58102
rect 220610 58046 220678 58102
rect 220734 58046 220802 58102
rect 220858 58046 220926 58102
rect 220982 58046 241238 58102
rect 241294 58046 241362 58102
rect 241418 58046 251274 58102
rect 251330 58046 251398 58102
rect 251454 58046 251522 58102
rect 251578 58046 251646 58102
rect 251702 58046 272518 58102
rect 272574 58046 272642 58102
rect 272698 58046 281994 58102
rect 282050 58046 282118 58102
rect 282174 58046 282242 58102
rect 282298 58046 282366 58102
rect 282422 58046 303238 58102
rect 303294 58046 303362 58102
rect 303418 58046 312714 58102
rect 312770 58046 312838 58102
rect 312894 58046 312962 58102
rect 313018 58046 313086 58102
rect 313142 58046 343434 58102
rect 343490 58046 343558 58102
rect 343614 58046 343682 58102
rect 343738 58046 343806 58102
rect 343862 58046 356518 58102
rect 356574 58046 356642 58102
rect 356698 58046 374154 58102
rect 374210 58046 374278 58102
rect 374334 58046 374402 58102
rect 374458 58046 374526 58102
rect 374582 58046 387238 58102
rect 387294 58046 387362 58102
rect 387418 58046 404874 58102
rect 404930 58046 404998 58102
rect 405054 58046 405122 58102
rect 405178 58046 405246 58102
rect 405302 58046 418518 58102
rect 418574 58046 418642 58102
rect 418698 58046 435594 58102
rect 435650 58046 435718 58102
rect 435774 58046 435842 58102
rect 435898 58046 435966 58102
rect 436022 58046 449238 58102
rect 449294 58046 449362 58102
rect 449418 58046 466314 58102
rect 466370 58046 466438 58102
rect 466494 58046 466562 58102
rect 466618 58046 466686 58102
rect 466742 58046 480518 58102
rect 480574 58046 480642 58102
rect 480698 58046 497034 58102
rect 497090 58046 497158 58102
rect 497214 58046 497282 58102
rect 497338 58046 497406 58102
rect 497462 58046 511238 58102
rect 511294 58046 511362 58102
rect 511418 58046 527754 58102
rect 527810 58046 527878 58102
rect 527934 58046 528002 58102
rect 528058 58046 528126 58102
rect 528182 58046 542518 58102
rect 542574 58046 542642 58102
rect 542698 58046 558474 58102
rect 558530 58046 558598 58102
rect 558654 58046 558722 58102
rect 558778 58046 558846 58102
rect 558902 58046 573238 58102
rect 573294 58046 573362 58102
rect 573418 58046 589194 58102
rect 589250 58046 589318 58102
rect 589374 58046 589442 58102
rect 589498 58046 589566 58102
rect 589622 58046 596496 58102
rect 596552 58046 596620 58102
rect 596676 58046 596744 58102
rect 596800 58046 596868 58102
rect 596924 58046 597980 58102
rect -1916 57978 597980 58046
rect -1916 57922 -860 57978
rect -804 57922 -736 57978
rect -680 57922 -612 57978
rect -556 57922 -488 57978
rect -432 57922 5514 57978
rect 5570 57922 5638 57978
rect 5694 57922 5762 57978
rect 5818 57922 5886 57978
rect 5942 57922 24518 57978
rect 24574 57922 24642 57978
rect 24698 57922 36234 57978
rect 36290 57922 36358 57978
rect 36414 57922 36482 57978
rect 36538 57922 36606 57978
rect 36662 57922 55238 57978
rect 55294 57922 55362 57978
rect 55418 57922 66954 57978
rect 67010 57922 67078 57978
rect 67134 57922 67202 57978
rect 67258 57922 67326 57978
rect 67382 57922 86518 57978
rect 86574 57922 86642 57978
rect 86698 57922 97674 57978
rect 97730 57922 97798 57978
rect 97854 57922 97922 57978
rect 97978 57922 98046 57978
rect 98102 57922 117238 57978
rect 117294 57922 117362 57978
rect 117418 57922 128394 57978
rect 128450 57922 128518 57978
rect 128574 57922 128642 57978
rect 128698 57922 128766 57978
rect 128822 57922 148518 57978
rect 148574 57922 148642 57978
rect 148698 57922 159114 57978
rect 159170 57922 159238 57978
rect 159294 57922 159362 57978
rect 159418 57922 159486 57978
rect 159542 57922 179238 57978
rect 179294 57922 179362 57978
rect 179418 57922 189834 57978
rect 189890 57922 189958 57978
rect 190014 57922 190082 57978
rect 190138 57922 190206 57978
rect 190262 57922 210518 57978
rect 210574 57922 210642 57978
rect 210698 57922 220554 57978
rect 220610 57922 220678 57978
rect 220734 57922 220802 57978
rect 220858 57922 220926 57978
rect 220982 57922 241238 57978
rect 241294 57922 241362 57978
rect 241418 57922 251274 57978
rect 251330 57922 251398 57978
rect 251454 57922 251522 57978
rect 251578 57922 251646 57978
rect 251702 57922 272518 57978
rect 272574 57922 272642 57978
rect 272698 57922 281994 57978
rect 282050 57922 282118 57978
rect 282174 57922 282242 57978
rect 282298 57922 282366 57978
rect 282422 57922 303238 57978
rect 303294 57922 303362 57978
rect 303418 57922 312714 57978
rect 312770 57922 312838 57978
rect 312894 57922 312962 57978
rect 313018 57922 313086 57978
rect 313142 57922 343434 57978
rect 343490 57922 343558 57978
rect 343614 57922 343682 57978
rect 343738 57922 343806 57978
rect 343862 57922 356518 57978
rect 356574 57922 356642 57978
rect 356698 57922 374154 57978
rect 374210 57922 374278 57978
rect 374334 57922 374402 57978
rect 374458 57922 374526 57978
rect 374582 57922 387238 57978
rect 387294 57922 387362 57978
rect 387418 57922 404874 57978
rect 404930 57922 404998 57978
rect 405054 57922 405122 57978
rect 405178 57922 405246 57978
rect 405302 57922 418518 57978
rect 418574 57922 418642 57978
rect 418698 57922 435594 57978
rect 435650 57922 435718 57978
rect 435774 57922 435842 57978
rect 435898 57922 435966 57978
rect 436022 57922 449238 57978
rect 449294 57922 449362 57978
rect 449418 57922 466314 57978
rect 466370 57922 466438 57978
rect 466494 57922 466562 57978
rect 466618 57922 466686 57978
rect 466742 57922 480518 57978
rect 480574 57922 480642 57978
rect 480698 57922 497034 57978
rect 497090 57922 497158 57978
rect 497214 57922 497282 57978
rect 497338 57922 497406 57978
rect 497462 57922 511238 57978
rect 511294 57922 511362 57978
rect 511418 57922 527754 57978
rect 527810 57922 527878 57978
rect 527934 57922 528002 57978
rect 528058 57922 528126 57978
rect 528182 57922 542518 57978
rect 542574 57922 542642 57978
rect 542698 57922 558474 57978
rect 558530 57922 558598 57978
rect 558654 57922 558722 57978
rect 558778 57922 558846 57978
rect 558902 57922 573238 57978
rect 573294 57922 573362 57978
rect 573418 57922 589194 57978
rect 589250 57922 589318 57978
rect 589374 57922 589442 57978
rect 589498 57922 589566 57978
rect 589622 57922 596496 57978
rect 596552 57922 596620 57978
rect 596676 57922 596744 57978
rect 596800 57922 596868 57978
rect 596924 57922 597980 57978
rect -1916 57826 597980 57922
rect 78916 56278 141108 56294
rect 78916 56222 82684 56278
rect 82740 56222 141036 56278
rect 141092 56222 141108 56278
rect 78916 56206 141108 56222
rect 144044 56278 203268 56294
rect 144044 56222 144060 56278
rect 144116 56222 203196 56278
rect 203252 56222 203268 56278
rect 144044 56206 203268 56222
rect 337636 56278 534340 56294
rect 337636 56222 349356 56278
rect 349412 56222 352716 56278
rect 352772 56222 414652 56278
rect 414708 56222 473676 56278
rect 473732 56222 534268 56278
rect 534324 56222 534340 56278
rect 337636 56206 534340 56222
rect 78916 55574 79004 56206
rect 206092 56098 208364 56114
rect 206092 56042 206108 56098
rect 206164 56042 208364 56098
rect 206092 56026 208364 56042
rect 18380 55558 79004 55574
rect 18380 55502 18396 55558
rect 18452 55502 79004 55558
rect 18380 55486 79004 55502
rect 208276 55574 208364 56026
rect 337636 55574 337724 56206
rect 208276 55558 337724 55574
rect 208276 55502 270060 55558
rect 270116 55502 337724 55558
rect 208276 55486 337724 55502
rect -1916 46350 597980 46446
rect -1916 46294 -1820 46350
rect -1764 46294 -1696 46350
rect -1640 46294 -1572 46350
rect -1516 46294 -1448 46350
rect -1392 46294 9234 46350
rect 9290 46294 9358 46350
rect 9414 46294 9482 46350
rect 9538 46294 9606 46350
rect 9662 46294 39878 46350
rect 39934 46294 40002 46350
rect 40058 46294 70674 46350
rect 70730 46294 70798 46350
rect 70854 46294 70922 46350
rect 70978 46294 71046 46350
rect 71102 46294 101878 46350
rect 101934 46294 102002 46350
rect 102058 46294 132114 46350
rect 132170 46294 132238 46350
rect 132294 46294 132362 46350
rect 132418 46294 132486 46350
rect 132542 46294 162834 46350
rect 162890 46294 162958 46350
rect 163014 46294 163082 46350
rect 163138 46294 163206 46350
rect 163262 46294 163878 46350
rect 163934 46294 164002 46350
rect 164058 46294 193554 46350
rect 193610 46294 193678 46350
rect 193734 46294 193802 46350
rect 193858 46294 193926 46350
rect 193982 46294 224274 46350
rect 224330 46294 224398 46350
rect 224454 46294 224522 46350
rect 224578 46294 224646 46350
rect 224702 46294 225878 46350
rect 225934 46294 226002 46350
rect 226058 46294 254994 46350
rect 255050 46294 255118 46350
rect 255174 46294 255242 46350
rect 255298 46294 255366 46350
rect 255422 46294 285714 46350
rect 285770 46294 285838 46350
rect 285894 46294 285962 46350
rect 286018 46294 286086 46350
rect 286142 46294 287878 46350
rect 287934 46294 288002 46350
rect 288058 46294 316434 46350
rect 316490 46294 316558 46350
rect 316614 46294 316682 46350
rect 316738 46294 316806 46350
rect 316862 46294 318598 46350
rect 318654 46294 318722 46350
rect 318778 46294 347154 46350
rect 347210 46294 347278 46350
rect 347334 46294 347402 46350
rect 347458 46294 347526 46350
rect 347582 46294 371878 46350
rect 371934 46294 372002 46350
rect 372058 46294 377874 46350
rect 377930 46294 377998 46350
rect 378054 46294 378122 46350
rect 378178 46294 378246 46350
rect 378302 46294 408594 46350
rect 408650 46294 408718 46350
rect 408774 46294 408842 46350
rect 408898 46294 408966 46350
rect 409022 46294 433878 46350
rect 433934 46294 434002 46350
rect 434058 46294 439314 46350
rect 439370 46294 439438 46350
rect 439494 46294 439562 46350
rect 439618 46294 439686 46350
rect 439742 46294 470034 46350
rect 470090 46294 470158 46350
rect 470214 46294 470282 46350
rect 470338 46294 470406 46350
rect 470462 46294 495878 46350
rect 495934 46294 496002 46350
rect 496058 46294 500754 46350
rect 500810 46294 500878 46350
rect 500934 46294 501002 46350
rect 501058 46294 501126 46350
rect 501182 46294 531474 46350
rect 531530 46294 531598 46350
rect 531654 46294 531722 46350
rect 531778 46294 531846 46350
rect 531902 46294 557878 46350
rect 557934 46294 558002 46350
rect 558058 46294 562194 46350
rect 562250 46294 562318 46350
rect 562374 46294 562442 46350
rect 562498 46294 562566 46350
rect 562622 46294 592914 46350
rect 592970 46294 593038 46350
rect 593094 46294 593162 46350
rect 593218 46294 593286 46350
rect 593342 46294 597456 46350
rect 597512 46294 597580 46350
rect 597636 46294 597704 46350
rect 597760 46294 597828 46350
rect 597884 46294 597980 46350
rect -1916 46226 597980 46294
rect -1916 46170 -1820 46226
rect -1764 46170 -1696 46226
rect -1640 46170 -1572 46226
rect -1516 46170 -1448 46226
rect -1392 46170 9234 46226
rect 9290 46170 9358 46226
rect 9414 46170 9482 46226
rect 9538 46170 9606 46226
rect 9662 46170 39878 46226
rect 39934 46170 40002 46226
rect 40058 46170 70674 46226
rect 70730 46170 70798 46226
rect 70854 46170 70922 46226
rect 70978 46170 71046 46226
rect 71102 46170 101878 46226
rect 101934 46170 102002 46226
rect 102058 46170 132114 46226
rect 132170 46170 132238 46226
rect 132294 46170 132362 46226
rect 132418 46170 132486 46226
rect 132542 46170 162834 46226
rect 162890 46170 162958 46226
rect 163014 46170 163082 46226
rect 163138 46170 163206 46226
rect 163262 46170 163878 46226
rect 163934 46170 164002 46226
rect 164058 46170 193554 46226
rect 193610 46170 193678 46226
rect 193734 46170 193802 46226
rect 193858 46170 193926 46226
rect 193982 46170 224274 46226
rect 224330 46170 224398 46226
rect 224454 46170 224522 46226
rect 224578 46170 224646 46226
rect 224702 46170 225878 46226
rect 225934 46170 226002 46226
rect 226058 46170 254994 46226
rect 255050 46170 255118 46226
rect 255174 46170 255242 46226
rect 255298 46170 255366 46226
rect 255422 46170 285714 46226
rect 285770 46170 285838 46226
rect 285894 46170 285962 46226
rect 286018 46170 286086 46226
rect 286142 46170 287878 46226
rect 287934 46170 288002 46226
rect 288058 46170 316434 46226
rect 316490 46170 316558 46226
rect 316614 46170 316682 46226
rect 316738 46170 316806 46226
rect 316862 46170 318598 46226
rect 318654 46170 318722 46226
rect 318778 46170 347154 46226
rect 347210 46170 347278 46226
rect 347334 46170 347402 46226
rect 347458 46170 347526 46226
rect 347582 46170 371878 46226
rect 371934 46170 372002 46226
rect 372058 46170 377874 46226
rect 377930 46170 377998 46226
rect 378054 46170 378122 46226
rect 378178 46170 378246 46226
rect 378302 46170 408594 46226
rect 408650 46170 408718 46226
rect 408774 46170 408842 46226
rect 408898 46170 408966 46226
rect 409022 46170 433878 46226
rect 433934 46170 434002 46226
rect 434058 46170 439314 46226
rect 439370 46170 439438 46226
rect 439494 46170 439562 46226
rect 439618 46170 439686 46226
rect 439742 46170 470034 46226
rect 470090 46170 470158 46226
rect 470214 46170 470282 46226
rect 470338 46170 470406 46226
rect 470462 46170 495878 46226
rect 495934 46170 496002 46226
rect 496058 46170 500754 46226
rect 500810 46170 500878 46226
rect 500934 46170 501002 46226
rect 501058 46170 501126 46226
rect 501182 46170 531474 46226
rect 531530 46170 531598 46226
rect 531654 46170 531722 46226
rect 531778 46170 531846 46226
rect 531902 46170 557878 46226
rect 557934 46170 558002 46226
rect 558058 46170 562194 46226
rect 562250 46170 562318 46226
rect 562374 46170 562442 46226
rect 562498 46170 562566 46226
rect 562622 46170 592914 46226
rect 592970 46170 593038 46226
rect 593094 46170 593162 46226
rect 593218 46170 593286 46226
rect 593342 46170 597456 46226
rect 597512 46170 597580 46226
rect 597636 46170 597704 46226
rect 597760 46170 597828 46226
rect 597884 46170 597980 46226
rect -1916 46102 597980 46170
rect -1916 46046 -1820 46102
rect -1764 46046 -1696 46102
rect -1640 46046 -1572 46102
rect -1516 46046 -1448 46102
rect -1392 46046 9234 46102
rect 9290 46046 9358 46102
rect 9414 46046 9482 46102
rect 9538 46046 9606 46102
rect 9662 46046 39878 46102
rect 39934 46046 40002 46102
rect 40058 46046 70674 46102
rect 70730 46046 70798 46102
rect 70854 46046 70922 46102
rect 70978 46046 71046 46102
rect 71102 46046 101878 46102
rect 101934 46046 102002 46102
rect 102058 46046 132114 46102
rect 132170 46046 132238 46102
rect 132294 46046 132362 46102
rect 132418 46046 132486 46102
rect 132542 46046 162834 46102
rect 162890 46046 162958 46102
rect 163014 46046 163082 46102
rect 163138 46046 163206 46102
rect 163262 46046 163878 46102
rect 163934 46046 164002 46102
rect 164058 46046 193554 46102
rect 193610 46046 193678 46102
rect 193734 46046 193802 46102
rect 193858 46046 193926 46102
rect 193982 46046 224274 46102
rect 224330 46046 224398 46102
rect 224454 46046 224522 46102
rect 224578 46046 224646 46102
rect 224702 46046 225878 46102
rect 225934 46046 226002 46102
rect 226058 46046 254994 46102
rect 255050 46046 255118 46102
rect 255174 46046 255242 46102
rect 255298 46046 255366 46102
rect 255422 46046 285714 46102
rect 285770 46046 285838 46102
rect 285894 46046 285962 46102
rect 286018 46046 286086 46102
rect 286142 46046 287878 46102
rect 287934 46046 288002 46102
rect 288058 46046 316434 46102
rect 316490 46046 316558 46102
rect 316614 46046 316682 46102
rect 316738 46046 316806 46102
rect 316862 46046 318598 46102
rect 318654 46046 318722 46102
rect 318778 46046 347154 46102
rect 347210 46046 347278 46102
rect 347334 46046 347402 46102
rect 347458 46046 347526 46102
rect 347582 46046 371878 46102
rect 371934 46046 372002 46102
rect 372058 46046 377874 46102
rect 377930 46046 377998 46102
rect 378054 46046 378122 46102
rect 378178 46046 378246 46102
rect 378302 46046 408594 46102
rect 408650 46046 408718 46102
rect 408774 46046 408842 46102
rect 408898 46046 408966 46102
rect 409022 46046 433878 46102
rect 433934 46046 434002 46102
rect 434058 46046 439314 46102
rect 439370 46046 439438 46102
rect 439494 46046 439562 46102
rect 439618 46046 439686 46102
rect 439742 46046 470034 46102
rect 470090 46046 470158 46102
rect 470214 46046 470282 46102
rect 470338 46046 470406 46102
rect 470462 46046 495878 46102
rect 495934 46046 496002 46102
rect 496058 46046 500754 46102
rect 500810 46046 500878 46102
rect 500934 46046 501002 46102
rect 501058 46046 501126 46102
rect 501182 46046 531474 46102
rect 531530 46046 531598 46102
rect 531654 46046 531722 46102
rect 531778 46046 531846 46102
rect 531902 46046 557878 46102
rect 557934 46046 558002 46102
rect 558058 46046 562194 46102
rect 562250 46046 562318 46102
rect 562374 46046 562442 46102
rect 562498 46046 562566 46102
rect 562622 46046 592914 46102
rect 592970 46046 593038 46102
rect 593094 46046 593162 46102
rect 593218 46046 593286 46102
rect 593342 46046 597456 46102
rect 597512 46046 597580 46102
rect 597636 46046 597704 46102
rect 597760 46046 597828 46102
rect 597884 46046 597980 46102
rect -1916 45978 597980 46046
rect -1916 45922 -1820 45978
rect -1764 45922 -1696 45978
rect -1640 45922 -1572 45978
rect -1516 45922 -1448 45978
rect -1392 45922 9234 45978
rect 9290 45922 9358 45978
rect 9414 45922 9482 45978
rect 9538 45922 9606 45978
rect 9662 45922 39878 45978
rect 39934 45922 40002 45978
rect 40058 45922 70674 45978
rect 70730 45922 70798 45978
rect 70854 45922 70922 45978
rect 70978 45922 71046 45978
rect 71102 45922 101878 45978
rect 101934 45922 102002 45978
rect 102058 45922 132114 45978
rect 132170 45922 132238 45978
rect 132294 45922 132362 45978
rect 132418 45922 132486 45978
rect 132542 45922 162834 45978
rect 162890 45922 162958 45978
rect 163014 45922 163082 45978
rect 163138 45922 163206 45978
rect 163262 45922 163878 45978
rect 163934 45922 164002 45978
rect 164058 45922 193554 45978
rect 193610 45922 193678 45978
rect 193734 45922 193802 45978
rect 193858 45922 193926 45978
rect 193982 45922 224274 45978
rect 224330 45922 224398 45978
rect 224454 45922 224522 45978
rect 224578 45922 224646 45978
rect 224702 45922 225878 45978
rect 225934 45922 226002 45978
rect 226058 45922 254994 45978
rect 255050 45922 255118 45978
rect 255174 45922 255242 45978
rect 255298 45922 255366 45978
rect 255422 45922 285714 45978
rect 285770 45922 285838 45978
rect 285894 45922 285962 45978
rect 286018 45922 286086 45978
rect 286142 45922 287878 45978
rect 287934 45922 288002 45978
rect 288058 45922 316434 45978
rect 316490 45922 316558 45978
rect 316614 45922 316682 45978
rect 316738 45922 316806 45978
rect 316862 45922 318598 45978
rect 318654 45922 318722 45978
rect 318778 45922 347154 45978
rect 347210 45922 347278 45978
rect 347334 45922 347402 45978
rect 347458 45922 347526 45978
rect 347582 45922 371878 45978
rect 371934 45922 372002 45978
rect 372058 45922 377874 45978
rect 377930 45922 377998 45978
rect 378054 45922 378122 45978
rect 378178 45922 378246 45978
rect 378302 45922 408594 45978
rect 408650 45922 408718 45978
rect 408774 45922 408842 45978
rect 408898 45922 408966 45978
rect 409022 45922 433878 45978
rect 433934 45922 434002 45978
rect 434058 45922 439314 45978
rect 439370 45922 439438 45978
rect 439494 45922 439562 45978
rect 439618 45922 439686 45978
rect 439742 45922 470034 45978
rect 470090 45922 470158 45978
rect 470214 45922 470282 45978
rect 470338 45922 470406 45978
rect 470462 45922 495878 45978
rect 495934 45922 496002 45978
rect 496058 45922 500754 45978
rect 500810 45922 500878 45978
rect 500934 45922 501002 45978
rect 501058 45922 501126 45978
rect 501182 45922 531474 45978
rect 531530 45922 531598 45978
rect 531654 45922 531722 45978
rect 531778 45922 531846 45978
rect 531902 45922 557878 45978
rect 557934 45922 558002 45978
rect 558058 45922 562194 45978
rect 562250 45922 562318 45978
rect 562374 45922 562442 45978
rect 562498 45922 562566 45978
rect 562622 45922 592914 45978
rect 592970 45922 593038 45978
rect 593094 45922 593162 45978
rect 593218 45922 593286 45978
rect 593342 45922 597456 45978
rect 597512 45922 597580 45978
rect 597636 45922 597704 45978
rect 597760 45922 597828 45978
rect 597884 45922 597980 45978
rect -1916 45826 597980 45922
rect -1916 40350 597980 40446
rect -1916 40294 -860 40350
rect -804 40294 -736 40350
rect -680 40294 -612 40350
rect -556 40294 -488 40350
rect -432 40294 5514 40350
rect 5570 40294 5638 40350
rect 5694 40294 5762 40350
rect 5818 40294 5886 40350
rect 5942 40294 24518 40350
rect 24574 40294 24642 40350
rect 24698 40294 36234 40350
rect 36290 40294 36358 40350
rect 36414 40294 36482 40350
rect 36538 40294 36606 40350
rect 36662 40294 55238 40350
rect 55294 40294 55362 40350
rect 55418 40294 66954 40350
rect 67010 40294 67078 40350
rect 67134 40294 67202 40350
rect 67258 40294 67326 40350
rect 67382 40294 86518 40350
rect 86574 40294 86642 40350
rect 86698 40294 97674 40350
rect 97730 40294 97798 40350
rect 97854 40294 97922 40350
rect 97978 40294 98046 40350
rect 98102 40294 117238 40350
rect 117294 40294 117362 40350
rect 117418 40294 128394 40350
rect 128450 40294 128518 40350
rect 128574 40294 128642 40350
rect 128698 40294 128766 40350
rect 128822 40294 148518 40350
rect 148574 40294 148642 40350
rect 148698 40294 159114 40350
rect 159170 40294 159238 40350
rect 159294 40294 159362 40350
rect 159418 40294 159486 40350
rect 159542 40294 179238 40350
rect 179294 40294 179362 40350
rect 179418 40294 189834 40350
rect 189890 40294 189958 40350
rect 190014 40294 190082 40350
rect 190138 40294 190206 40350
rect 190262 40294 210518 40350
rect 210574 40294 210642 40350
rect 210698 40294 220554 40350
rect 220610 40294 220678 40350
rect 220734 40294 220802 40350
rect 220858 40294 220926 40350
rect 220982 40294 241238 40350
rect 241294 40294 241362 40350
rect 241418 40294 251274 40350
rect 251330 40294 251398 40350
rect 251454 40294 251522 40350
rect 251578 40294 251646 40350
rect 251702 40294 272518 40350
rect 272574 40294 272642 40350
rect 272698 40294 281994 40350
rect 282050 40294 282118 40350
rect 282174 40294 282242 40350
rect 282298 40294 282366 40350
rect 282422 40294 303238 40350
rect 303294 40294 303362 40350
rect 303418 40294 312714 40350
rect 312770 40294 312838 40350
rect 312894 40294 312962 40350
rect 313018 40294 313086 40350
rect 313142 40294 343434 40350
rect 343490 40294 343558 40350
rect 343614 40294 343682 40350
rect 343738 40294 343806 40350
rect 343862 40294 356518 40350
rect 356574 40294 356642 40350
rect 356698 40294 374154 40350
rect 374210 40294 374278 40350
rect 374334 40294 374402 40350
rect 374458 40294 374526 40350
rect 374582 40294 387238 40350
rect 387294 40294 387362 40350
rect 387418 40294 404874 40350
rect 404930 40294 404998 40350
rect 405054 40294 405122 40350
rect 405178 40294 405246 40350
rect 405302 40294 418518 40350
rect 418574 40294 418642 40350
rect 418698 40294 435594 40350
rect 435650 40294 435718 40350
rect 435774 40294 435842 40350
rect 435898 40294 435966 40350
rect 436022 40294 449238 40350
rect 449294 40294 449362 40350
rect 449418 40294 466314 40350
rect 466370 40294 466438 40350
rect 466494 40294 466562 40350
rect 466618 40294 466686 40350
rect 466742 40294 480518 40350
rect 480574 40294 480642 40350
rect 480698 40294 497034 40350
rect 497090 40294 497158 40350
rect 497214 40294 497282 40350
rect 497338 40294 497406 40350
rect 497462 40294 511238 40350
rect 511294 40294 511362 40350
rect 511418 40294 527754 40350
rect 527810 40294 527878 40350
rect 527934 40294 528002 40350
rect 528058 40294 528126 40350
rect 528182 40294 542518 40350
rect 542574 40294 542642 40350
rect 542698 40294 558474 40350
rect 558530 40294 558598 40350
rect 558654 40294 558722 40350
rect 558778 40294 558846 40350
rect 558902 40294 573238 40350
rect 573294 40294 573362 40350
rect 573418 40294 589194 40350
rect 589250 40294 589318 40350
rect 589374 40294 589442 40350
rect 589498 40294 589566 40350
rect 589622 40294 596496 40350
rect 596552 40294 596620 40350
rect 596676 40294 596744 40350
rect 596800 40294 596868 40350
rect 596924 40294 597980 40350
rect -1916 40226 597980 40294
rect -1916 40170 -860 40226
rect -804 40170 -736 40226
rect -680 40170 -612 40226
rect -556 40170 -488 40226
rect -432 40170 5514 40226
rect 5570 40170 5638 40226
rect 5694 40170 5762 40226
rect 5818 40170 5886 40226
rect 5942 40170 24518 40226
rect 24574 40170 24642 40226
rect 24698 40170 36234 40226
rect 36290 40170 36358 40226
rect 36414 40170 36482 40226
rect 36538 40170 36606 40226
rect 36662 40170 55238 40226
rect 55294 40170 55362 40226
rect 55418 40170 66954 40226
rect 67010 40170 67078 40226
rect 67134 40170 67202 40226
rect 67258 40170 67326 40226
rect 67382 40170 86518 40226
rect 86574 40170 86642 40226
rect 86698 40170 97674 40226
rect 97730 40170 97798 40226
rect 97854 40170 97922 40226
rect 97978 40170 98046 40226
rect 98102 40170 117238 40226
rect 117294 40170 117362 40226
rect 117418 40170 128394 40226
rect 128450 40170 128518 40226
rect 128574 40170 128642 40226
rect 128698 40170 128766 40226
rect 128822 40170 148518 40226
rect 148574 40170 148642 40226
rect 148698 40170 159114 40226
rect 159170 40170 159238 40226
rect 159294 40170 159362 40226
rect 159418 40170 159486 40226
rect 159542 40170 179238 40226
rect 179294 40170 179362 40226
rect 179418 40170 189834 40226
rect 189890 40170 189958 40226
rect 190014 40170 190082 40226
rect 190138 40170 190206 40226
rect 190262 40170 210518 40226
rect 210574 40170 210642 40226
rect 210698 40170 220554 40226
rect 220610 40170 220678 40226
rect 220734 40170 220802 40226
rect 220858 40170 220926 40226
rect 220982 40170 241238 40226
rect 241294 40170 241362 40226
rect 241418 40170 251274 40226
rect 251330 40170 251398 40226
rect 251454 40170 251522 40226
rect 251578 40170 251646 40226
rect 251702 40170 272518 40226
rect 272574 40170 272642 40226
rect 272698 40170 281994 40226
rect 282050 40170 282118 40226
rect 282174 40170 282242 40226
rect 282298 40170 282366 40226
rect 282422 40170 303238 40226
rect 303294 40170 303362 40226
rect 303418 40170 312714 40226
rect 312770 40170 312838 40226
rect 312894 40170 312962 40226
rect 313018 40170 313086 40226
rect 313142 40170 343434 40226
rect 343490 40170 343558 40226
rect 343614 40170 343682 40226
rect 343738 40170 343806 40226
rect 343862 40170 356518 40226
rect 356574 40170 356642 40226
rect 356698 40170 374154 40226
rect 374210 40170 374278 40226
rect 374334 40170 374402 40226
rect 374458 40170 374526 40226
rect 374582 40170 387238 40226
rect 387294 40170 387362 40226
rect 387418 40170 404874 40226
rect 404930 40170 404998 40226
rect 405054 40170 405122 40226
rect 405178 40170 405246 40226
rect 405302 40170 418518 40226
rect 418574 40170 418642 40226
rect 418698 40170 435594 40226
rect 435650 40170 435718 40226
rect 435774 40170 435842 40226
rect 435898 40170 435966 40226
rect 436022 40170 449238 40226
rect 449294 40170 449362 40226
rect 449418 40170 466314 40226
rect 466370 40170 466438 40226
rect 466494 40170 466562 40226
rect 466618 40170 466686 40226
rect 466742 40170 480518 40226
rect 480574 40170 480642 40226
rect 480698 40170 497034 40226
rect 497090 40170 497158 40226
rect 497214 40170 497282 40226
rect 497338 40170 497406 40226
rect 497462 40170 511238 40226
rect 511294 40170 511362 40226
rect 511418 40170 527754 40226
rect 527810 40170 527878 40226
rect 527934 40170 528002 40226
rect 528058 40170 528126 40226
rect 528182 40170 542518 40226
rect 542574 40170 542642 40226
rect 542698 40170 558474 40226
rect 558530 40170 558598 40226
rect 558654 40170 558722 40226
rect 558778 40170 558846 40226
rect 558902 40170 573238 40226
rect 573294 40170 573362 40226
rect 573418 40170 589194 40226
rect 589250 40170 589318 40226
rect 589374 40170 589442 40226
rect 589498 40170 589566 40226
rect 589622 40170 596496 40226
rect 596552 40170 596620 40226
rect 596676 40170 596744 40226
rect 596800 40170 596868 40226
rect 596924 40170 597980 40226
rect -1916 40102 597980 40170
rect -1916 40046 -860 40102
rect -804 40046 -736 40102
rect -680 40046 -612 40102
rect -556 40046 -488 40102
rect -432 40046 5514 40102
rect 5570 40046 5638 40102
rect 5694 40046 5762 40102
rect 5818 40046 5886 40102
rect 5942 40046 24518 40102
rect 24574 40046 24642 40102
rect 24698 40046 36234 40102
rect 36290 40046 36358 40102
rect 36414 40046 36482 40102
rect 36538 40046 36606 40102
rect 36662 40046 55238 40102
rect 55294 40046 55362 40102
rect 55418 40046 66954 40102
rect 67010 40046 67078 40102
rect 67134 40046 67202 40102
rect 67258 40046 67326 40102
rect 67382 40046 86518 40102
rect 86574 40046 86642 40102
rect 86698 40046 97674 40102
rect 97730 40046 97798 40102
rect 97854 40046 97922 40102
rect 97978 40046 98046 40102
rect 98102 40046 117238 40102
rect 117294 40046 117362 40102
rect 117418 40046 128394 40102
rect 128450 40046 128518 40102
rect 128574 40046 128642 40102
rect 128698 40046 128766 40102
rect 128822 40046 148518 40102
rect 148574 40046 148642 40102
rect 148698 40046 159114 40102
rect 159170 40046 159238 40102
rect 159294 40046 159362 40102
rect 159418 40046 159486 40102
rect 159542 40046 179238 40102
rect 179294 40046 179362 40102
rect 179418 40046 189834 40102
rect 189890 40046 189958 40102
rect 190014 40046 190082 40102
rect 190138 40046 190206 40102
rect 190262 40046 210518 40102
rect 210574 40046 210642 40102
rect 210698 40046 220554 40102
rect 220610 40046 220678 40102
rect 220734 40046 220802 40102
rect 220858 40046 220926 40102
rect 220982 40046 241238 40102
rect 241294 40046 241362 40102
rect 241418 40046 251274 40102
rect 251330 40046 251398 40102
rect 251454 40046 251522 40102
rect 251578 40046 251646 40102
rect 251702 40046 272518 40102
rect 272574 40046 272642 40102
rect 272698 40046 281994 40102
rect 282050 40046 282118 40102
rect 282174 40046 282242 40102
rect 282298 40046 282366 40102
rect 282422 40046 303238 40102
rect 303294 40046 303362 40102
rect 303418 40046 312714 40102
rect 312770 40046 312838 40102
rect 312894 40046 312962 40102
rect 313018 40046 313086 40102
rect 313142 40046 343434 40102
rect 343490 40046 343558 40102
rect 343614 40046 343682 40102
rect 343738 40046 343806 40102
rect 343862 40046 356518 40102
rect 356574 40046 356642 40102
rect 356698 40046 374154 40102
rect 374210 40046 374278 40102
rect 374334 40046 374402 40102
rect 374458 40046 374526 40102
rect 374582 40046 387238 40102
rect 387294 40046 387362 40102
rect 387418 40046 404874 40102
rect 404930 40046 404998 40102
rect 405054 40046 405122 40102
rect 405178 40046 405246 40102
rect 405302 40046 418518 40102
rect 418574 40046 418642 40102
rect 418698 40046 435594 40102
rect 435650 40046 435718 40102
rect 435774 40046 435842 40102
rect 435898 40046 435966 40102
rect 436022 40046 449238 40102
rect 449294 40046 449362 40102
rect 449418 40046 466314 40102
rect 466370 40046 466438 40102
rect 466494 40046 466562 40102
rect 466618 40046 466686 40102
rect 466742 40046 480518 40102
rect 480574 40046 480642 40102
rect 480698 40046 497034 40102
rect 497090 40046 497158 40102
rect 497214 40046 497282 40102
rect 497338 40046 497406 40102
rect 497462 40046 511238 40102
rect 511294 40046 511362 40102
rect 511418 40046 527754 40102
rect 527810 40046 527878 40102
rect 527934 40046 528002 40102
rect 528058 40046 528126 40102
rect 528182 40046 542518 40102
rect 542574 40046 542642 40102
rect 542698 40046 558474 40102
rect 558530 40046 558598 40102
rect 558654 40046 558722 40102
rect 558778 40046 558846 40102
rect 558902 40046 573238 40102
rect 573294 40046 573362 40102
rect 573418 40046 589194 40102
rect 589250 40046 589318 40102
rect 589374 40046 589442 40102
rect 589498 40046 589566 40102
rect 589622 40046 596496 40102
rect 596552 40046 596620 40102
rect 596676 40046 596744 40102
rect 596800 40046 596868 40102
rect 596924 40046 597980 40102
rect -1916 39978 597980 40046
rect -1916 39922 -860 39978
rect -804 39922 -736 39978
rect -680 39922 -612 39978
rect -556 39922 -488 39978
rect -432 39922 5514 39978
rect 5570 39922 5638 39978
rect 5694 39922 5762 39978
rect 5818 39922 5886 39978
rect 5942 39922 24518 39978
rect 24574 39922 24642 39978
rect 24698 39922 36234 39978
rect 36290 39922 36358 39978
rect 36414 39922 36482 39978
rect 36538 39922 36606 39978
rect 36662 39922 55238 39978
rect 55294 39922 55362 39978
rect 55418 39922 66954 39978
rect 67010 39922 67078 39978
rect 67134 39922 67202 39978
rect 67258 39922 67326 39978
rect 67382 39922 86518 39978
rect 86574 39922 86642 39978
rect 86698 39922 97674 39978
rect 97730 39922 97798 39978
rect 97854 39922 97922 39978
rect 97978 39922 98046 39978
rect 98102 39922 117238 39978
rect 117294 39922 117362 39978
rect 117418 39922 128394 39978
rect 128450 39922 128518 39978
rect 128574 39922 128642 39978
rect 128698 39922 128766 39978
rect 128822 39922 148518 39978
rect 148574 39922 148642 39978
rect 148698 39922 159114 39978
rect 159170 39922 159238 39978
rect 159294 39922 159362 39978
rect 159418 39922 159486 39978
rect 159542 39922 179238 39978
rect 179294 39922 179362 39978
rect 179418 39922 189834 39978
rect 189890 39922 189958 39978
rect 190014 39922 190082 39978
rect 190138 39922 190206 39978
rect 190262 39922 210518 39978
rect 210574 39922 210642 39978
rect 210698 39922 220554 39978
rect 220610 39922 220678 39978
rect 220734 39922 220802 39978
rect 220858 39922 220926 39978
rect 220982 39922 241238 39978
rect 241294 39922 241362 39978
rect 241418 39922 251274 39978
rect 251330 39922 251398 39978
rect 251454 39922 251522 39978
rect 251578 39922 251646 39978
rect 251702 39922 272518 39978
rect 272574 39922 272642 39978
rect 272698 39922 281994 39978
rect 282050 39922 282118 39978
rect 282174 39922 282242 39978
rect 282298 39922 282366 39978
rect 282422 39922 303238 39978
rect 303294 39922 303362 39978
rect 303418 39922 312714 39978
rect 312770 39922 312838 39978
rect 312894 39922 312962 39978
rect 313018 39922 313086 39978
rect 313142 39922 343434 39978
rect 343490 39922 343558 39978
rect 343614 39922 343682 39978
rect 343738 39922 343806 39978
rect 343862 39922 356518 39978
rect 356574 39922 356642 39978
rect 356698 39922 374154 39978
rect 374210 39922 374278 39978
rect 374334 39922 374402 39978
rect 374458 39922 374526 39978
rect 374582 39922 387238 39978
rect 387294 39922 387362 39978
rect 387418 39922 404874 39978
rect 404930 39922 404998 39978
rect 405054 39922 405122 39978
rect 405178 39922 405246 39978
rect 405302 39922 418518 39978
rect 418574 39922 418642 39978
rect 418698 39922 435594 39978
rect 435650 39922 435718 39978
rect 435774 39922 435842 39978
rect 435898 39922 435966 39978
rect 436022 39922 449238 39978
rect 449294 39922 449362 39978
rect 449418 39922 466314 39978
rect 466370 39922 466438 39978
rect 466494 39922 466562 39978
rect 466618 39922 466686 39978
rect 466742 39922 480518 39978
rect 480574 39922 480642 39978
rect 480698 39922 497034 39978
rect 497090 39922 497158 39978
rect 497214 39922 497282 39978
rect 497338 39922 497406 39978
rect 497462 39922 511238 39978
rect 511294 39922 511362 39978
rect 511418 39922 527754 39978
rect 527810 39922 527878 39978
rect 527934 39922 528002 39978
rect 528058 39922 528126 39978
rect 528182 39922 542518 39978
rect 542574 39922 542642 39978
rect 542698 39922 558474 39978
rect 558530 39922 558598 39978
rect 558654 39922 558722 39978
rect 558778 39922 558846 39978
rect 558902 39922 573238 39978
rect 573294 39922 573362 39978
rect 573418 39922 589194 39978
rect 589250 39922 589318 39978
rect 589374 39922 589442 39978
rect 589498 39922 589566 39978
rect 589622 39922 596496 39978
rect 596552 39922 596620 39978
rect 596676 39922 596744 39978
rect 596800 39922 596868 39978
rect 596924 39922 597980 39978
rect -1916 39826 597980 39922
rect -1916 28350 597980 28446
rect -1916 28294 -1820 28350
rect -1764 28294 -1696 28350
rect -1640 28294 -1572 28350
rect -1516 28294 -1448 28350
rect -1392 28294 9234 28350
rect 9290 28294 9358 28350
rect 9414 28294 9482 28350
rect 9538 28294 9606 28350
rect 9662 28294 39954 28350
rect 40010 28294 40078 28350
rect 40134 28294 40202 28350
rect 40258 28294 40326 28350
rect 40382 28294 70674 28350
rect 70730 28294 70798 28350
rect 70854 28294 70922 28350
rect 70978 28294 71046 28350
rect 71102 28294 101394 28350
rect 101450 28294 101518 28350
rect 101574 28294 101642 28350
rect 101698 28294 101766 28350
rect 101822 28294 132114 28350
rect 132170 28294 132238 28350
rect 132294 28294 132362 28350
rect 132418 28294 132486 28350
rect 132542 28294 162834 28350
rect 162890 28294 162958 28350
rect 163014 28294 163082 28350
rect 163138 28294 163206 28350
rect 163262 28294 193554 28350
rect 193610 28294 193678 28350
rect 193734 28294 193802 28350
rect 193858 28294 193926 28350
rect 193982 28294 224274 28350
rect 224330 28294 224398 28350
rect 224454 28294 224522 28350
rect 224578 28294 224646 28350
rect 224702 28294 254994 28350
rect 255050 28294 255118 28350
rect 255174 28294 255242 28350
rect 255298 28294 255366 28350
rect 255422 28294 285714 28350
rect 285770 28294 285838 28350
rect 285894 28294 285962 28350
rect 286018 28294 286086 28350
rect 286142 28294 316434 28350
rect 316490 28294 316558 28350
rect 316614 28294 316682 28350
rect 316738 28294 316806 28350
rect 316862 28294 347154 28350
rect 347210 28294 347278 28350
rect 347334 28294 347402 28350
rect 347458 28294 347526 28350
rect 347582 28294 377874 28350
rect 377930 28294 377998 28350
rect 378054 28294 378122 28350
rect 378178 28294 378246 28350
rect 378302 28294 408594 28350
rect 408650 28294 408718 28350
rect 408774 28294 408842 28350
rect 408898 28294 408966 28350
rect 409022 28294 439314 28350
rect 439370 28294 439438 28350
rect 439494 28294 439562 28350
rect 439618 28294 439686 28350
rect 439742 28294 470034 28350
rect 470090 28294 470158 28350
rect 470214 28294 470282 28350
rect 470338 28294 470406 28350
rect 470462 28294 500754 28350
rect 500810 28294 500878 28350
rect 500934 28294 501002 28350
rect 501058 28294 501126 28350
rect 501182 28294 531474 28350
rect 531530 28294 531598 28350
rect 531654 28294 531722 28350
rect 531778 28294 531846 28350
rect 531902 28294 562194 28350
rect 562250 28294 562318 28350
rect 562374 28294 562442 28350
rect 562498 28294 562566 28350
rect 562622 28294 592914 28350
rect 592970 28294 593038 28350
rect 593094 28294 593162 28350
rect 593218 28294 593286 28350
rect 593342 28294 597456 28350
rect 597512 28294 597580 28350
rect 597636 28294 597704 28350
rect 597760 28294 597828 28350
rect 597884 28294 597980 28350
rect -1916 28226 597980 28294
rect -1916 28170 -1820 28226
rect -1764 28170 -1696 28226
rect -1640 28170 -1572 28226
rect -1516 28170 -1448 28226
rect -1392 28170 9234 28226
rect 9290 28170 9358 28226
rect 9414 28170 9482 28226
rect 9538 28170 9606 28226
rect 9662 28170 39954 28226
rect 40010 28170 40078 28226
rect 40134 28170 40202 28226
rect 40258 28170 40326 28226
rect 40382 28170 70674 28226
rect 70730 28170 70798 28226
rect 70854 28170 70922 28226
rect 70978 28170 71046 28226
rect 71102 28170 101394 28226
rect 101450 28170 101518 28226
rect 101574 28170 101642 28226
rect 101698 28170 101766 28226
rect 101822 28170 132114 28226
rect 132170 28170 132238 28226
rect 132294 28170 132362 28226
rect 132418 28170 132486 28226
rect 132542 28170 162834 28226
rect 162890 28170 162958 28226
rect 163014 28170 163082 28226
rect 163138 28170 163206 28226
rect 163262 28170 193554 28226
rect 193610 28170 193678 28226
rect 193734 28170 193802 28226
rect 193858 28170 193926 28226
rect 193982 28170 224274 28226
rect 224330 28170 224398 28226
rect 224454 28170 224522 28226
rect 224578 28170 224646 28226
rect 224702 28170 254994 28226
rect 255050 28170 255118 28226
rect 255174 28170 255242 28226
rect 255298 28170 255366 28226
rect 255422 28170 285714 28226
rect 285770 28170 285838 28226
rect 285894 28170 285962 28226
rect 286018 28170 286086 28226
rect 286142 28170 316434 28226
rect 316490 28170 316558 28226
rect 316614 28170 316682 28226
rect 316738 28170 316806 28226
rect 316862 28170 347154 28226
rect 347210 28170 347278 28226
rect 347334 28170 347402 28226
rect 347458 28170 347526 28226
rect 347582 28170 377874 28226
rect 377930 28170 377998 28226
rect 378054 28170 378122 28226
rect 378178 28170 378246 28226
rect 378302 28170 408594 28226
rect 408650 28170 408718 28226
rect 408774 28170 408842 28226
rect 408898 28170 408966 28226
rect 409022 28170 439314 28226
rect 439370 28170 439438 28226
rect 439494 28170 439562 28226
rect 439618 28170 439686 28226
rect 439742 28170 470034 28226
rect 470090 28170 470158 28226
rect 470214 28170 470282 28226
rect 470338 28170 470406 28226
rect 470462 28170 500754 28226
rect 500810 28170 500878 28226
rect 500934 28170 501002 28226
rect 501058 28170 501126 28226
rect 501182 28170 531474 28226
rect 531530 28170 531598 28226
rect 531654 28170 531722 28226
rect 531778 28170 531846 28226
rect 531902 28170 562194 28226
rect 562250 28170 562318 28226
rect 562374 28170 562442 28226
rect 562498 28170 562566 28226
rect 562622 28170 592914 28226
rect 592970 28170 593038 28226
rect 593094 28170 593162 28226
rect 593218 28170 593286 28226
rect 593342 28170 597456 28226
rect 597512 28170 597580 28226
rect 597636 28170 597704 28226
rect 597760 28170 597828 28226
rect 597884 28170 597980 28226
rect -1916 28102 597980 28170
rect -1916 28046 -1820 28102
rect -1764 28046 -1696 28102
rect -1640 28046 -1572 28102
rect -1516 28046 -1448 28102
rect -1392 28046 9234 28102
rect 9290 28046 9358 28102
rect 9414 28046 9482 28102
rect 9538 28046 9606 28102
rect 9662 28046 39954 28102
rect 40010 28046 40078 28102
rect 40134 28046 40202 28102
rect 40258 28046 40326 28102
rect 40382 28046 70674 28102
rect 70730 28046 70798 28102
rect 70854 28046 70922 28102
rect 70978 28046 71046 28102
rect 71102 28046 101394 28102
rect 101450 28046 101518 28102
rect 101574 28046 101642 28102
rect 101698 28046 101766 28102
rect 101822 28046 132114 28102
rect 132170 28046 132238 28102
rect 132294 28046 132362 28102
rect 132418 28046 132486 28102
rect 132542 28046 162834 28102
rect 162890 28046 162958 28102
rect 163014 28046 163082 28102
rect 163138 28046 163206 28102
rect 163262 28046 193554 28102
rect 193610 28046 193678 28102
rect 193734 28046 193802 28102
rect 193858 28046 193926 28102
rect 193982 28046 224274 28102
rect 224330 28046 224398 28102
rect 224454 28046 224522 28102
rect 224578 28046 224646 28102
rect 224702 28046 254994 28102
rect 255050 28046 255118 28102
rect 255174 28046 255242 28102
rect 255298 28046 255366 28102
rect 255422 28046 285714 28102
rect 285770 28046 285838 28102
rect 285894 28046 285962 28102
rect 286018 28046 286086 28102
rect 286142 28046 316434 28102
rect 316490 28046 316558 28102
rect 316614 28046 316682 28102
rect 316738 28046 316806 28102
rect 316862 28046 347154 28102
rect 347210 28046 347278 28102
rect 347334 28046 347402 28102
rect 347458 28046 347526 28102
rect 347582 28046 377874 28102
rect 377930 28046 377998 28102
rect 378054 28046 378122 28102
rect 378178 28046 378246 28102
rect 378302 28046 408594 28102
rect 408650 28046 408718 28102
rect 408774 28046 408842 28102
rect 408898 28046 408966 28102
rect 409022 28046 439314 28102
rect 439370 28046 439438 28102
rect 439494 28046 439562 28102
rect 439618 28046 439686 28102
rect 439742 28046 470034 28102
rect 470090 28046 470158 28102
rect 470214 28046 470282 28102
rect 470338 28046 470406 28102
rect 470462 28046 500754 28102
rect 500810 28046 500878 28102
rect 500934 28046 501002 28102
rect 501058 28046 501126 28102
rect 501182 28046 531474 28102
rect 531530 28046 531598 28102
rect 531654 28046 531722 28102
rect 531778 28046 531846 28102
rect 531902 28046 562194 28102
rect 562250 28046 562318 28102
rect 562374 28046 562442 28102
rect 562498 28046 562566 28102
rect 562622 28046 592914 28102
rect 592970 28046 593038 28102
rect 593094 28046 593162 28102
rect 593218 28046 593286 28102
rect 593342 28046 597456 28102
rect 597512 28046 597580 28102
rect 597636 28046 597704 28102
rect 597760 28046 597828 28102
rect 597884 28046 597980 28102
rect -1916 27978 597980 28046
rect -1916 27922 -1820 27978
rect -1764 27922 -1696 27978
rect -1640 27922 -1572 27978
rect -1516 27922 -1448 27978
rect -1392 27922 9234 27978
rect 9290 27922 9358 27978
rect 9414 27922 9482 27978
rect 9538 27922 9606 27978
rect 9662 27922 39954 27978
rect 40010 27922 40078 27978
rect 40134 27922 40202 27978
rect 40258 27922 40326 27978
rect 40382 27922 70674 27978
rect 70730 27922 70798 27978
rect 70854 27922 70922 27978
rect 70978 27922 71046 27978
rect 71102 27922 101394 27978
rect 101450 27922 101518 27978
rect 101574 27922 101642 27978
rect 101698 27922 101766 27978
rect 101822 27922 132114 27978
rect 132170 27922 132238 27978
rect 132294 27922 132362 27978
rect 132418 27922 132486 27978
rect 132542 27922 162834 27978
rect 162890 27922 162958 27978
rect 163014 27922 163082 27978
rect 163138 27922 163206 27978
rect 163262 27922 193554 27978
rect 193610 27922 193678 27978
rect 193734 27922 193802 27978
rect 193858 27922 193926 27978
rect 193982 27922 224274 27978
rect 224330 27922 224398 27978
rect 224454 27922 224522 27978
rect 224578 27922 224646 27978
rect 224702 27922 254994 27978
rect 255050 27922 255118 27978
rect 255174 27922 255242 27978
rect 255298 27922 255366 27978
rect 255422 27922 285714 27978
rect 285770 27922 285838 27978
rect 285894 27922 285962 27978
rect 286018 27922 286086 27978
rect 286142 27922 316434 27978
rect 316490 27922 316558 27978
rect 316614 27922 316682 27978
rect 316738 27922 316806 27978
rect 316862 27922 347154 27978
rect 347210 27922 347278 27978
rect 347334 27922 347402 27978
rect 347458 27922 347526 27978
rect 347582 27922 377874 27978
rect 377930 27922 377998 27978
rect 378054 27922 378122 27978
rect 378178 27922 378246 27978
rect 378302 27922 408594 27978
rect 408650 27922 408718 27978
rect 408774 27922 408842 27978
rect 408898 27922 408966 27978
rect 409022 27922 439314 27978
rect 439370 27922 439438 27978
rect 439494 27922 439562 27978
rect 439618 27922 439686 27978
rect 439742 27922 470034 27978
rect 470090 27922 470158 27978
rect 470214 27922 470282 27978
rect 470338 27922 470406 27978
rect 470462 27922 500754 27978
rect 500810 27922 500878 27978
rect 500934 27922 501002 27978
rect 501058 27922 501126 27978
rect 501182 27922 531474 27978
rect 531530 27922 531598 27978
rect 531654 27922 531722 27978
rect 531778 27922 531846 27978
rect 531902 27922 562194 27978
rect 562250 27922 562318 27978
rect 562374 27922 562442 27978
rect 562498 27922 562566 27978
rect 562622 27922 592914 27978
rect 592970 27922 593038 27978
rect 593094 27922 593162 27978
rect 593218 27922 593286 27978
rect 593342 27922 597456 27978
rect 597512 27922 597580 27978
rect 597636 27922 597704 27978
rect 597760 27922 597828 27978
rect 597884 27922 597980 27978
rect -1916 27826 597980 27922
rect -1916 22350 597980 22446
rect -1916 22294 -860 22350
rect -804 22294 -736 22350
rect -680 22294 -612 22350
rect -556 22294 -488 22350
rect -432 22294 5514 22350
rect 5570 22294 5638 22350
rect 5694 22294 5762 22350
rect 5818 22294 5886 22350
rect 5942 22294 36234 22350
rect 36290 22294 36358 22350
rect 36414 22294 36482 22350
rect 36538 22294 36606 22350
rect 36662 22294 66954 22350
rect 67010 22294 67078 22350
rect 67134 22294 67202 22350
rect 67258 22294 67326 22350
rect 67382 22294 97674 22350
rect 97730 22294 97798 22350
rect 97854 22294 97922 22350
rect 97978 22294 98046 22350
rect 98102 22294 128394 22350
rect 128450 22294 128518 22350
rect 128574 22294 128642 22350
rect 128698 22294 128766 22350
rect 128822 22294 159114 22350
rect 159170 22294 159238 22350
rect 159294 22294 159362 22350
rect 159418 22294 159486 22350
rect 159542 22294 189834 22350
rect 189890 22294 189958 22350
rect 190014 22294 190082 22350
rect 190138 22294 190206 22350
rect 190262 22294 220554 22350
rect 220610 22294 220678 22350
rect 220734 22294 220802 22350
rect 220858 22294 220926 22350
rect 220982 22294 251274 22350
rect 251330 22294 251398 22350
rect 251454 22294 251522 22350
rect 251578 22294 251646 22350
rect 251702 22294 281994 22350
rect 282050 22294 282118 22350
rect 282174 22294 282242 22350
rect 282298 22294 282366 22350
rect 282422 22294 312714 22350
rect 312770 22294 312838 22350
rect 312894 22294 312962 22350
rect 313018 22294 313086 22350
rect 313142 22294 343434 22350
rect 343490 22294 343558 22350
rect 343614 22294 343682 22350
rect 343738 22294 343806 22350
rect 343862 22294 374154 22350
rect 374210 22294 374278 22350
rect 374334 22294 374402 22350
rect 374458 22294 374526 22350
rect 374582 22294 404874 22350
rect 404930 22294 404998 22350
rect 405054 22294 405122 22350
rect 405178 22294 405246 22350
rect 405302 22294 435594 22350
rect 435650 22294 435718 22350
rect 435774 22294 435842 22350
rect 435898 22294 435966 22350
rect 436022 22294 466314 22350
rect 466370 22294 466438 22350
rect 466494 22294 466562 22350
rect 466618 22294 466686 22350
rect 466742 22294 497034 22350
rect 497090 22294 497158 22350
rect 497214 22294 497282 22350
rect 497338 22294 497406 22350
rect 497462 22294 527754 22350
rect 527810 22294 527878 22350
rect 527934 22294 528002 22350
rect 528058 22294 528126 22350
rect 528182 22294 558474 22350
rect 558530 22294 558598 22350
rect 558654 22294 558722 22350
rect 558778 22294 558846 22350
rect 558902 22294 589194 22350
rect 589250 22294 589318 22350
rect 589374 22294 589442 22350
rect 589498 22294 589566 22350
rect 589622 22294 596496 22350
rect 596552 22294 596620 22350
rect 596676 22294 596744 22350
rect 596800 22294 596868 22350
rect 596924 22294 597980 22350
rect -1916 22226 597980 22294
rect -1916 22170 -860 22226
rect -804 22170 -736 22226
rect -680 22170 -612 22226
rect -556 22170 -488 22226
rect -432 22170 5514 22226
rect 5570 22170 5638 22226
rect 5694 22170 5762 22226
rect 5818 22170 5886 22226
rect 5942 22170 36234 22226
rect 36290 22170 36358 22226
rect 36414 22170 36482 22226
rect 36538 22170 36606 22226
rect 36662 22170 66954 22226
rect 67010 22170 67078 22226
rect 67134 22170 67202 22226
rect 67258 22170 67326 22226
rect 67382 22170 97674 22226
rect 97730 22170 97798 22226
rect 97854 22170 97922 22226
rect 97978 22170 98046 22226
rect 98102 22170 128394 22226
rect 128450 22170 128518 22226
rect 128574 22170 128642 22226
rect 128698 22170 128766 22226
rect 128822 22170 159114 22226
rect 159170 22170 159238 22226
rect 159294 22170 159362 22226
rect 159418 22170 159486 22226
rect 159542 22170 189834 22226
rect 189890 22170 189958 22226
rect 190014 22170 190082 22226
rect 190138 22170 190206 22226
rect 190262 22170 220554 22226
rect 220610 22170 220678 22226
rect 220734 22170 220802 22226
rect 220858 22170 220926 22226
rect 220982 22170 251274 22226
rect 251330 22170 251398 22226
rect 251454 22170 251522 22226
rect 251578 22170 251646 22226
rect 251702 22170 281994 22226
rect 282050 22170 282118 22226
rect 282174 22170 282242 22226
rect 282298 22170 282366 22226
rect 282422 22170 312714 22226
rect 312770 22170 312838 22226
rect 312894 22170 312962 22226
rect 313018 22170 313086 22226
rect 313142 22170 343434 22226
rect 343490 22170 343558 22226
rect 343614 22170 343682 22226
rect 343738 22170 343806 22226
rect 343862 22170 374154 22226
rect 374210 22170 374278 22226
rect 374334 22170 374402 22226
rect 374458 22170 374526 22226
rect 374582 22170 404874 22226
rect 404930 22170 404998 22226
rect 405054 22170 405122 22226
rect 405178 22170 405246 22226
rect 405302 22170 435594 22226
rect 435650 22170 435718 22226
rect 435774 22170 435842 22226
rect 435898 22170 435966 22226
rect 436022 22170 466314 22226
rect 466370 22170 466438 22226
rect 466494 22170 466562 22226
rect 466618 22170 466686 22226
rect 466742 22170 497034 22226
rect 497090 22170 497158 22226
rect 497214 22170 497282 22226
rect 497338 22170 497406 22226
rect 497462 22170 527754 22226
rect 527810 22170 527878 22226
rect 527934 22170 528002 22226
rect 528058 22170 528126 22226
rect 528182 22170 558474 22226
rect 558530 22170 558598 22226
rect 558654 22170 558722 22226
rect 558778 22170 558846 22226
rect 558902 22170 589194 22226
rect 589250 22170 589318 22226
rect 589374 22170 589442 22226
rect 589498 22170 589566 22226
rect 589622 22170 596496 22226
rect 596552 22170 596620 22226
rect 596676 22170 596744 22226
rect 596800 22170 596868 22226
rect 596924 22170 597980 22226
rect -1916 22102 597980 22170
rect -1916 22046 -860 22102
rect -804 22046 -736 22102
rect -680 22046 -612 22102
rect -556 22046 -488 22102
rect -432 22046 5514 22102
rect 5570 22046 5638 22102
rect 5694 22046 5762 22102
rect 5818 22046 5886 22102
rect 5942 22046 36234 22102
rect 36290 22046 36358 22102
rect 36414 22046 36482 22102
rect 36538 22046 36606 22102
rect 36662 22046 66954 22102
rect 67010 22046 67078 22102
rect 67134 22046 67202 22102
rect 67258 22046 67326 22102
rect 67382 22046 97674 22102
rect 97730 22046 97798 22102
rect 97854 22046 97922 22102
rect 97978 22046 98046 22102
rect 98102 22046 128394 22102
rect 128450 22046 128518 22102
rect 128574 22046 128642 22102
rect 128698 22046 128766 22102
rect 128822 22046 159114 22102
rect 159170 22046 159238 22102
rect 159294 22046 159362 22102
rect 159418 22046 159486 22102
rect 159542 22046 189834 22102
rect 189890 22046 189958 22102
rect 190014 22046 190082 22102
rect 190138 22046 190206 22102
rect 190262 22046 220554 22102
rect 220610 22046 220678 22102
rect 220734 22046 220802 22102
rect 220858 22046 220926 22102
rect 220982 22046 251274 22102
rect 251330 22046 251398 22102
rect 251454 22046 251522 22102
rect 251578 22046 251646 22102
rect 251702 22046 281994 22102
rect 282050 22046 282118 22102
rect 282174 22046 282242 22102
rect 282298 22046 282366 22102
rect 282422 22046 312714 22102
rect 312770 22046 312838 22102
rect 312894 22046 312962 22102
rect 313018 22046 313086 22102
rect 313142 22046 343434 22102
rect 343490 22046 343558 22102
rect 343614 22046 343682 22102
rect 343738 22046 343806 22102
rect 343862 22046 374154 22102
rect 374210 22046 374278 22102
rect 374334 22046 374402 22102
rect 374458 22046 374526 22102
rect 374582 22046 404874 22102
rect 404930 22046 404998 22102
rect 405054 22046 405122 22102
rect 405178 22046 405246 22102
rect 405302 22046 435594 22102
rect 435650 22046 435718 22102
rect 435774 22046 435842 22102
rect 435898 22046 435966 22102
rect 436022 22046 466314 22102
rect 466370 22046 466438 22102
rect 466494 22046 466562 22102
rect 466618 22046 466686 22102
rect 466742 22046 497034 22102
rect 497090 22046 497158 22102
rect 497214 22046 497282 22102
rect 497338 22046 497406 22102
rect 497462 22046 527754 22102
rect 527810 22046 527878 22102
rect 527934 22046 528002 22102
rect 528058 22046 528126 22102
rect 528182 22046 558474 22102
rect 558530 22046 558598 22102
rect 558654 22046 558722 22102
rect 558778 22046 558846 22102
rect 558902 22046 589194 22102
rect 589250 22046 589318 22102
rect 589374 22046 589442 22102
rect 589498 22046 589566 22102
rect 589622 22046 596496 22102
rect 596552 22046 596620 22102
rect 596676 22046 596744 22102
rect 596800 22046 596868 22102
rect 596924 22046 597980 22102
rect -1916 21978 597980 22046
rect -1916 21922 -860 21978
rect -804 21922 -736 21978
rect -680 21922 -612 21978
rect -556 21922 -488 21978
rect -432 21922 5514 21978
rect 5570 21922 5638 21978
rect 5694 21922 5762 21978
rect 5818 21922 5886 21978
rect 5942 21922 36234 21978
rect 36290 21922 36358 21978
rect 36414 21922 36482 21978
rect 36538 21922 36606 21978
rect 36662 21922 66954 21978
rect 67010 21922 67078 21978
rect 67134 21922 67202 21978
rect 67258 21922 67326 21978
rect 67382 21922 97674 21978
rect 97730 21922 97798 21978
rect 97854 21922 97922 21978
rect 97978 21922 98046 21978
rect 98102 21922 128394 21978
rect 128450 21922 128518 21978
rect 128574 21922 128642 21978
rect 128698 21922 128766 21978
rect 128822 21922 159114 21978
rect 159170 21922 159238 21978
rect 159294 21922 159362 21978
rect 159418 21922 159486 21978
rect 159542 21922 189834 21978
rect 189890 21922 189958 21978
rect 190014 21922 190082 21978
rect 190138 21922 190206 21978
rect 190262 21922 220554 21978
rect 220610 21922 220678 21978
rect 220734 21922 220802 21978
rect 220858 21922 220926 21978
rect 220982 21922 251274 21978
rect 251330 21922 251398 21978
rect 251454 21922 251522 21978
rect 251578 21922 251646 21978
rect 251702 21922 281994 21978
rect 282050 21922 282118 21978
rect 282174 21922 282242 21978
rect 282298 21922 282366 21978
rect 282422 21922 312714 21978
rect 312770 21922 312838 21978
rect 312894 21922 312962 21978
rect 313018 21922 313086 21978
rect 313142 21922 343434 21978
rect 343490 21922 343558 21978
rect 343614 21922 343682 21978
rect 343738 21922 343806 21978
rect 343862 21922 374154 21978
rect 374210 21922 374278 21978
rect 374334 21922 374402 21978
rect 374458 21922 374526 21978
rect 374582 21922 404874 21978
rect 404930 21922 404998 21978
rect 405054 21922 405122 21978
rect 405178 21922 405246 21978
rect 405302 21922 435594 21978
rect 435650 21922 435718 21978
rect 435774 21922 435842 21978
rect 435898 21922 435966 21978
rect 436022 21922 466314 21978
rect 466370 21922 466438 21978
rect 466494 21922 466562 21978
rect 466618 21922 466686 21978
rect 466742 21922 497034 21978
rect 497090 21922 497158 21978
rect 497214 21922 497282 21978
rect 497338 21922 497406 21978
rect 497462 21922 527754 21978
rect 527810 21922 527878 21978
rect 527934 21922 528002 21978
rect 528058 21922 528126 21978
rect 528182 21922 558474 21978
rect 558530 21922 558598 21978
rect 558654 21922 558722 21978
rect 558778 21922 558846 21978
rect 558902 21922 589194 21978
rect 589250 21922 589318 21978
rect 589374 21922 589442 21978
rect 589498 21922 589566 21978
rect 589622 21922 596496 21978
rect 596552 21922 596620 21978
rect 596676 21922 596744 21978
rect 596800 21922 596868 21978
rect 596924 21922 597980 21978
rect -1916 21826 597980 21922
rect -1916 10350 597980 10446
rect -1916 10294 -1820 10350
rect -1764 10294 -1696 10350
rect -1640 10294 -1572 10350
rect -1516 10294 -1448 10350
rect -1392 10294 9234 10350
rect 9290 10294 9358 10350
rect 9414 10294 9482 10350
rect 9538 10294 9606 10350
rect 9662 10294 39954 10350
rect 40010 10294 40078 10350
rect 40134 10294 40202 10350
rect 40258 10294 40326 10350
rect 40382 10294 70674 10350
rect 70730 10294 70798 10350
rect 70854 10294 70922 10350
rect 70978 10294 71046 10350
rect 71102 10294 101394 10350
rect 101450 10294 101518 10350
rect 101574 10294 101642 10350
rect 101698 10294 101766 10350
rect 101822 10294 132114 10350
rect 132170 10294 132238 10350
rect 132294 10294 132362 10350
rect 132418 10294 132486 10350
rect 132542 10294 162834 10350
rect 162890 10294 162958 10350
rect 163014 10294 163082 10350
rect 163138 10294 163206 10350
rect 163262 10294 193554 10350
rect 193610 10294 193678 10350
rect 193734 10294 193802 10350
rect 193858 10294 193926 10350
rect 193982 10294 224274 10350
rect 224330 10294 224398 10350
rect 224454 10294 224522 10350
rect 224578 10294 224646 10350
rect 224702 10294 254994 10350
rect 255050 10294 255118 10350
rect 255174 10294 255242 10350
rect 255298 10294 255366 10350
rect 255422 10294 285714 10350
rect 285770 10294 285838 10350
rect 285894 10294 285962 10350
rect 286018 10294 286086 10350
rect 286142 10294 316434 10350
rect 316490 10294 316558 10350
rect 316614 10294 316682 10350
rect 316738 10294 316806 10350
rect 316862 10294 347154 10350
rect 347210 10294 347278 10350
rect 347334 10294 347402 10350
rect 347458 10294 347526 10350
rect 347582 10294 377874 10350
rect 377930 10294 377998 10350
rect 378054 10294 378122 10350
rect 378178 10294 378246 10350
rect 378302 10294 408594 10350
rect 408650 10294 408718 10350
rect 408774 10294 408842 10350
rect 408898 10294 408966 10350
rect 409022 10294 439314 10350
rect 439370 10294 439438 10350
rect 439494 10294 439562 10350
rect 439618 10294 439686 10350
rect 439742 10294 470034 10350
rect 470090 10294 470158 10350
rect 470214 10294 470282 10350
rect 470338 10294 470406 10350
rect 470462 10294 500754 10350
rect 500810 10294 500878 10350
rect 500934 10294 501002 10350
rect 501058 10294 501126 10350
rect 501182 10294 531474 10350
rect 531530 10294 531598 10350
rect 531654 10294 531722 10350
rect 531778 10294 531846 10350
rect 531902 10294 562194 10350
rect 562250 10294 562318 10350
rect 562374 10294 562442 10350
rect 562498 10294 562566 10350
rect 562622 10294 592914 10350
rect 592970 10294 593038 10350
rect 593094 10294 593162 10350
rect 593218 10294 593286 10350
rect 593342 10294 597456 10350
rect 597512 10294 597580 10350
rect 597636 10294 597704 10350
rect 597760 10294 597828 10350
rect 597884 10294 597980 10350
rect -1916 10226 597980 10294
rect -1916 10170 -1820 10226
rect -1764 10170 -1696 10226
rect -1640 10170 -1572 10226
rect -1516 10170 -1448 10226
rect -1392 10170 9234 10226
rect 9290 10170 9358 10226
rect 9414 10170 9482 10226
rect 9538 10170 9606 10226
rect 9662 10170 39954 10226
rect 40010 10170 40078 10226
rect 40134 10170 40202 10226
rect 40258 10170 40326 10226
rect 40382 10170 70674 10226
rect 70730 10170 70798 10226
rect 70854 10170 70922 10226
rect 70978 10170 71046 10226
rect 71102 10170 101394 10226
rect 101450 10170 101518 10226
rect 101574 10170 101642 10226
rect 101698 10170 101766 10226
rect 101822 10170 132114 10226
rect 132170 10170 132238 10226
rect 132294 10170 132362 10226
rect 132418 10170 132486 10226
rect 132542 10170 162834 10226
rect 162890 10170 162958 10226
rect 163014 10170 163082 10226
rect 163138 10170 163206 10226
rect 163262 10170 193554 10226
rect 193610 10170 193678 10226
rect 193734 10170 193802 10226
rect 193858 10170 193926 10226
rect 193982 10170 224274 10226
rect 224330 10170 224398 10226
rect 224454 10170 224522 10226
rect 224578 10170 224646 10226
rect 224702 10170 254994 10226
rect 255050 10170 255118 10226
rect 255174 10170 255242 10226
rect 255298 10170 255366 10226
rect 255422 10170 285714 10226
rect 285770 10170 285838 10226
rect 285894 10170 285962 10226
rect 286018 10170 286086 10226
rect 286142 10170 316434 10226
rect 316490 10170 316558 10226
rect 316614 10170 316682 10226
rect 316738 10170 316806 10226
rect 316862 10170 347154 10226
rect 347210 10170 347278 10226
rect 347334 10170 347402 10226
rect 347458 10170 347526 10226
rect 347582 10170 377874 10226
rect 377930 10170 377998 10226
rect 378054 10170 378122 10226
rect 378178 10170 378246 10226
rect 378302 10170 408594 10226
rect 408650 10170 408718 10226
rect 408774 10170 408842 10226
rect 408898 10170 408966 10226
rect 409022 10170 439314 10226
rect 439370 10170 439438 10226
rect 439494 10170 439562 10226
rect 439618 10170 439686 10226
rect 439742 10170 470034 10226
rect 470090 10170 470158 10226
rect 470214 10170 470282 10226
rect 470338 10170 470406 10226
rect 470462 10170 500754 10226
rect 500810 10170 500878 10226
rect 500934 10170 501002 10226
rect 501058 10170 501126 10226
rect 501182 10170 531474 10226
rect 531530 10170 531598 10226
rect 531654 10170 531722 10226
rect 531778 10170 531846 10226
rect 531902 10170 562194 10226
rect 562250 10170 562318 10226
rect 562374 10170 562442 10226
rect 562498 10170 562566 10226
rect 562622 10170 592914 10226
rect 592970 10170 593038 10226
rect 593094 10170 593162 10226
rect 593218 10170 593286 10226
rect 593342 10170 597456 10226
rect 597512 10170 597580 10226
rect 597636 10170 597704 10226
rect 597760 10170 597828 10226
rect 597884 10170 597980 10226
rect -1916 10102 597980 10170
rect -1916 10046 -1820 10102
rect -1764 10046 -1696 10102
rect -1640 10046 -1572 10102
rect -1516 10046 -1448 10102
rect -1392 10046 9234 10102
rect 9290 10046 9358 10102
rect 9414 10046 9482 10102
rect 9538 10046 9606 10102
rect 9662 10046 39954 10102
rect 40010 10046 40078 10102
rect 40134 10046 40202 10102
rect 40258 10046 40326 10102
rect 40382 10046 70674 10102
rect 70730 10046 70798 10102
rect 70854 10046 70922 10102
rect 70978 10046 71046 10102
rect 71102 10046 101394 10102
rect 101450 10046 101518 10102
rect 101574 10046 101642 10102
rect 101698 10046 101766 10102
rect 101822 10046 132114 10102
rect 132170 10046 132238 10102
rect 132294 10046 132362 10102
rect 132418 10046 132486 10102
rect 132542 10046 162834 10102
rect 162890 10046 162958 10102
rect 163014 10046 163082 10102
rect 163138 10046 163206 10102
rect 163262 10046 193554 10102
rect 193610 10046 193678 10102
rect 193734 10046 193802 10102
rect 193858 10046 193926 10102
rect 193982 10046 224274 10102
rect 224330 10046 224398 10102
rect 224454 10046 224522 10102
rect 224578 10046 224646 10102
rect 224702 10046 254994 10102
rect 255050 10046 255118 10102
rect 255174 10046 255242 10102
rect 255298 10046 255366 10102
rect 255422 10046 285714 10102
rect 285770 10046 285838 10102
rect 285894 10046 285962 10102
rect 286018 10046 286086 10102
rect 286142 10046 316434 10102
rect 316490 10046 316558 10102
rect 316614 10046 316682 10102
rect 316738 10046 316806 10102
rect 316862 10046 347154 10102
rect 347210 10046 347278 10102
rect 347334 10046 347402 10102
rect 347458 10046 347526 10102
rect 347582 10046 377874 10102
rect 377930 10046 377998 10102
rect 378054 10046 378122 10102
rect 378178 10046 378246 10102
rect 378302 10046 408594 10102
rect 408650 10046 408718 10102
rect 408774 10046 408842 10102
rect 408898 10046 408966 10102
rect 409022 10046 439314 10102
rect 439370 10046 439438 10102
rect 439494 10046 439562 10102
rect 439618 10046 439686 10102
rect 439742 10046 470034 10102
rect 470090 10046 470158 10102
rect 470214 10046 470282 10102
rect 470338 10046 470406 10102
rect 470462 10046 500754 10102
rect 500810 10046 500878 10102
rect 500934 10046 501002 10102
rect 501058 10046 501126 10102
rect 501182 10046 531474 10102
rect 531530 10046 531598 10102
rect 531654 10046 531722 10102
rect 531778 10046 531846 10102
rect 531902 10046 562194 10102
rect 562250 10046 562318 10102
rect 562374 10046 562442 10102
rect 562498 10046 562566 10102
rect 562622 10046 592914 10102
rect 592970 10046 593038 10102
rect 593094 10046 593162 10102
rect 593218 10046 593286 10102
rect 593342 10046 597456 10102
rect 597512 10046 597580 10102
rect 597636 10046 597704 10102
rect 597760 10046 597828 10102
rect 597884 10046 597980 10102
rect -1916 9978 597980 10046
rect -1916 9922 -1820 9978
rect -1764 9922 -1696 9978
rect -1640 9922 -1572 9978
rect -1516 9922 -1448 9978
rect -1392 9922 9234 9978
rect 9290 9922 9358 9978
rect 9414 9922 9482 9978
rect 9538 9922 9606 9978
rect 9662 9922 39954 9978
rect 40010 9922 40078 9978
rect 40134 9922 40202 9978
rect 40258 9922 40326 9978
rect 40382 9922 70674 9978
rect 70730 9922 70798 9978
rect 70854 9922 70922 9978
rect 70978 9922 71046 9978
rect 71102 9922 101394 9978
rect 101450 9922 101518 9978
rect 101574 9922 101642 9978
rect 101698 9922 101766 9978
rect 101822 9922 132114 9978
rect 132170 9922 132238 9978
rect 132294 9922 132362 9978
rect 132418 9922 132486 9978
rect 132542 9922 162834 9978
rect 162890 9922 162958 9978
rect 163014 9922 163082 9978
rect 163138 9922 163206 9978
rect 163262 9922 193554 9978
rect 193610 9922 193678 9978
rect 193734 9922 193802 9978
rect 193858 9922 193926 9978
rect 193982 9922 224274 9978
rect 224330 9922 224398 9978
rect 224454 9922 224522 9978
rect 224578 9922 224646 9978
rect 224702 9922 254994 9978
rect 255050 9922 255118 9978
rect 255174 9922 255242 9978
rect 255298 9922 255366 9978
rect 255422 9922 285714 9978
rect 285770 9922 285838 9978
rect 285894 9922 285962 9978
rect 286018 9922 286086 9978
rect 286142 9922 316434 9978
rect 316490 9922 316558 9978
rect 316614 9922 316682 9978
rect 316738 9922 316806 9978
rect 316862 9922 347154 9978
rect 347210 9922 347278 9978
rect 347334 9922 347402 9978
rect 347458 9922 347526 9978
rect 347582 9922 377874 9978
rect 377930 9922 377998 9978
rect 378054 9922 378122 9978
rect 378178 9922 378246 9978
rect 378302 9922 408594 9978
rect 408650 9922 408718 9978
rect 408774 9922 408842 9978
rect 408898 9922 408966 9978
rect 409022 9922 439314 9978
rect 439370 9922 439438 9978
rect 439494 9922 439562 9978
rect 439618 9922 439686 9978
rect 439742 9922 470034 9978
rect 470090 9922 470158 9978
rect 470214 9922 470282 9978
rect 470338 9922 470406 9978
rect 470462 9922 500754 9978
rect 500810 9922 500878 9978
rect 500934 9922 501002 9978
rect 501058 9922 501126 9978
rect 501182 9922 531474 9978
rect 531530 9922 531598 9978
rect 531654 9922 531722 9978
rect 531778 9922 531846 9978
rect 531902 9922 562194 9978
rect 562250 9922 562318 9978
rect 562374 9922 562442 9978
rect 562498 9922 562566 9978
rect 562622 9922 592914 9978
rect 592970 9922 593038 9978
rect 593094 9922 593162 9978
rect 593218 9922 593286 9978
rect 593342 9922 597456 9978
rect 597512 9922 597580 9978
rect 597636 9922 597704 9978
rect 597760 9922 597828 9978
rect 597884 9922 597980 9978
rect -1916 9826 597980 9922
rect -1916 4350 597980 4446
rect -1916 4294 -860 4350
rect -804 4294 -736 4350
rect -680 4294 -612 4350
rect -556 4294 -488 4350
rect -432 4294 5514 4350
rect 5570 4294 5638 4350
rect 5694 4294 5762 4350
rect 5818 4294 5886 4350
rect 5942 4294 36234 4350
rect 36290 4294 36358 4350
rect 36414 4294 36482 4350
rect 36538 4294 36606 4350
rect 36662 4294 66954 4350
rect 67010 4294 67078 4350
rect 67134 4294 67202 4350
rect 67258 4294 67326 4350
rect 67382 4294 97674 4350
rect 97730 4294 97798 4350
rect 97854 4294 97922 4350
rect 97978 4294 98046 4350
rect 98102 4294 128394 4350
rect 128450 4294 128518 4350
rect 128574 4294 128642 4350
rect 128698 4294 128766 4350
rect 128822 4294 159114 4350
rect 159170 4294 159238 4350
rect 159294 4294 159362 4350
rect 159418 4294 159486 4350
rect 159542 4294 189834 4350
rect 189890 4294 189958 4350
rect 190014 4294 190082 4350
rect 190138 4294 190206 4350
rect 190262 4294 220554 4350
rect 220610 4294 220678 4350
rect 220734 4294 220802 4350
rect 220858 4294 220926 4350
rect 220982 4294 251274 4350
rect 251330 4294 251398 4350
rect 251454 4294 251522 4350
rect 251578 4294 251646 4350
rect 251702 4294 281994 4350
rect 282050 4294 282118 4350
rect 282174 4294 282242 4350
rect 282298 4294 282366 4350
rect 282422 4294 312714 4350
rect 312770 4294 312838 4350
rect 312894 4294 312962 4350
rect 313018 4294 313086 4350
rect 313142 4294 343434 4350
rect 343490 4294 343558 4350
rect 343614 4294 343682 4350
rect 343738 4294 343806 4350
rect 343862 4294 374154 4350
rect 374210 4294 374278 4350
rect 374334 4294 374402 4350
rect 374458 4294 374526 4350
rect 374582 4294 404874 4350
rect 404930 4294 404998 4350
rect 405054 4294 405122 4350
rect 405178 4294 405246 4350
rect 405302 4294 435594 4350
rect 435650 4294 435718 4350
rect 435774 4294 435842 4350
rect 435898 4294 435966 4350
rect 436022 4294 466314 4350
rect 466370 4294 466438 4350
rect 466494 4294 466562 4350
rect 466618 4294 466686 4350
rect 466742 4294 497034 4350
rect 497090 4294 497158 4350
rect 497214 4294 497282 4350
rect 497338 4294 497406 4350
rect 497462 4294 527754 4350
rect 527810 4294 527878 4350
rect 527934 4294 528002 4350
rect 528058 4294 528126 4350
rect 528182 4294 558474 4350
rect 558530 4294 558598 4350
rect 558654 4294 558722 4350
rect 558778 4294 558846 4350
rect 558902 4294 589194 4350
rect 589250 4294 589318 4350
rect 589374 4294 589442 4350
rect 589498 4294 589566 4350
rect 589622 4294 596496 4350
rect 596552 4294 596620 4350
rect 596676 4294 596744 4350
rect 596800 4294 596868 4350
rect 596924 4294 597980 4350
rect -1916 4226 597980 4294
rect -1916 4170 -860 4226
rect -804 4170 -736 4226
rect -680 4170 -612 4226
rect -556 4170 -488 4226
rect -432 4170 5514 4226
rect 5570 4170 5638 4226
rect 5694 4170 5762 4226
rect 5818 4170 5886 4226
rect 5942 4170 36234 4226
rect 36290 4170 36358 4226
rect 36414 4170 36482 4226
rect 36538 4170 36606 4226
rect 36662 4170 66954 4226
rect 67010 4170 67078 4226
rect 67134 4170 67202 4226
rect 67258 4170 67326 4226
rect 67382 4170 97674 4226
rect 97730 4170 97798 4226
rect 97854 4170 97922 4226
rect 97978 4170 98046 4226
rect 98102 4170 128394 4226
rect 128450 4170 128518 4226
rect 128574 4170 128642 4226
rect 128698 4170 128766 4226
rect 128822 4170 159114 4226
rect 159170 4170 159238 4226
rect 159294 4170 159362 4226
rect 159418 4170 159486 4226
rect 159542 4170 189834 4226
rect 189890 4170 189958 4226
rect 190014 4170 190082 4226
rect 190138 4170 190206 4226
rect 190262 4170 220554 4226
rect 220610 4170 220678 4226
rect 220734 4170 220802 4226
rect 220858 4170 220926 4226
rect 220982 4170 251274 4226
rect 251330 4170 251398 4226
rect 251454 4170 251522 4226
rect 251578 4170 251646 4226
rect 251702 4170 281994 4226
rect 282050 4170 282118 4226
rect 282174 4170 282242 4226
rect 282298 4170 282366 4226
rect 282422 4170 312714 4226
rect 312770 4170 312838 4226
rect 312894 4170 312962 4226
rect 313018 4170 313086 4226
rect 313142 4170 343434 4226
rect 343490 4170 343558 4226
rect 343614 4170 343682 4226
rect 343738 4170 343806 4226
rect 343862 4170 374154 4226
rect 374210 4170 374278 4226
rect 374334 4170 374402 4226
rect 374458 4170 374526 4226
rect 374582 4170 404874 4226
rect 404930 4170 404998 4226
rect 405054 4170 405122 4226
rect 405178 4170 405246 4226
rect 405302 4170 435594 4226
rect 435650 4170 435718 4226
rect 435774 4170 435842 4226
rect 435898 4170 435966 4226
rect 436022 4170 466314 4226
rect 466370 4170 466438 4226
rect 466494 4170 466562 4226
rect 466618 4170 466686 4226
rect 466742 4170 497034 4226
rect 497090 4170 497158 4226
rect 497214 4170 497282 4226
rect 497338 4170 497406 4226
rect 497462 4170 527754 4226
rect 527810 4170 527878 4226
rect 527934 4170 528002 4226
rect 528058 4170 528126 4226
rect 528182 4170 558474 4226
rect 558530 4170 558598 4226
rect 558654 4170 558722 4226
rect 558778 4170 558846 4226
rect 558902 4170 589194 4226
rect 589250 4170 589318 4226
rect 589374 4170 589442 4226
rect 589498 4170 589566 4226
rect 589622 4170 596496 4226
rect 596552 4170 596620 4226
rect 596676 4170 596744 4226
rect 596800 4170 596868 4226
rect 596924 4170 597980 4226
rect -1916 4102 597980 4170
rect -1916 4046 -860 4102
rect -804 4046 -736 4102
rect -680 4046 -612 4102
rect -556 4046 -488 4102
rect -432 4046 5514 4102
rect 5570 4046 5638 4102
rect 5694 4046 5762 4102
rect 5818 4046 5886 4102
rect 5942 4046 36234 4102
rect 36290 4046 36358 4102
rect 36414 4046 36482 4102
rect 36538 4046 36606 4102
rect 36662 4046 66954 4102
rect 67010 4046 67078 4102
rect 67134 4046 67202 4102
rect 67258 4046 67326 4102
rect 67382 4046 97674 4102
rect 97730 4046 97798 4102
rect 97854 4046 97922 4102
rect 97978 4046 98046 4102
rect 98102 4046 128394 4102
rect 128450 4046 128518 4102
rect 128574 4046 128642 4102
rect 128698 4046 128766 4102
rect 128822 4046 159114 4102
rect 159170 4046 159238 4102
rect 159294 4046 159362 4102
rect 159418 4046 159486 4102
rect 159542 4046 189834 4102
rect 189890 4046 189958 4102
rect 190014 4046 190082 4102
rect 190138 4046 190206 4102
rect 190262 4046 220554 4102
rect 220610 4046 220678 4102
rect 220734 4046 220802 4102
rect 220858 4046 220926 4102
rect 220982 4046 251274 4102
rect 251330 4046 251398 4102
rect 251454 4046 251522 4102
rect 251578 4046 251646 4102
rect 251702 4046 281994 4102
rect 282050 4046 282118 4102
rect 282174 4046 282242 4102
rect 282298 4046 282366 4102
rect 282422 4046 312714 4102
rect 312770 4046 312838 4102
rect 312894 4046 312962 4102
rect 313018 4046 313086 4102
rect 313142 4046 343434 4102
rect 343490 4046 343558 4102
rect 343614 4046 343682 4102
rect 343738 4046 343806 4102
rect 343862 4046 374154 4102
rect 374210 4046 374278 4102
rect 374334 4046 374402 4102
rect 374458 4046 374526 4102
rect 374582 4046 404874 4102
rect 404930 4046 404998 4102
rect 405054 4046 405122 4102
rect 405178 4046 405246 4102
rect 405302 4046 435594 4102
rect 435650 4046 435718 4102
rect 435774 4046 435842 4102
rect 435898 4046 435966 4102
rect 436022 4046 466314 4102
rect 466370 4046 466438 4102
rect 466494 4046 466562 4102
rect 466618 4046 466686 4102
rect 466742 4046 497034 4102
rect 497090 4046 497158 4102
rect 497214 4046 497282 4102
rect 497338 4046 497406 4102
rect 497462 4046 527754 4102
rect 527810 4046 527878 4102
rect 527934 4046 528002 4102
rect 528058 4046 528126 4102
rect 528182 4046 558474 4102
rect 558530 4046 558598 4102
rect 558654 4046 558722 4102
rect 558778 4046 558846 4102
rect 558902 4046 589194 4102
rect 589250 4046 589318 4102
rect 589374 4046 589442 4102
rect 589498 4046 589566 4102
rect 589622 4046 596496 4102
rect 596552 4046 596620 4102
rect 596676 4046 596744 4102
rect 596800 4046 596868 4102
rect 596924 4046 597980 4102
rect -1916 3978 597980 4046
rect -1916 3922 -860 3978
rect -804 3922 -736 3978
rect -680 3922 -612 3978
rect -556 3922 -488 3978
rect -432 3922 5514 3978
rect 5570 3922 5638 3978
rect 5694 3922 5762 3978
rect 5818 3922 5886 3978
rect 5942 3922 36234 3978
rect 36290 3922 36358 3978
rect 36414 3922 36482 3978
rect 36538 3922 36606 3978
rect 36662 3922 66954 3978
rect 67010 3922 67078 3978
rect 67134 3922 67202 3978
rect 67258 3922 67326 3978
rect 67382 3922 97674 3978
rect 97730 3922 97798 3978
rect 97854 3922 97922 3978
rect 97978 3922 98046 3978
rect 98102 3922 128394 3978
rect 128450 3922 128518 3978
rect 128574 3922 128642 3978
rect 128698 3922 128766 3978
rect 128822 3922 159114 3978
rect 159170 3922 159238 3978
rect 159294 3922 159362 3978
rect 159418 3922 159486 3978
rect 159542 3922 189834 3978
rect 189890 3922 189958 3978
rect 190014 3922 190082 3978
rect 190138 3922 190206 3978
rect 190262 3922 220554 3978
rect 220610 3922 220678 3978
rect 220734 3922 220802 3978
rect 220858 3922 220926 3978
rect 220982 3922 251274 3978
rect 251330 3922 251398 3978
rect 251454 3922 251522 3978
rect 251578 3922 251646 3978
rect 251702 3922 281994 3978
rect 282050 3922 282118 3978
rect 282174 3922 282242 3978
rect 282298 3922 282366 3978
rect 282422 3922 312714 3978
rect 312770 3922 312838 3978
rect 312894 3922 312962 3978
rect 313018 3922 313086 3978
rect 313142 3922 343434 3978
rect 343490 3922 343558 3978
rect 343614 3922 343682 3978
rect 343738 3922 343806 3978
rect 343862 3922 374154 3978
rect 374210 3922 374278 3978
rect 374334 3922 374402 3978
rect 374458 3922 374526 3978
rect 374582 3922 404874 3978
rect 404930 3922 404998 3978
rect 405054 3922 405122 3978
rect 405178 3922 405246 3978
rect 405302 3922 435594 3978
rect 435650 3922 435718 3978
rect 435774 3922 435842 3978
rect 435898 3922 435966 3978
rect 436022 3922 466314 3978
rect 466370 3922 466438 3978
rect 466494 3922 466562 3978
rect 466618 3922 466686 3978
rect 466742 3922 497034 3978
rect 497090 3922 497158 3978
rect 497214 3922 497282 3978
rect 497338 3922 497406 3978
rect 497462 3922 527754 3978
rect 527810 3922 527878 3978
rect 527934 3922 528002 3978
rect 528058 3922 528126 3978
rect 528182 3922 558474 3978
rect 558530 3922 558598 3978
rect 558654 3922 558722 3978
rect 558778 3922 558846 3978
rect 558902 3922 589194 3978
rect 589250 3922 589318 3978
rect 589374 3922 589442 3978
rect 589498 3922 589566 3978
rect 589622 3922 596496 3978
rect 596552 3922 596620 3978
rect 596676 3922 596744 3978
rect 596800 3922 596868 3978
rect 596924 3922 597980 3978
rect -1916 3826 597980 3922
rect -956 -160 597020 -64
rect -956 -216 -860 -160
rect -804 -216 -736 -160
rect -680 -216 -612 -160
rect -556 -216 -488 -160
rect -432 -216 5514 -160
rect 5570 -216 5638 -160
rect 5694 -216 5762 -160
rect 5818 -216 5886 -160
rect 5942 -216 36234 -160
rect 36290 -216 36358 -160
rect 36414 -216 36482 -160
rect 36538 -216 36606 -160
rect 36662 -216 66954 -160
rect 67010 -216 67078 -160
rect 67134 -216 67202 -160
rect 67258 -216 67326 -160
rect 67382 -216 97674 -160
rect 97730 -216 97798 -160
rect 97854 -216 97922 -160
rect 97978 -216 98046 -160
rect 98102 -216 128394 -160
rect 128450 -216 128518 -160
rect 128574 -216 128642 -160
rect 128698 -216 128766 -160
rect 128822 -216 159114 -160
rect 159170 -216 159238 -160
rect 159294 -216 159362 -160
rect 159418 -216 159486 -160
rect 159542 -216 189834 -160
rect 189890 -216 189958 -160
rect 190014 -216 190082 -160
rect 190138 -216 190206 -160
rect 190262 -216 220554 -160
rect 220610 -216 220678 -160
rect 220734 -216 220802 -160
rect 220858 -216 220926 -160
rect 220982 -216 251274 -160
rect 251330 -216 251398 -160
rect 251454 -216 251522 -160
rect 251578 -216 251646 -160
rect 251702 -216 281994 -160
rect 282050 -216 282118 -160
rect 282174 -216 282242 -160
rect 282298 -216 282366 -160
rect 282422 -216 312714 -160
rect 312770 -216 312838 -160
rect 312894 -216 312962 -160
rect 313018 -216 313086 -160
rect 313142 -216 343434 -160
rect 343490 -216 343558 -160
rect 343614 -216 343682 -160
rect 343738 -216 343806 -160
rect 343862 -216 374154 -160
rect 374210 -216 374278 -160
rect 374334 -216 374402 -160
rect 374458 -216 374526 -160
rect 374582 -216 404874 -160
rect 404930 -216 404998 -160
rect 405054 -216 405122 -160
rect 405178 -216 405246 -160
rect 405302 -216 435594 -160
rect 435650 -216 435718 -160
rect 435774 -216 435842 -160
rect 435898 -216 435966 -160
rect 436022 -216 466314 -160
rect 466370 -216 466438 -160
rect 466494 -216 466562 -160
rect 466618 -216 466686 -160
rect 466742 -216 497034 -160
rect 497090 -216 497158 -160
rect 497214 -216 497282 -160
rect 497338 -216 497406 -160
rect 497462 -216 527754 -160
rect 527810 -216 527878 -160
rect 527934 -216 528002 -160
rect 528058 -216 528126 -160
rect 528182 -216 558474 -160
rect 558530 -216 558598 -160
rect 558654 -216 558722 -160
rect 558778 -216 558846 -160
rect 558902 -216 589194 -160
rect 589250 -216 589318 -160
rect 589374 -216 589442 -160
rect 589498 -216 589566 -160
rect 589622 -216 596496 -160
rect 596552 -216 596620 -160
rect 596676 -216 596744 -160
rect 596800 -216 596868 -160
rect 596924 -216 597020 -160
rect -956 -284 597020 -216
rect -956 -340 -860 -284
rect -804 -340 -736 -284
rect -680 -340 -612 -284
rect -556 -340 -488 -284
rect -432 -340 5514 -284
rect 5570 -340 5638 -284
rect 5694 -340 5762 -284
rect 5818 -340 5886 -284
rect 5942 -340 36234 -284
rect 36290 -340 36358 -284
rect 36414 -340 36482 -284
rect 36538 -340 36606 -284
rect 36662 -340 66954 -284
rect 67010 -340 67078 -284
rect 67134 -340 67202 -284
rect 67258 -340 67326 -284
rect 67382 -340 97674 -284
rect 97730 -340 97798 -284
rect 97854 -340 97922 -284
rect 97978 -340 98046 -284
rect 98102 -340 128394 -284
rect 128450 -340 128518 -284
rect 128574 -340 128642 -284
rect 128698 -340 128766 -284
rect 128822 -340 159114 -284
rect 159170 -340 159238 -284
rect 159294 -340 159362 -284
rect 159418 -340 159486 -284
rect 159542 -340 189834 -284
rect 189890 -340 189958 -284
rect 190014 -340 190082 -284
rect 190138 -340 190206 -284
rect 190262 -340 220554 -284
rect 220610 -340 220678 -284
rect 220734 -340 220802 -284
rect 220858 -340 220926 -284
rect 220982 -340 251274 -284
rect 251330 -340 251398 -284
rect 251454 -340 251522 -284
rect 251578 -340 251646 -284
rect 251702 -340 281994 -284
rect 282050 -340 282118 -284
rect 282174 -340 282242 -284
rect 282298 -340 282366 -284
rect 282422 -340 312714 -284
rect 312770 -340 312838 -284
rect 312894 -340 312962 -284
rect 313018 -340 313086 -284
rect 313142 -340 343434 -284
rect 343490 -340 343558 -284
rect 343614 -340 343682 -284
rect 343738 -340 343806 -284
rect 343862 -340 374154 -284
rect 374210 -340 374278 -284
rect 374334 -340 374402 -284
rect 374458 -340 374526 -284
rect 374582 -340 404874 -284
rect 404930 -340 404998 -284
rect 405054 -340 405122 -284
rect 405178 -340 405246 -284
rect 405302 -340 435594 -284
rect 435650 -340 435718 -284
rect 435774 -340 435842 -284
rect 435898 -340 435966 -284
rect 436022 -340 466314 -284
rect 466370 -340 466438 -284
rect 466494 -340 466562 -284
rect 466618 -340 466686 -284
rect 466742 -340 497034 -284
rect 497090 -340 497158 -284
rect 497214 -340 497282 -284
rect 497338 -340 497406 -284
rect 497462 -340 527754 -284
rect 527810 -340 527878 -284
rect 527934 -340 528002 -284
rect 528058 -340 528126 -284
rect 528182 -340 558474 -284
rect 558530 -340 558598 -284
rect 558654 -340 558722 -284
rect 558778 -340 558846 -284
rect 558902 -340 589194 -284
rect 589250 -340 589318 -284
rect 589374 -340 589442 -284
rect 589498 -340 589566 -284
rect 589622 -340 596496 -284
rect 596552 -340 596620 -284
rect 596676 -340 596744 -284
rect 596800 -340 596868 -284
rect 596924 -340 597020 -284
rect -956 -408 597020 -340
rect -956 -464 -860 -408
rect -804 -464 -736 -408
rect -680 -464 -612 -408
rect -556 -464 -488 -408
rect -432 -464 5514 -408
rect 5570 -464 5638 -408
rect 5694 -464 5762 -408
rect 5818 -464 5886 -408
rect 5942 -464 36234 -408
rect 36290 -464 36358 -408
rect 36414 -464 36482 -408
rect 36538 -464 36606 -408
rect 36662 -464 66954 -408
rect 67010 -464 67078 -408
rect 67134 -464 67202 -408
rect 67258 -464 67326 -408
rect 67382 -464 97674 -408
rect 97730 -464 97798 -408
rect 97854 -464 97922 -408
rect 97978 -464 98046 -408
rect 98102 -464 128394 -408
rect 128450 -464 128518 -408
rect 128574 -464 128642 -408
rect 128698 -464 128766 -408
rect 128822 -464 159114 -408
rect 159170 -464 159238 -408
rect 159294 -464 159362 -408
rect 159418 -464 159486 -408
rect 159542 -464 189834 -408
rect 189890 -464 189958 -408
rect 190014 -464 190082 -408
rect 190138 -464 190206 -408
rect 190262 -464 220554 -408
rect 220610 -464 220678 -408
rect 220734 -464 220802 -408
rect 220858 -464 220926 -408
rect 220982 -464 251274 -408
rect 251330 -464 251398 -408
rect 251454 -464 251522 -408
rect 251578 -464 251646 -408
rect 251702 -464 281994 -408
rect 282050 -464 282118 -408
rect 282174 -464 282242 -408
rect 282298 -464 282366 -408
rect 282422 -464 312714 -408
rect 312770 -464 312838 -408
rect 312894 -464 312962 -408
rect 313018 -464 313086 -408
rect 313142 -464 343434 -408
rect 343490 -464 343558 -408
rect 343614 -464 343682 -408
rect 343738 -464 343806 -408
rect 343862 -464 374154 -408
rect 374210 -464 374278 -408
rect 374334 -464 374402 -408
rect 374458 -464 374526 -408
rect 374582 -464 404874 -408
rect 404930 -464 404998 -408
rect 405054 -464 405122 -408
rect 405178 -464 405246 -408
rect 405302 -464 435594 -408
rect 435650 -464 435718 -408
rect 435774 -464 435842 -408
rect 435898 -464 435966 -408
rect 436022 -464 466314 -408
rect 466370 -464 466438 -408
rect 466494 -464 466562 -408
rect 466618 -464 466686 -408
rect 466742 -464 497034 -408
rect 497090 -464 497158 -408
rect 497214 -464 497282 -408
rect 497338 -464 497406 -408
rect 497462 -464 527754 -408
rect 527810 -464 527878 -408
rect 527934 -464 528002 -408
rect 528058 -464 528126 -408
rect 528182 -464 558474 -408
rect 558530 -464 558598 -408
rect 558654 -464 558722 -408
rect 558778 -464 558846 -408
rect 558902 -464 589194 -408
rect 589250 -464 589318 -408
rect 589374 -464 589442 -408
rect 589498 -464 589566 -408
rect 589622 -464 596496 -408
rect 596552 -464 596620 -408
rect 596676 -464 596744 -408
rect 596800 -464 596868 -408
rect 596924 -464 597020 -408
rect -956 -532 597020 -464
rect -956 -588 -860 -532
rect -804 -588 -736 -532
rect -680 -588 -612 -532
rect -556 -588 -488 -532
rect -432 -588 5514 -532
rect 5570 -588 5638 -532
rect 5694 -588 5762 -532
rect 5818 -588 5886 -532
rect 5942 -588 36234 -532
rect 36290 -588 36358 -532
rect 36414 -588 36482 -532
rect 36538 -588 36606 -532
rect 36662 -588 66954 -532
rect 67010 -588 67078 -532
rect 67134 -588 67202 -532
rect 67258 -588 67326 -532
rect 67382 -588 97674 -532
rect 97730 -588 97798 -532
rect 97854 -588 97922 -532
rect 97978 -588 98046 -532
rect 98102 -588 128394 -532
rect 128450 -588 128518 -532
rect 128574 -588 128642 -532
rect 128698 -588 128766 -532
rect 128822 -588 159114 -532
rect 159170 -588 159238 -532
rect 159294 -588 159362 -532
rect 159418 -588 159486 -532
rect 159542 -588 189834 -532
rect 189890 -588 189958 -532
rect 190014 -588 190082 -532
rect 190138 -588 190206 -532
rect 190262 -588 220554 -532
rect 220610 -588 220678 -532
rect 220734 -588 220802 -532
rect 220858 -588 220926 -532
rect 220982 -588 251274 -532
rect 251330 -588 251398 -532
rect 251454 -588 251522 -532
rect 251578 -588 251646 -532
rect 251702 -588 281994 -532
rect 282050 -588 282118 -532
rect 282174 -588 282242 -532
rect 282298 -588 282366 -532
rect 282422 -588 312714 -532
rect 312770 -588 312838 -532
rect 312894 -588 312962 -532
rect 313018 -588 313086 -532
rect 313142 -588 343434 -532
rect 343490 -588 343558 -532
rect 343614 -588 343682 -532
rect 343738 -588 343806 -532
rect 343862 -588 374154 -532
rect 374210 -588 374278 -532
rect 374334 -588 374402 -532
rect 374458 -588 374526 -532
rect 374582 -588 404874 -532
rect 404930 -588 404998 -532
rect 405054 -588 405122 -532
rect 405178 -588 405246 -532
rect 405302 -588 435594 -532
rect 435650 -588 435718 -532
rect 435774 -588 435842 -532
rect 435898 -588 435966 -532
rect 436022 -588 466314 -532
rect 466370 -588 466438 -532
rect 466494 -588 466562 -532
rect 466618 -588 466686 -532
rect 466742 -588 497034 -532
rect 497090 -588 497158 -532
rect 497214 -588 497282 -532
rect 497338 -588 497406 -532
rect 497462 -588 527754 -532
rect 527810 -588 527878 -532
rect 527934 -588 528002 -532
rect 528058 -588 528126 -532
rect 528182 -588 558474 -532
rect 558530 -588 558598 -532
rect 558654 -588 558722 -532
rect 558778 -588 558846 -532
rect 558902 -588 589194 -532
rect 589250 -588 589318 -532
rect 589374 -588 589442 -532
rect 589498 -588 589566 -532
rect 589622 -588 596496 -532
rect 596552 -588 596620 -532
rect 596676 -588 596744 -532
rect 596800 -588 596868 -532
rect 596924 -588 597020 -532
rect -956 -684 597020 -588
rect -1916 -1120 597980 -1024
rect -1916 -1176 -1820 -1120
rect -1764 -1176 -1696 -1120
rect -1640 -1176 -1572 -1120
rect -1516 -1176 -1448 -1120
rect -1392 -1176 9234 -1120
rect 9290 -1176 9358 -1120
rect 9414 -1176 9482 -1120
rect 9538 -1176 9606 -1120
rect 9662 -1176 39954 -1120
rect 40010 -1176 40078 -1120
rect 40134 -1176 40202 -1120
rect 40258 -1176 40326 -1120
rect 40382 -1176 70674 -1120
rect 70730 -1176 70798 -1120
rect 70854 -1176 70922 -1120
rect 70978 -1176 71046 -1120
rect 71102 -1176 101394 -1120
rect 101450 -1176 101518 -1120
rect 101574 -1176 101642 -1120
rect 101698 -1176 101766 -1120
rect 101822 -1176 132114 -1120
rect 132170 -1176 132238 -1120
rect 132294 -1176 132362 -1120
rect 132418 -1176 132486 -1120
rect 132542 -1176 162834 -1120
rect 162890 -1176 162958 -1120
rect 163014 -1176 163082 -1120
rect 163138 -1176 163206 -1120
rect 163262 -1176 193554 -1120
rect 193610 -1176 193678 -1120
rect 193734 -1176 193802 -1120
rect 193858 -1176 193926 -1120
rect 193982 -1176 224274 -1120
rect 224330 -1176 224398 -1120
rect 224454 -1176 224522 -1120
rect 224578 -1176 224646 -1120
rect 224702 -1176 254994 -1120
rect 255050 -1176 255118 -1120
rect 255174 -1176 255242 -1120
rect 255298 -1176 255366 -1120
rect 255422 -1176 285714 -1120
rect 285770 -1176 285838 -1120
rect 285894 -1176 285962 -1120
rect 286018 -1176 286086 -1120
rect 286142 -1176 316434 -1120
rect 316490 -1176 316558 -1120
rect 316614 -1176 316682 -1120
rect 316738 -1176 316806 -1120
rect 316862 -1176 347154 -1120
rect 347210 -1176 347278 -1120
rect 347334 -1176 347402 -1120
rect 347458 -1176 347526 -1120
rect 347582 -1176 377874 -1120
rect 377930 -1176 377998 -1120
rect 378054 -1176 378122 -1120
rect 378178 -1176 378246 -1120
rect 378302 -1176 408594 -1120
rect 408650 -1176 408718 -1120
rect 408774 -1176 408842 -1120
rect 408898 -1176 408966 -1120
rect 409022 -1176 439314 -1120
rect 439370 -1176 439438 -1120
rect 439494 -1176 439562 -1120
rect 439618 -1176 439686 -1120
rect 439742 -1176 470034 -1120
rect 470090 -1176 470158 -1120
rect 470214 -1176 470282 -1120
rect 470338 -1176 470406 -1120
rect 470462 -1176 500754 -1120
rect 500810 -1176 500878 -1120
rect 500934 -1176 501002 -1120
rect 501058 -1176 501126 -1120
rect 501182 -1176 531474 -1120
rect 531530 -1176 531598 -1120
rect 531654 -1176 531722 -1120
rect 531778 -1176 531846 -1120
rect 531902 -1176 562194 -1120
rect 562250 -1176 562318 -1120
rect 562374 -1176 562442 -1120
rect 562498 -1176 562566 -1120
rect 562622 -1176 592914 -1120
rect 592970 -1176 593038 -1120
rect 593094 -1176 593162 -1120
rect 593218 -1176 593286 -1120
rect 593342 -1176 597456 -1120
rect 597512 -1176 597580 -1120
rect 597636 -1176 597704 -1120
rect 597760 -1176 597828 -1120
rect 597884 -1176 597980 -1120
rect -1916 -1244 597980 -1176
rect -1916 -1300 -1820 -1244
rect -1764 -1300 -1696 -1244
rect -1640 -1300 -1572 -1244
rect -1516 -1300 -1448 -1244
rect -1392 -1300 9234 -1244
rect 9290 -1300 9358 -1244
rect 9414 -1300 9482 -1244
rect 9538 -1300 9606 -1244
rect 9662 -1300 39954 -1244
rect 40010 -1300 40078 -1244
rect 40134 -1300 40202 -1244
rect 40258 -1300 40326 -1244
rect 40382 -1300 70674 -1244
rect 70730 -1300 70798 -1244
rect 70854 -1300 70922 -1244
rect 70978 -1300 71046 -1244
rect 71102 -1300 101394 -1244
rect 101450 -1300 101518 -1244
rect 101574 -1300 101642 -1244
rect 101698 -1300 101766 -1244
rect 101822 -1300 132114 -1244
rect 132170 -1300 132238 -1244
rect 132294 -1300 132362 -1244
rect 132418 -1300 132486 -1244
rect 132542 -1300 162834 -1244
rect 162890 -1300 162958 -1244
rect 163014 -1300 163082 -1244
rect 163138 -1300 163206 -1244
rect 163262 -1300 193554 -1244
rect 193610 -1300 193678 -1244
rect 193734 -1300 193802 -1244
rect 193858 -1300 193926 -1244
rect 193982 -1300 224274 -1244
rect 224330 -1300 224398 -1244
rect 224454 -1300 224522 -1244
rect 224578 -1300 224646 -1244
rect 224702 -1300 254994 -1244
rect 255050 -1300 255118 -1244
rect 255174 -1300 255242 -1244
rect 255298 -1300 255366 -1244
rect 255422 -1300 285714 -1244
rect 285770 -1300 285838 -1244
rect 285894 -1300 285962 -1244
rect 286018 -1300 286086 -1244
rect 286142 -1300 316434 -1244
rect 316490 -1300 316558 -1244
rect 316614 -1300 316682 -1244
rect 316738 -1300 316806 -1244
rect 316862 -1300 347154 -1244
rect 347210 -1300 347278 -1244
rect 347334 -1300 347402 -1244
rect 347458 -1300 347526 -1244
rect 347582 -1300 377874 -1244
rect 377930 -1300 377998 -1244
rect 378054 -1300 378122 -1244
rect 378178 -1300 378246 -1244
rect 378302 -1300 408594 -1244
rect 408650 -1300 408718 -1244
rect 408774 -1300 408842 -1244
rect 408898 -1300 408966 -1244
rect 409022 -1300 439314 -1244
rect 439370 -1300 439438 -1244
rect 439494 -1300 439562 -1244
rect 439618 -1300 439686 -1244
rect 439742 -1300 470034 -1244
rect 470090 -1300 470158 -1244
rect 470214 -1300 470282 -1244
rect 470338 -1300 470406 -1244
rect 470462 -1300 500754 -1244
rect 500810 -1300 500878 -1244
rect 500934 -1300 501002 -1244
rect 501058 -1300 501126 -1244
rect 501182 -1300 531474 -1244
rect 531530 -1300 531598 -1244
rect 531654 -1300 531722 -1244
rect 531778 -1300 531846 -1244
rect 531902 -1300 562194 -1244
rect 562250 -1300 562318 -1244
rect 562374 -1300 562442 -1244
rect 562498 -1300 562566 -1244
rect 562622 -1300 592914 -1244
rect 592970 -1300 593038 -1244
rect 593094 -1300 593162 -1244
rect 593218 -1300 593286 -1244
rect 593342 -1300 597456 -1244
rect 597512 -1300 597580 -1244
rect 597636 -1300 597704 -1244
rect 597760 -1300 597828 -1244
rect 597884 -1300 597980 -1244
rect -1916 -1368 597980 -1300
rect -1916 -1424 -1820 -1368
rect -1764 -1424 -1696 -1368
rect -1640 -1424 -1572 -1368
rect -1516 -1424 -1448 -1368
rect -1392 -1424 9234 -1368
rect 9290 -1424 9358 -1368
rect 9414 -1424 9482 -1368
rect 9538 -1424 9606 -1368
rect 9662 -1424 39954 -1368
rect 40010 -1424 40078 -1368
rect 40134 -1424 40202 -1368
rect 40258 -1424 40326 -1368
rect 40382 -1424 70674 -1368
rect 70730 -1424 70798 -1368
rect 70854 -1424 70922 -1368
rect 70978 -1424 71046 -1368
rect 71102 -1424 101394 -1368
rect 101450 -1424 101518 -1368
rect 101574 -1424 101642 -1368
rect 101698 -1424 101766 -1368
rect 101822 -1424 132114 -1368
rect 132170 -1424 132238 -1368
rect 132294 -1424 132362 -1368
rect 132418 -1424 132486 -1368
rect 132542 -1424 162834 -1368
rect 162890 -1424 162958 -1368
rect 163014 -1424 163082 -1368
rect 163138 -1424 163206 -1368
rect 163262 -1424 193554 -1368
rect 193610 -1424 193678 -1368
rect 193734 -1424 193802 -1368
rect 193858 -1424 193926 -1368
rect 193982 -1424 224274 -1368
rect 224330 -1424 224398 -1368
rect 224454 -1424 224522 -1368
rect 224578 -1424 224646 -1368
rect 224702 -1424 254994 -1368
rect 255050 -1424 255118 -1368
rect 255174 -1424 255242 -1368
rect 255298 -1424 255366 -1368
rect 255422 -1424 285714 -1368
rect 285770 -1424 285838 -1368
rect 285894 -1424 285962 -1368
rect 286018 -1424 286086 -1368
rect 286142 -1424 316434 -1368
rect 316490 -1424 316558 -1368
rect 316614 -1424 316682 -1368
rect 316738 -1424 316806 -1368
rect 316862 -1424 347154 -1368
rect 347210 -1424 347278 -1368
rect 347334 -1424 347402 -1368
rect 347458 -1424 347526 -1368
rect 347582 -1424 377874 -1368
rect 377930 -1424 377998 -1368
rect 378054 -1424 378122 -1368
rect 378178 -1424 378246 -1368
rect 378302 -1424 408594 -1368
rect 408650 -1424 408718 -1368
rect 408774 -1424 408842 -1368
rect 408898 -1424 408966 -1368
rect 409022 -1424 439314 -1368
rect 439370 -1424 439438 -1368
rect 439494 -1424 439562 -1368
rect 439618 -1424 439686 -1368
rect 439742 -1424 470034 -1368
rect 470090 -1424 470158 -1368
rect 470214 -1424 470282 -1368
rect 470338 -1424 470406 -1368
rect 470462 -1424 500754 -1368
rect 500810 -1424 500878 -1368
rect 500934 -1424 501002 -1368
rect 501058 -1424 501126 -1368
rect 501182 -1424 531474 -1368
rect 531530 -1424 531598 -1368
rect 531654 -1424 531722 -1368
rect 531778 -1424 531846 -1368
rect 531902 -1424 562194 -1368
rect 562250 -1424 562318 -1368
rect 562374 -1424 562442 -1368
rect 562498 -1424 562566 -1368
rect 562622 -1424 592914 -1368
rect 592970 -1424 593038 -1368
rect 593094 -1424 593162 -1368
rect 593218 -1424 593286 -1368
rect 593342 -1424 597456 -1368
rect 597512 -1424 597580 -1368
rect 597636 -1424 597704 -1368
rect 597760 -1424 597828 -1368
rect 597884 -1424 597980 -1368
rect -1916 -1492 597980 -1424
rect -1916 -1548 -1820 -1492
rect -1764 -1548 -1696 -1492
rect -1640 -1548 -1572 -1492
rect -1516 -1548 -1448 -1492
rect -1392 -1548 9234 -1492
rect 9290 -1548 9358 -1492
rect 9414 -1548 9482 -1492
rect 9538 -1548 9606 -1492
rect 9662 -1548 39954 -1492
rect 40010 -1548 40078 -1492
rect 40134 -1548 40202 -1492
rect 40258 -1548 40326 -1492
rect 40382 -1548 70674 -1492
rect 70730 -1548 70798 -1492
rect 70854 -1548 70922 -1492
rect 70978 -1548 71046 -1492
rect 71102 -1548 101394 -1492
rect 101450 -1548 101518 -1492
rect 101574 -1548 101642 -1492
rect 101698 -1548 101766 -1492
rect 101822 -1548 132114 -1492
rect 132170 -1548 132238 -1492
rect 132294 -1548 132362 -1492
rect 132418 -1548 132486 -1492
rect 132542 -1548 162834 -1492
rect 162890 -1548 162958 -1492
rect 163014 -1548 163082 -1492
rect 163138 -1548 163206 -1492
rect 163262 -1548 193554 -1492
rect 193610 -1548 193678 -1492
rect 193734 -1548 193802 -1492
rect 193858 -1548 193926 -1492
rect 193982 -1548 224274 -1492
rect 224330 -1548 224398 -1492
rect 224454 -1548 224522 -1492
rect 224578 -1548 224646 -1492
rect 224702 -1548 254994 -1492
rect 255050 -1548 255118 -1492
rect 255174 -1548 255242 -1492
rect 255298 -1548 255366 -1492
rect 255422 -1548 285714 -1492
rect 285770 -1548 285838 -1492
rect 285894 -1548 285962 -1492
rect 286018 -1548 286086 -1492
rect 286142 -1548 316434 -1492
rect 316490 -1548 316558 -1492
rect 316614 -1548 316682 -1492
rect 316738 -1548 316806 -1492
rect 316862 -1548 347154 -1492
rect 347210 -1548 347278 -1492
rect 347334 -1548 347402 -1492
rect 347458 -1548 347526 -1492
rect 347582 -1548 377874 -1492
rect 377930 -1548 377998 -1492
rect 378054 -1548 378122 -1492
rect 378178 -1548 378246 -1492
rect 378302 -1548 408594 -1492
rect 408650 -1548 408718 -1492
rect 408774 -1548 408842 -1492
rect 408898 -1548 408966 -1492
rect 409022 -1548 439314 -1492
rect 439370 -1548 439438 -1492
rect 439494 -1548 439562 -1492
rect 439618 -1548 439686 -1492
rect 439742 -1548 470034 -1492
rect 470090 -1548 470158 -1492
rect 470214 -1548 470282 -1492
rect 470338 -1548 470406 -1492
rect 470462 -1548 500754 -1492
rect 500810 -1548 500878 -1492
rect 500934 -1548 501002 -1492
rect 501058 -1548 501126 -1492
rect 501182 -1548 531474 -1492
rect 531530 -1548 531598 -1492
rect 531654 -1548 531722 -1492
rect 531778 -1548 531846 -1492
rect 531902 -1548 562194 -1492
rect 562250 -1548 562318 -1492
rect 562374 -1548 562442 -1492
rect 562498 -1548 562566 -1492
rect 562622 -1548 592914 -1492
rect 592970 -1548 593038 -1492
rect 593094 -1548 593162 -1492
rect 593218 -1548 593286 -1492
rect 593342 -1548 597456 -1492
rect 597512 -1548 597580 -1492
rect 597636 -1548 597704 -1492
rect 597760 -1548 597828 -1492
rect 597884 -1548 597980 -1492
rect -1916 -1644 597980 -1548
use ita1  ita1
timestamp 0
transform 1 0 20000 0 1 29200
box 0 0 42000 42000
use ita2  ita2
timestamp 0
transform 1 0 82000 0 1 29200
box 0 0 42000 42000
use ita3  ita3
timestamp 0
transform 1 0 144000 0 1 29200
box 0 0 42000 42000
use ita4  ita4
timestamp 0
transform 1 0 206000 0 1 29200
box 0 0 42000 42000
use ita5  ita5
timestamp 0
transform 1 0 352000 0 1 29200
box 0 0 42000 42000
use ita6  ita6
timestamp 0
transform 1 0 414000 0 1 29200
box 0 0 42000 42000
use ita7  ita7
timestamp 0
transform 1 0 476000 0 1 29200
box 0 0 42000 42000
use ita8  ita8
timestamp 0
transform 1 0 538000 0 1 29200
box 0 0 42000 42000
use ita9  ita9
timestamp 0
transform 1 0 20000 0 1 100400
box 0 0 42000 42000
use ita10  ita10
timestamp 0
transform 1 0 82000 0 1 100400
box 0 0 42000 42000
use ita11  ita11
timestamp 0
transform 1 0 144000 0 1 100400
box 0 0 42000 42000
use ita12  ita12
timestamp 0
transform 1 0 206000 0 1 100400
box 0 0 42000 42000
use ita13  ita13
timestamp 0
transform 1 0 352000 0 1 100400
box 0 0 42000 42000
use ita14  ita14
timestamp 0
transform 1 0 414000 0 1 100400
box 0 0 42000 42000
use ita15  ita15
timestamp 0
transform 1 0 476000 0 1 100400
box 0 0 42000 42000
use ita16  ita16
timestamp 0
transform 1 0 538000 0 1 100400
box 0 0 42000 42000
use ita17  ita17
timestamp 0
transform 1 0 20000 0 1 171600
box 0 0 42000 42000
use ita18  ita18
timestamp 0
transform 1 0 82000 0 1 171600
box 0 0 42000 42000
use ita19  ita19
timestamp 0
transform 1 0 144000 0 1 171600
box 0 0 42000 42000
use ita20  ita20
timestamp 0
transform 1 0 206000 0 1 171600
box 0 0 42000 42000
use ita21  ita21
timestamp 0
transform 1 0 352000 0 1 171600
box 0 0 42000 42000
use ita22  ita22
timestamp 0
transform 1 0 414000 0 1 171600
box 0 0 42000 42000
use ita23  ita23
timestamp 0
transform 1 0 476000 0 1 171600
box 0 0 42000 42000
use ita24  ita24
timestamp 0
transform 1 0 538000 0 1 171600
box 0 0 42000 42000
use ita25  ita25
timestamp 0
transform 1 0 20000 0 1 242800
box 0 0 42000 42000
use ita26  ita26
timestamp 0
transform 1 0 82000 0 1 242800
box 0 0 42000 42000
use ita27  ita27
timestamp 0
transform 1 0 144000 0 1 242800
box 0 0 42000 42000
use ita28  ita28
timestamp 0
transform 1 0 206000 0 1 242800
box 0 0 42000 42000
use ita29  ita29
timestamp 0
transform 1 0 352000 0 1 242800
box 0 0 42000 42000
use ita30  ita30
timestamp 0
transform 1 0 414000 0 1 242800
box 0 0 42000 42000
use ita31  ita31
timestamp 0
transform 1 0 476000 0 1 242800
box 0 0 42000 42000
use ita32  ita32
timestamp 0
transform 1 0 538000 0 1 242800
box 0 0 42000 42000
use ita33  ita33
timestamp 0
transform 1 0 20000 0 1 314000
box 0 0 42000 42000
use ita34  ita34
timestamp 0
transform 1 0 82000 0 1 314000
box 0 0 42000 42000
use ita35  ita35
timestamp 0
transform 1 0 144000 0 1 314000
box 0 0 42000 42000
use ita36  ita36
timestamp 0
transform 1 0 206000 0 1 314000
box 0 0 42000 42000
use ita37  ita37
timestamp 0
transform 1 0 352000 0 1 314000
box 0 0 42000 42000
use ita38  ita38
timestamp 0
transform 1 0 414000 0 1 314000
box 0 0 42000 42000
use ita39  ita39
timestamp 0
transform 1 0 476000 0 1 314000
box 0 0 42000 42000
use ita40  ita40
timestamp 0
transform 1 0 538000 0 1 314000
box 0 0 42000 42000
use ita41  ita41
timestamp 0
transform 1 0 20000 0 1 385200
box 0 0 42000 42000
use ita42  ita42
timestamp 0
transform 1 0 82000 0 1 385200
box 0 0 42000 42000
use ita43  ita43
timestamp 0
transform 1 0 144000 0 1 385200
box 0 0 42000 42000
use ita44  ita44
timestamp 0
transform 1 0 206000 0 1 385200
box 0 0 42000 42000
use ita45  ita45
timestamp 0
transform 1 0 352000 0 1 385200
box 0 0 42000 42000
use ita46  ita46
timestamp 0
transform 1 0 414000 0 1 385200
box 0 0 42000 42000
use ita47  ita47
timestamp 0
transform 1 0 476000 0 1 385200
box 0 0 42000 42000
use ita48  ita48
timestamp 0
transform 1 0 538000 0 1 385200
box 0 0 42000 42000
use ita49  ita49
timestamp 0
transform 1 0 20000 0 1 456400
box 0 0 42000 42000
use ita50  ita50
timestamp 0
transform 1 0 82000 0 1 456400
box 0 0 42000 42000
use ita51  ita51
timestamp 0
transform 1 0 144000 0 1 456400
box 0 0 42000 42000
use ita52  ita52
timestamp 0
transform 1 0 206000 0 1 456400
box 0 0 42000 42000
use ita53  ita53
timestamp 0
transform 1 0 352000 0 1 456400
box 0 0 42000 42000
use ita54  ita54
timestamp 0
transform 1 0 414000 0 1 456400
box 0 0 42000 42000
use ita55  ita55
timestamp 0
transform 1 0 476000 0 1 456400
box 0 0 42000 42000
use ita56  ita56
timestamp 0
transform 1 0 538000 0 1 456400
box 0 0 42000 42000
use ita57  ita57
timestamp 0
transform 1 0 20000 0 1 527600
box 0 0 42000 42000
use ita58  ita58
timestamp 0
transform 1 0 82000 0 1 527600
box 0 0 42000 42000
use ita59  ita59
timestamp 0
transform 1 0 144000 0 1 527600
box 0 0 42000 42000
use ita60  ita60
timestamp 0
transform 1 0 206000 0 1 527600
box 0 0 42000 42000
use ita61  ita61
timestamp 0
transform 1 0 352000 0 1 527600
box 0 0 42000 42000
use ita62  ita62
timestamp 0
transform 1 0 414000 0 1 527600
box 0 0 42000 42000
use ita63  ita63
timestamp 0
transform 1 0 476000 0 1 527600
box 0 0 42000 42000
use ita64  ita64
timestamp 0
transform 1 0 538000 0 1 527600
box 0 0 42000 42000
use ita  ita
timestamp 0
transform 1 0 268000 0 1 29200
box 0 0 64000 540400
<< labels >>
flabel metal3 s 595560 7112 597000 7336 0 FreeSans 896 0 0 0 io_in[0]
port 0 nsew signal input
flabel metal3 s 595560 403592 597000 403816 0 FreeSans 896 0 0 0 io_in[10]
port 1 nsew signal input
flabel metal3 s 595560 443240 597000 443464 0 FreeSans 896 0 0 0 io_in[11]
port 2 nsew signal input
flabel metal3 s 595560 482888 597000 483112 0 FreeSans 896 0 0 0 io_in[12]
port 3 nsew signal input
flabel metal3 s 595560 522536 597000 522760 0 FreeSans 896 0 0 0 io_in[13]
port 4 nsew signal input
flabel metal3 s 595560 562184 597000 562408 0 FreeSans 896 0 0 0 io_in[14]
port 5 nsew signal input
flabel metal2 s 584696 595560 584920 597000 0 FreeSans 896 90 0 0 io_in[15]
port 6 nsew signal input
flabel metal2 s 518504 595560 518728 597000 0 FreeSans 896 90 0 0 io_in[16]
port 7 nsew signal input
flabel metal2 s 452312 595560 452536 597000 0 FreeSans 896 90 0 0 io_in[17]
port 8 nsew signal input
flabel metal2 s 386120 595560 386344 597000 0 FreeSans 896 90 0 0 io_in[18]
port 9 nsew signal input
flabel metal2 s 319928 595560 320152 597000 0 FreeSans 896 90 0 0 io_in[19]
port 10 nsew signal input
flabel metal3 s 595560 46760 597000 46984 0 FreeSans 896 0 0 0 io_in[1]
port 11 nsew signal input
flabel metal2 s 253736 595560 253960 597000 0 FreeSans 896 90 0 0 io_in[20]
port 12 nsew signal input
flabel metal2 s 187544 595560 187768 597000 0 FreeSans 896 90 0 0 io_in[21]
port 13 nsew signal input
flabel metal2 s 121352 595560 121576 597000 0 FreeSans 896 90 0 0 io_in[22]
port 14 nsew signal input
flabel metal2 s 55160 595560 55384 597000 0 FreeSans 896 90 0 0 io_in[23]
port 15 nsew signal input
flabel metal3 s -960 587160 480 587384 0 FreeSans 896 0 0 0 io_in[24]
port 16 nsew signal input
flabel metal3 s -960 544824 480 545048 0 FreeSans 896 0 0 0 io_in[25]
port 17 nsew signal input
flabel metal3 s -960 502488 480 502712 0 FreeSans 896 0 0 0 io_in[26]
port 18 nsew signal input
flabel metal3 s -960 460152 480 460376 0 FreeSans 896 0 0 0 io_in[27]
port 19 nsew signal input
flabel metal3 s -960 417816 480 418040 0 FreeSans 896 0 0 0 io_in[28]
port 20 nsew signal input
flabel metal3 s -960 375480 480 375704 0 FreeSans 896 0 0 0 io_in[29]
port 21 nsew signal input
flabel metal3 s 595560 86408 597000 86632 0 FreeSans 896 0 0 0 io_in[2]
port 22 nsew signal input
flabel metal3 s -960 333144 480 333368 0 FreeSans 896 0 0 0 io_in[30]
port 23 nsew signal input
flabel metal3 s -960 290808 480 291032 0 FreeSans 896 0 0 0 io_in[31]
port 24 nsew signal input
flabel metal3 s -960 248472 480 248696 0 FreeSans 896 0 0 0 io_in[32]
port 25 nsew signal input
flabel metal3 s -960 206136 480 206360 0 FreeSans 896 0 0 0 io_in[33]
port 26 nsew signal input
flabel metal3 s -960 163800 480 164024 0 FreeSans 896 0 0 0 io_in[34]
port 27 nsew signal input
flabel metal3 s -960 121464 480 121688 0 FreeSans 896 0 0 0 io_in[35]
port 28 nsew signal input
flabel metal3 s -960 79128 480 79352 0 FreeSans 896 0 0 0 io_in[36]
port 29 nsew signal input
flabel metal3 s -960 36792 480 37016 0 FreeSans 896 0 0 0 io_in[37]
port 30 nsew signal input
flabel metal3 s 595560 126056 597000 126280 0 FreeSans 896 0 0 0 io_in[3]
port 31 nsew signal input
flabel metal3 s 595560 165704 597000 165928 0 FreeSans 896 0 0 0 io_in[4]
port 32 nsew signal input
flabel metal3 s 595560 205352 597000 205576 0 FreeSans 896 0 0 0 io_in[5]
port 33 nsew signal input
flabel metal3 s 595560 245000 597000 245224 0 FreeSans 896 0 0 0 io_in[6]
port 34 nsew signal input
flabel metal3 s 595560 284648 597000 284872 0 FreeSans 896 0 0 0 io_in[7]
port 35 nsew signal input
flabel metal3 s 595560 324296 597000 324520 0 FreeSans 896 0 0 0 io_in[8]
port 36 nsew signal input
flabel metal3 s 595560 363944 597000 364168 0 FreeSans 896 0 0 0 io_in[9]
port 37 nsew signal input
flabel metal3 s 595560 33544 597000 33768 0 FreeSans 896 0 0 0 io_oeb[0]
port 38 nsew signal tristate
flabel metal3 s 595560 430024 597000 430248 0 FreeSans 896 0 0 0 io_oeb[10]
port 39 nsew signal tristate
flabel metal3 s 595560 469672 597000 469896 0 FreeSans 896 0 0 0 io_oeb[11]
port 40 nsew signal tristate
flabel metal3 s 595560 509320 597000 509544 0 FreeSans 896 0 0 0 io_oeb[12]
port 41 nsew signal tristate
flabel metal3 s 595560 548968 597000 549192 0 FreeSans 896 0 0 0 io_oeb[13]
port 42 nsew signal tristate
flabel metal3 s 595560 588616 597000 588840 0 FreeSans 896 0 0 0 io_oeb[14]
port 43 nsew signal tristate
flabel metal2 s 540568 595560 540792 597000 0 FreeSans 896 90 0 0 io_oeb[15]
port 44 nsew signal tristate
flabel metal2 s 474376 595560 474600 597000 0 FreeSans 896 90 0 0 io_oeb[16]
port 45 nsew signal tristate
flabel metal2 s 408184 595560 408408 597000 0 FreeSans 896 90 0 0 io_oeb[17]
port 46 nsew signal tristate
flabel metal2 s 341992 595560 342216 597000 0 FreeSans 896 90 0 0 io_oeb[18]
port 47 nsew signal tristate
flabel metal2 s 275800 595560 276024 597000 0 FreeSans 896 90 0 0 io_oeb[19]
port 48 nsew signal tristate
flabel metal3 s 595560 73192 597000 73416 0 FreeSans 896 0 0 0 io_oeb[1]
port 49 nsew signal tristate
flabel metal2 s 209608 595560 209832 597000 0 FreeSans 896 90 0 0 io_oeb[20]
port 50 nsew signal tristate
flabel metal2 s 143416 595560 143640 597000 0 FreeSans 896 90 0 0 io_oeb[21]
port 51 nsew signal tristate
flabel metal2 s 77224 595560 77448 597000 0 FreeSans 896 90 0 0 io_oeb[22]
port 52 nsew signal tristate
flabel metal2 s 11032 595560 11256 597000 0 FreeSans 896 90 0 0 io_oeb[23]
port 53 nsew signal tristate
flabel metal3 s -960 558936 480 559160 0 FreeSans 896 0 0 0 io_oeb[24]
port 54 nsew signal tristate
flabel metal3 s -960 516600 480 516824 0 FreeSans 896 0 0 0 io_oeb[25]
port 55 nsew signal tristate
flabel metal3 s -960 474264 480 474488 0 FreeSans 896 0 0 0 io_oeb[26]
port 56 nsew signal tristate
flabel metal3 s -960 431928 480 432152 0 FreeSans 896 0 0 0 io_oeb[27]
port 57 nsew signal tristate
flabel metal3 s -960 389592 480 389816 0 FreeSans 896 0 0 0 io_oeb[28]
port 58 nsew signal tristate
flabel metal3 s -960 347256 480 347480 0 FreeSans 896 0 0 0 io_oeb[29]
port 59 nsew signal tristate
flabel metal3 s 595560 112840 597000 113064 0 FreeSans 896 0 0 0 io_oeb[2]
port 60 nsew signal tristate
flabel metal3 s -960 304920 480 305144 0 FreeSans 896 0 0 0 io_oeb[30]
port 61 nsew signal tristate
flabel metal3 s -960 262584 480 262808 0 FreeSans 896 0 0 0 io_oeb[31]
port 62 nsew signal tristate
flabel metal3 s -960 220248 480 220472 0 FreeSans 896 0 0 0 io_oeb[32]
port 63 nsew signal tristate
flabel metal3 s -960 177912 480 178136 0 FreeSans 896 0 0 0 io_oeb[33]
port 64 nsew signal tristate
flabel metal3 s -960 135576 480 135800 0 FreeSans 896 0 0 0 io_oeb[34]
port 65 nsew signal tristate
flabel metal3 s -960 93240 480 93464 0 FreeSans 896 0 0 0 io_oeb[35]
port 66 nsew signal tristate
flabel metal3 s -960 50904 480 51128 0 FreeSans 896 0 0 0 io_oeb[36]
port 67 nsew signal tristate
flabel metal3 s -960 8568 480 8792 0 FreeSans 896 0 0 0 io_oeb[37]
port 68 nsew signal tristate
flabel metal3 s 595560 152488 597000 152712 0 FreeSans 896 0 0 0 io_oeb[3]
port 69 nsew signal tristate
flabel metal3 s 595560 192136 597000 192360 0 FreeSans 896 0 0 0 io_oeb[4]
port 70 nsew signal tristate
flabel metal3 s 595560 231784 597000 232008 0 FreeSans 896 0 0 0 io_oeb[5]
port 71 nsew signal tristate
flabel metal3 s 595560 271432 597000 271656 0 FreeSans 896 0 0 0 io_oeb[6]
port 72 nsew signal tristate
flabel metal3 s 595560 311080 597000 311304 0 FreeSans 896 0 0 0 io_oeb[7]
port 73 nsew signal tristate
flabel metal3 s 595560 350728 597000 350952 0 FreeSans 896 0 0 0 io_oeb[8]
port 74 nsew signal tristate
flabel metal3 s 595560 390376 597000 390600 0 FreeSans 896 0 0 0 io_oeb[9]
port 75 nsew signal tristate
flabel metal3 s 595560 20328 597000 20552 0 FreeSans 896 0 0 0 io_out[0]
port 76 nsew signal tristate
flabel metal3 s 595560 416808 597000 417032 0 FreeSans 896 0 0 0 io_out[10]
port 77 nsew signal tristate
flabel metal3 s 595560 456456 597000 456680 0 FreeSans 896 0 0 0 io_out[11]
port 78 nsew signal tristate
flabel metal3 s 595560 496104 597000 496328 0 FreeSans 896 0 0 0 io_out[12]
port 79 nsew signal tristate
flabel metal3 s 595560 535752 597000 535976 0 FreeSans 896 0 0 0 io_out[13]
port 80 nsew signal tristate
flabel metal3 s 595560 575400 597000 575624 0 FreeSans 896 0 0 0 io_out[14]
port 81 nsew signal tristate
flabel metal2 s 562632 595560 562856 597000 0 FreeSans 896 90 0 0 io_out[15]
port 82 nsew signal tristate
flabel metal2 s 496440 595560 496664 597000 0 FreeSans 896 90 0 0 io_out[16]
port 83 nsew signal tristate
flabel metal2 s 430248 595560 430472 597000 0 FreeSans 896 90 0 0 io_out[17]
port 84 nsew signal tristate
flabel metal2 s 364056 595560 364280 597000 0 FreeSans 896 90 0 0 io_out[18]
port 85 nsew signal tristate
flabel metal2 s 297864 595560 298088 597000 0 FreeSans 896 90 0 0 io_out[19]
port 86 nsew signal tristate
flabel metal3 s 595560 59976 597000 60200 0 FreeSans 896 0 0 0 io_out[1]
port 87 nsew signal tristate
flabel metal2 s 231672 595560 231896 597000 0 FreeSans 896 90 0 0 io_out[20]
port 88 nsew signal tristate
flabel metal2 s 165480 595560 165704 597000 0 FreeSans 896 90 0 0 io_out[21]
port 89 nsew signal tristate
flabel metal2 s 99288 595560 99512 597000 0 FreeSans 896 90 0 0 io_out[22]
port 90 nsew signal tristate
flabel metal2 s 33096 595560 33320 597000 0 FreeSans 896 90 0 0 io_out[23]
port 91 nsew signal tristate
flabel metal3 s -960 573048 480 573272 0 FreeSans 896 0 0 0 io_out[24]
port 92 nsew signal tristate
flabel metal3 s -960 530712 480 530936 0 FreeSans 896 0 0 0 io_out[25]
port 93 nsew signal tristate
flabel metal3 s -960 488376 480 488600 0 FreeSans 896 0 0 0 io_out[26]
port 94 nsew signal tristate
flabel metal3 s -960 446040 480 446264 0 FreeSans 896 0 0 0 io_out[27]
port 95 nsew signal tristate
flabel metal3 s -960 403704 480 403928 0 FreeSans 896 0 0 0 io_out[28]
port 96 nsew signal tristate
flabel metal3 s -960 361368 480 361592 0 FreeSans 896 0 0 0 io_out[29]
port 97 nsew signal tristate
flabel metal3 s 595560 99624 597000 99848 0 FreeSans 896 0 0 0 io_out[2]
port 98 nsew signal tristate
flabel metal3 s -960 319032 480 319256 0 FreeSans 896 0 0 0 io_out[30]
port 99 nsew signal tristate
flabel metal3 s -960 276696 480 276920 0 FreeSans 896 0 0 0 io_out[31]
port 100 nsew signal tristate
flabel metal3 s -960 234360 480 234584 0 FreeSans 896 0 0 0 io_out[32]
port 101 nsew signal tristate
flabel metal3 s -960 192024 480 192248 0 FreeSans 896 0 0 0 io_out[33]
port 102 nsew signal tristate
flabel metal3 s -960 149688 480 149912 0 FreeSans 896 0 0 0 io_out[34]
port 103 nsew signal tristate
flabel metal3 s -960 107352 480 107576 0 FreeSans 896 0 0 0 io_out[35]
port 104 nsew signal tristate
flabel metal3 s -960 65016 480 65240 0 FreeSans 896 0 0 0 io_out[36]
port 105 nsew signal tristate
flabel metal3 s -960 22680 480 22904 0 FreeSans 896 0 0 0 io_out[37]
port 106 nsew signal tristate
flabel metal3 s 595560 139272 597000 139496 0 FreeSans 896 0 0 0 io_out[3]
port 107 nsew signal tristate
flabel metal3 s 595560 178920 597000 179144 0 FreeSans 896 0 0 0 io_out[4]
port 108 nsew signal tristate
flabel metal3 s 595560 218568 597000 218792 0 FreeSans 896 0 0 0 io_out[5]
port 109 nsew signal tristate
flabel metal3 s 595560 258216 597000 258440 0 FreeSans 896 0 0 0 io_out[6]
port 110 nsew signal tristate
flabel metal3 s 595560 297864 597000 298088 0 FreeSans 896 0 0 0 io_out[7]
port 111 nsew signal tristate
flabel metal3 s 595560 337512 597000 337736 0 FreeSans 896 0 0 0 io_out[8]
port 112 nsew signal tristate
flabel metal3 s 595560 377160 597000 377384 0 FreeSans 896 0 0 0 io_out[9]
port 113 nsew signal tristate
flabel metal2 s 213192 -960 213416 480 0 FreeSans 896 90 0 0 la_data_in[0]
port 114 nsew signal input
flabel metal2 s 270312 -960 270536 480 0 FreeSans 896 90 0 0 la_data_in[10]
port 115 nsew signal input
flabel metal2 s 276024 -960 276248 480 0 FreeSans 896 90 0 0 la_data_in[11]
port 116 nsew signal input
flabel metal2 s 281736 -960 281960 480 0 FreeSans 896 90 0 0 la_data_in[12]
port 117 nsew signal input
flabel metal2 s 287448 -960 287672 480 0 FreeSans 896 90 0 0 la_data_in[13]
port 118 nsew signal input
flabel metal2 s 293160 -960 293384 480 0 FreeSans 896 90 0 0 la_data_in[14]
port 119 nsew signal input
flabel metal2 s 298872 -960 299096 480 0 FreeSans 896 90 0 0 la_data_in[15]
port 120 nsew signal input
flabel metal2 s 304584 -960 304808 480 0 FreeSans 896 90 0 0 la_data_in[16]
port 121 nsew signal input
flabel metal2 s 310296 -960 310520 480 0 FreeSans 896 90 0 0 la_data_in[17]
port 122 nsew signal input
flabel metal2 s 316008 -960 316232 480 0 FreeSans 896 90 0 0 la_data_in[18]
port 123 nsew signal input
flabel metal2 s 321720 -960 321944 480 0 FreeSans 896 90 0 0 la_data_in[19]
port 124 nsew signal input
flabel metal2 s 218904 -960 219128 480 0 FreeSans 896 90 0 0 la_data_in[1]
port 125 nsew signal input
flabel metal2 s 327432 -960 327656 480 0 FreeSans 896 90 0 0 la_data_in[20]
port 126 nsew signal input
flabel metal2 s 333144 -960 333368 480 0 FreeSans 896 90 0 0 la_data_in[21]
port 127 nsew signal input
flabel metal2 s 338856 -960 339080 480 0 FreeSans 896 90 0 0 la_data_in[22]
port 128 nsew signal input
flabel metal2 s 344568 -960 344792 480 0 FreeSans 896 90 0 0 la_data_in[23]
port 129 nsew signal input
flabel metal2 s 350280 -960 350504 480 0 FreeSans 896 90 0 0 la_data_in[24]
port 130 nsew signal input
flabel metal2 s 355992 -960 356216 480 0 FreeSans 896 90 0 0 la_data_in[25]
port 131 nsew signal input
flabel metal2 s 361704 -960 361928 480 0 FreeSans 896 90 0 0 la_data_in[26]
port 132 nsew signal input
flabel metal2 s 367416 -960 367640 480 0 FreeSans 896 90 0 0 la_data_in[27]
port 133 nsew signal input
flabel metal2 s 373128 -960 373352 480 0 FreeSans 896 90 0 0 la_data_in[28]
port 134 nsew signal input
flabel metal2 s 378840 -960 379064 480 0 FreeSans 896 90 0 0 la_data_in[29]
port 135 nsew signal input
flabel metal2 s 224616 -960 224840 480 0 FreeSans 896 90 0 0 la_data_in[2]
port 136 nsew signal input
flabel metal2 s 384552 -960 384776 480 0 FreeSans 896 90 0 0 la_data_in[30]
port 137 nsew signal input
flabel metal2 s 390264 -960 390488 480 0 FreeSans 896 90 0 0 la_data_in[31]
port 138 nsew signal input
flabel metal2 s 395976 -960 396200 480 0 FreeSans 896 90 0 0 la_data_in[32]
port 139 nsew signal input
flabel metal2 s 401688 -960 401912 480 0 FreeSans 896 90 0 0 la_data_in[33]
port 140 nsew signal input
flabel metal2 s 407400 -960 407624 480 0 FreeSans 896 90 0 0 la_data_in[34]
port 141 nsew signal input
flabel metal2 s 413112 -960 413336 480 0 FreeSans 896 90 0 0 la_data_in[35]
port 142 nsew signal input
flabel metal2 s 418824 -960 419048 480 0 FreeSans 896 90 0 0 la_data_in[36]
port 143 nsew signal input
flabel metal2 s 424536 -960 424760 480 0 FreeSans 896 90 0 0 la_data_in[37]
port 144 nsew signal input
flabel metal2 s 430248 -960 430472 480 0 FreeSans 896 90 0 0 la_data_in[38]
port 145 nsew signal input
flabel metal2 s 435960 -960 436184 480 0 FreeSans 896 90 0 0 la_data_in[39]
port 146 nsew signal input
flabel metal2 s 230328 -960 230552 480 0 FreeSans 896 90 0 0 la_data_in[3]
port 147 nsew signal input
flabel metal2 s 441672 -960 441896 480 0 FreeSans 896 90 0 0 la_data_in[40]
port 148 nsew signal input
flabel metal2 s 447384 -960 447608 480 0 FreeSans 896 90 0 0 la_data_in[41]
port 149 nsew signal input
flabel metal2 s 453096 -960 453320 480 0 FreeSans 896 90 0 0 la_data_in[42]
port 150 nsew signal input
flabel metal2 s 458808 -960 459032 480 0 FreeSans 896 90 0 0 la_data_in[43]
port 151 nsew signal input
flabel metal2 s 464520 -960 464744 480 0 FreeSans 896 90 0 0 la_data_in[44]
port 152 nsew signal input
flabel metal2 s 470232 -960 470456 480 0 FreeSans 896 90 0 0 la_data_in[45]
port 153 nsew signal input
flabel metal2 s 475944 -960 476168 480 0 FreeSans 896 90 0 0 la_data_in[46]
port 154 nsew signal input
flabel metal2 s 481656 -960 481880 480 0 FreeSans 896 90 0 0 la_data_in[47]
port 155 nsew signal input
flabel metal2 s 487368 -960 487592 480 0 FreeSans 896 90 0 0 la_data_in[48]
port 156 nsew signal input
flabel metal2 s 493080 -960 493304 480 0 FreeSans 896 90 0 0 la_data_in[49]
port 157 nsew signal input
flabel metal2 s 236040 -960 236264 480 0 FreeSans 896 90 0 0 la_data_in[4]
port 158 nsew signal input
flabel metal2 s 498792 -960 499016 480 0 FreeSans 896 90 0 0 la_data_in[50]
port 159 nsew signal input
flabel metal2 s 504504 -960 504728 480 0 FreeSans 896 90 0 0 la_data_in[51]
port 160 nsew signal input
flabel metal2 s 510216 -960 510440 480 0 FreeSans 896 90 0 0 la_data_in[52]
port 161 nsew signal input
flabel metal2 s 515928 -960 516152 480 0 FreeSans 896 90 0 0 la_data_in[53]
port 162 nsew signal input
flabel metal2 s 521640 -960 521864 480 0 FreeSans 896 90 0 0 la_data_in[54]
port 163 nsew signal input
flabel metal2 s 527352 -960 527576 480 0 FreeSans 896 90 0 0 la_data_in[55]
port 164 nsew signal input
flabel metal2 s 533064 -960 533288 480 0 FreeSans 896 90 0 0 la_data_in[56]
port 165 nsew signal input
flabel metal2 s 538776 -960 539000 480 0 FreeSans 896 90 0 0 la_data_in[57]
port 166 nsew signal input
flabel metal2 s 544488 -960 544712 480 0 FreeSans 896 90 0 0 la_data_in[58]
port 167 nsew signal input
flabel metal2 s 550200 -960 550424 480 0 FreeSans 896 90 0 0 la_data_in[59]
port 168 nsew signal input
flabel metal2 s 241752 -960 241976 480 0 FreeSans 896 90 0 0 la_data_in[5]
port 169 nsew signal input
flabel metal2 s 555912 -960 556136 480 0 FreeSans 896 90 0 0 la_data_in[60]
port 170 nsew signal input
flabel metal2 s 561624 -960 561848 480 0 FreeSans 896 90 0 0 la_data_in[61]
port 171 nsew signal input
flabel metal2 s 567336 -960 567560 480 0 FreeSans 896 90 0 0 la_data_in[62]
port 172 nsew signal input
flabel metal2 s 573048 -960 573272 480 0 FreeSans 896 90 0 0 la_data_in[63]
port 173 nsew signal input
flabel metal2 s 247464 -960 247688 480 0 FreeSans 896 90 0 0 la_data_in[6]
port 174 nsew signal input
flabel metal2 s 253176 -960 253400 480 0 FreeSans 896 90 0 0 la_data_in[7]
port 175 nsew signal input
flabel metal2 s 258888 -960 259112 480 0 FreeSans 896 90 0 0 la_data_in[8]
port 176 nsew signal input
flabel metal2 s 264600 -960 264824 480 0 FreeSans 896 90 0 0 la_data_in[9]
port 177 nsew signal input
flabel metal2 s 215096 -960 215320 480 0 FreeSans 896 90 0 0 la_data_out[0]
port 178 nsew signal tristate
flabel metal2 s 272216 -960 272440 480 0 FreeSans 896 90 0 0 la_data_out[10]
port 179 nsew signal tristate
flabel metal2 s 277928 -960 278152 480 0 FreeSans 896 90 0 0 la_data_out[11]
port 180 nsew signal tristate
flabel metal2 s 283640 -960 283864 480 0 FreeSans 896 90 0 0 la_data_out[12]
port 181 nsew signal tristate
flabel metal2 s 289352 -960 289576 480 0 FreeSans 896 90 0 0 la_data_out[13]
port 182 nsew signal tristate
flabel metal2 s 295064 -960 295288 480 0 FreeSans 896 90 0 0 la_data_out[14]
port 183 nsew signal tristate
flabel metal2 s 300776 -960 301000 480 0 FreeSans 896 90 0 0 la_data_out[15]
port 184 nsew signal tristate
flabel metal2 s 306488 -960 306712 480 0 FreeSans 896 90 0 0 la_data_out[16]
port 185 nsew signal tristate
flabel metal2 s 312200 -960 312424 480 0 FreeSans 896 90 0 0 la_data_out[17]
port 186 nsew signal tristate
flabel metal2 s 317912 -960 318136 480 0 FreeSans 896 90 0 0 la_data_out[18]
port 187 nsew signal tristate
flabel metal2 s 323624 -960 323848 480 0 FreeSans 896 90 0 0 la_data_out[19]
port 188 nsew signal tristate
flabel metal2 s 220808 -960 221032 480 0 FreeSans 896 90 0 0 la_data_out[1]
port 189 nsew signal tristate
flabel metal2 s 329336 -960 329560 480 0 FreeSans 896 90 0 0 la_data_out[20]
port 190 nsew signal tristate
flabel metal2 s 335048 -960 335272 480 0 FreeSans 896 90 0 0 la_data_out[21]
port 191 nsew signal tristate
flabel metal2 s 340760 -960 340984 480 0 FreeSans 896 90 0 0 la_data_out[22]
port 192 nsew signal tristate
flabel metal2 s 346472 -960 346696 480 0 FreeSans 896 90 0 0 la_data_out[23]
port 193 nsew signal tristate
flabel metal2 s 352184 -960 352408 480 0 FreeSans 896 90 0 0 la_data_out[24]
port 194 nsew signal tristate
flabel metal2 s 357896 -960 358120 480 0 FreeSans 896 90 0 0 la_data_out[25]
port 195 nsew signal tristate
flabel metal2 s 363608 -960 363832 480 0 FreeSans 896 90 0 0 la_data_out[26]
port 196 nsew signal tristate
flabel metal2 s 369320 -960 369544 480 0 FreeSans 896 90 0 0 la_data_out[27]
port 197 nsew signal tristate
flabel metal2 s 375032 -960 375256 480 0 FreeSans 896 90 0 0 la_data_out[28]
port 198 nsew signal tristate
flabel metal2 s 380744 -960 380968 480 0 FreeSans 896 90 0 0 la_data_out[29]
port 199 nsew signal tristate
flabel metal2 s 226520 -960 226744 480 0 FreeSans 896 90 0 0 la_data_out[2]
port 200 nsew signal tristate
flabel metal2 s 386456 -960 386680 480 0 FreeSans 896 90 0 0 la_data_out[30]
port 201 nsew signal tristate
flabel metal2 s 392168 -960 392392 480 0 FreeSans 896 90 0 0 la_data_out[31]
port 202 nsew signal tristate
flabel metal2 s 397880 -960 398104 480 0 FreeSans 896 90 0 0 la_data_out[32]
port 203 nsew signal tristate
flabel metal2 s 403592 -960 403816 480 0 FreeSans 896 90 0 0 la_data_out[33]
port 204 nsew signal tristate
flabel metal2 s 409304 -960 409528 480 0 FreeSans 896 90 0 0 la_data_out[34]
port 205 nsew signal tristate
flabel metal2 s 415016 -960 415240 480 0 FreeSans 896 90 0 0 la_data_out[35]
port 206 nsew signal tristate
flabel metal2 s 420728 -960 420952 480 0 FreeSans 896 90 0 0 la_data_out[36]
port 207 nsew signal tristate
flabel metal2 s 426440 -960 426664 480 0 FreeSans 896 90 0 0 la_data_out[37]
port 208 nsew signal tristate
flabel metal2 s 432152 -960 432376 480 0 FreeSans 896 90 0 0 la_data_out[38]
port 209 nsew signal tristate
flabel metal2 s 437864 -960 438088 480 0 FreeSans 896 90 0 0 la_data_out[39]
port 210 nsew signal tristate
flabel metal2 s 232232 -960 232456 480 0 FreeSans 896 90 0 0 la_data_out[3]
port 211 nsew signal tristate
flabel metal2 s 443576 -960 443800 480 0 FreeSans 896 90 0 0 la_data_out[40]
port 212 nsew signal tristate
flabel metal2 s 449288 -960 449512 480 0 FreeSans 896 90 0 0 la_data_out[41]
port 213 nsew signal tristate
flabel metal2 s 455000 -960 455224 480 0 FreeSans 896 90 0 0 la_data_out[42]
port 214 nsew signal tristate
flabel metal2 s 460712 -960 460936 480 0 FreeSans 896 90 0 0 la_data_out[43]
port 215 nsew signal tristate
flabel metal2 s 466424 -960 466648 480 0 FreeSans 896 90 0 0 la_data_out[44]
port 216 nsew signal tristate
flabel metal2 s 472136 -960 472360 480 0 FreeSans 896 90 0 0 la_data_out[45]
port 217 nsew signal tristate
flabel metal2 s 477848 -960 478072 480 0 FreeSans 896 90 0 0 la_data_out[46]
port 218 nsew signal tristate
flabel metal2 s 483560 -960 483784 480 0 FreeSans 896 90 0 0 la_data_out[47]
port 219 nsew signal tristate
flabel metal2 s 489272 -960 489496 480 0 FreeSans 896 90 0 0 la_data_out[48]
port 220 nsew signal tristate
flabel metal2 s 494984 -960 495208 480 0 FreeSans 896 90 0 0 la_data_out[49]
port 221 nsew signal tristate
flabel metal2 s 237944 -960 238168 480 0 FreeSans 896 90 0 0 la_data_out[4]
port 222 nsew signal tristate
flabel metal2 s 500696 -960 500920 480 0 FreeSans 896 90 0 0 la_data_out[50]
port 223 nsew signal tristate
flabel metal2 s 506408 -960 506632 480 0 FreeSans 896 90 0 0 la_data_out[51]
port 224 nsew signal tristate
flabel metal2 s 512120 -960 512344 480 0 FreeSans 896 90 0 0 la_data_out[52]
port 225 nsew signal tristate
flabel metal2 s 517832 -960 518056 480 0 FreeSans 896 90 0 0 la_data_out[53]
port 226 nsew signal tristate
flabel metal2 s 523544 -960 523768 480 0 FreeSans 896 90 0 0 la_data_out[54]
port 227 nsew signal tristate
flabel metal2 s 529256 -960 529480 480 0 FreeSans 896 90 0 0 la_data_out[55]
port 228 nsew signal tristate
flabel metal2 s 534968 -960 535192 480 0 FreeSans 896 90 0 0 la_data_out[56]
port 229 nsew signal tristate
flabel metal2 s 540680 -960 540904 480 0 FreeSans 896 90 0 0 la_data_out[57]
port 230 nsew signal tristate
flabel metal2 s 546392 -960 546616 480 0 FreeSans 896 90 0 0 la_data_out[58]
port 231 nsew signal tristate
flabel metal2 s 552104 -960 552328 480 0 FreeSans 896 90 0 0 la_data_out[59]
port 232 nsew signal tristate
flabel metal2 s 243656 -960 243880 480 0 FreeSans 896 90 0 0 la_data_out[5]
port 233 nsew signal tristate
flabel metal2 s 557816 -960 558040 480 0 FreeSans 896 90 0 0 la_data_out[60]
port 234 nsew signal tristate
flabel metal2 s 563528 -960 563752 480 0 FreeSans 896 90 0 0 la_data_out[61]
port 235 nsew signal tristate
flabel metal2 s 569240 -960 569464 480 0 FreeSans 896 90 0 0 la_data_out[62]
port 236 nsew signal tristate
flabel metal2 s 574952 -960 575176 480 0 FreeSans 896 90 0 0 la_data_out[63]
port 237 nsew signal tristate
flabel metal2 s 249368 -960 249592 480 0 FreeSans 896 90 0 0 la_data_out[6]
port 238 nsew signal tristate
flabel metal2 s 255080 -960 255304 480 0 FreeSans 896 90 0 0 la_data_out[7]
port 239 nsew signal tristate
flabel metal2 s 260792 -960 261016 480 0 FreeSans 896 90 0 0 la_data_out[8]
port 240 nsew signal tristate
flabel metal2 s 266504 -960 266728 480 0 FreeSans 896 90 0 0 la_data_out[9]
port 241 nsew signal tristate
flabel metal2 s 217000 -960 217224 480 0 FreeSans 896 90 0 0 la_oenb[0]
port 242 nsew signal input
flabel metal2 s 274120 -960 274344 480 0 FreeSans 896 90 0 0 la_oenb[10]
port 243 nsew signal input
flabel metal2 s 279832 -960 280056 480 0 FreeSans 896 90 0 0 la_oenb[11]
port 244 nsew signal input
flabel metal2 s 285544 -960 285768 480 0 FreeSans 896 90 0 0 la_oenb[12]
port 245 nsew signal input
flabel metal2 s 291256 -960 291480 480 0 FreeSans 896 90 0 0 la_oenb[13]
port 246 nsew signal input
flabel metal2 s 296968 -960 297192 480 0 FreeSans 896 90 0 0 la_oenb[14]
port 247 nsew signal input
flabel metal2 s 302680 -960 302904 480 0 FreeSans 896 90 0 0 la_oenb[15]
port 248 nsew signal input
flabel metal2 s 308392 -960 308616 480 0 FreeSans 896 90 0 0 la_oenb[16]
port 249 nsew signal input
flabel metal2 s 314104 -960 314328 480 0 FreeSans 896 90 0 0 la_oenb[17]
port 250 nsew signal input
flabel metal2 s 319816 -960 320040 480 0 FreeSans 896 90 0 0 la_oenb[18]
port 251 nsew signal input
flabel metal2 s 325528 -960 325752 480 0 FreeSans 896 90 0 0 la_oenb[19]
port 252 nsew signal input
flabel metal2 s 222712 -960 222936 480 0 FreeSans 896 90 0 0 la_oenb[1]
port 253 nsew signal input
flabel metal2 s 331240 -960 331464 480 0 FreeSans 896 90 0 0 la_oenb[20]
port 254 nsew signal input
flabel metal2 s 336952 -960 337176 480 0 FreeSans 896 90 0 0 la_oenb[21]
port 255 nsew signal input
flabel metal2 s 342664 -960 342888 480 0 FreeSans 896 90 0 0 la_oenb[22]
port 256 nsew signal input
flabel metal2 s 348376 -960 348600 480 0 FreeSans 896 90 0 0 la_oenb[23]
port 257 nsew signal input
flabel metal2 s 354088 -960 354312 480 0 FreeSans 896 90 0 0 la_oenb[24]
port 258 nsew signal input
flabel metal2 s 359800 -960 360024 480 0 FreeSans 896 90 0 0 la_oenb[25]
port 259 nsew signal input
flabel metal2 s 365512 -960 365736 480 0 FreeSans 896 90 0 0 la_oenb[26]
port 260 nsew signal input
flabel metal2 s 371224 -960 371448 480 0 FreeSans 896 90 0 0 la_oenb[27]
port 261 nsew signal input
flabel metal2 s 376936 -960 377160 480 0 FreeSans 896 90 0 0 la_oenb[28]
port 262 nsew signal input
flabel metal2 s 382648 -960 382872 480 0 FreeSans 896 90 0 0 la_oenb[29]
port 263 nsew signal input
flabel metal2 s 228424 -960 228648 480 0 FreeSans 896 90 0 0 la_oenb[2]
port 264 nsew signal input
flabel metal2 s 388360 -960 388584 480 0 FreeSans 896 90 0 0 la_oenb[30]
port 265 nsew signal input
flabel metal2 s 394072 -960 394296 480 0 FreeSans 896 90 0 0 la_oenb[31]
port 266 nsew signal input
flabel metal2 s 399784 -960 400008 480 0 FreeSans 896 90 0 0 la_oenb[32]
port 267 nsew signal input
flabel metal2 s 405496 -960 405720 480 0 FreeSans 896 90 0 0 la_oenb[33]
port 268 nsew signal input
flabel metal2 s 411208 -960 411432 480 0 FreeSans 896 90 0 0 la_oenb[34]
port 269 nsew signal input
flabel metal2 s 416920 -960 417144 480 0 FreeSans 896 90 0 0 la_oenb[35]
port 270 nsew signal input
flabel metal2 s 422632 -960 422856 480 0 FreeSans 896 90 0 0 la_oenb[36]
port 271 nsew signal input
flabel metal2 s 428344 -960 428568 480 0 FreeSans 896 90 0 0 la_oenb[37]
port 272 nsew signal input
flabel metal2 s 434056 -960 434280 480 0 FreeSans 896 90 0 0 la_oenb[38]
port 273 nsew signal input
flabel metal2 s 439768 -960 439992 480 0 FreeSans 896 90 0 0 la_oenb[39]
port 274 nsew signal input
flabel metal2 s 234136 -960 234360 480 0 FreeSans 896 90 0 0 la_oenb[3]
port 275 nsew signal input
flabel metal2 s 445480 -960 445704 480 0 FreeSans 896 90 0 0 la_oenb[40]
port 276 nsew signal input
flabel metal2 s 451192 -960 451416 480 0 FreeSans 896 90 0 0 la_oenb[41]
port 277 nsew signal input
flabel metal2 s 456904 -960 457128 480 0 FreeSans 896 90 0 0 la_oenb[42]
port 278 nsew signal input
flabel metal2 s 462616 -960 462840 480 0 FreeSans 896 90 0 0 la_oenb[43]
port 279 nsew signal input
flabel metal2 s 468328 -960 468552 480 0 FreeSans 896 90 0 0 la_oenb[44]
port 280 nsew signal input
flabel metal2 s 474040 -960 474264 480 0 FreeSans 896 90 0 0 la_oenb[45]
port 281 nsew signal input
flabel metal2 s 479752 -960 479976 480 0 FreeSans 896 90 0 0 la_oenb[46]
port 282 nsew signal input
flabel metal2 s 485464 -960 485688 480 0 FreeSans 896 90 0 0 la_oenb[47]
port 283 nsew signal input
flabel metal2 s 491176 -960 491400 480 0 FreeSans 896 90 0 0 la_oenb[48]
port 284 nsew signal input
flabel metal2 s 496888 -960 497112 480 0 FreeSans 896 90 0 0 la_oenb[49]
port 285 nsew signal input
flabel metal2 s 239848 -960 240072 480 0 FreeSans 896 90 0 0 la_oenb[4]
port 286 nsew signal input
flabel metal2 s 502600 -960 502824 480 0 FreeSans 896 90 0 0 la_oenb[50]
port 287 nsew signal input
flabel metal2 s 508312 -960 508536 480 0 FreeSans 896 90 0 0 la_oenb[51]
port 288 nsew signal input
flabel metal2 s 514024 -960 514248 480 0 FreeSans 896 90 0 0 la_oenb[52]
port 289 nsew signal input
flabel metal2 s 519736 -960 519960 480 0 FreeSans 896 90 0 0 la_oenb[53]
port 290 nsew signal input
flabel metal2 s 525448 -960 525672 480 0 FreeSans 896 90 0 0 la_oenb[54]
port 291 nsew signal input
flabel metal2 s 531160 -960 531384 480 0 FreeSans 896 90 0 0 la_oenb[55]
port 292 nsew signal input
flabel metal2 s 536872 -960 537096 480 0 FreeSans 896 90 0 0 la_oenb[56]
port 293 nsew signal input
flabel metal2 s 542584 -960 542808 480 0 FreeSans 896 90 0 0 la_oenb[57]
port 294 nsew signal input
flabel metal2 s 548296 -960 548520 480 0 FreeSans 896 90 0 0 la_oenb[58]
port 295 nsew signal input
flabel metal2 s 554008 -960 554232 480 0 FreeSans 896 90 0 0 la_oenb[59]
port 296 nsew signal input
flabel metal2 s 245560 -960 245784 480 0 FreeSans 896 90 0 0 la_oenb[5]
port 297 nsew signal input
flabel metal2 s 559720 -960 559944 480 0 FreeSans 896 90 0 0 la_oenb[60]
port 298 nsew signal input
flabel metal2 s 565432 -960 565656 480 0 FreeSans 896 90 0 0 la_oenb[61]
port 299 nsew signal input
flabel metal2 s 571144 -960 571368 480 0 FreeSans 896 90 0 0 la_oenb[62]
port 300 nsew signal input
flabel metal2 s 576856 -960 577080 480 0 FreeSans 896 90 0 0 la_oenb[63]
port 301 nsew signal input
flabel metal2 s 251272 -960 251496 480 0 FreeSans 896 90 0 0 la_oenb[6]
port 302 nsew signal input
flabel metal2 s 256984 -960 257208 480 0 FreeSans 896 90 0 0 la_oenb[7]
port 303 nsew signal input
flabel metal2 s 262696 -960 262920 480 0 FreeSans 896 90 0 0 la_oenb[8]
port 304 nsew signal input
flabel metal2 s 268408 -960 268632 480 0 FreeSans 896 90 0 0 la_oenb[9]
port 305 nsew signal input
flabel metal2 s 578760 -960 578984 480 0 FreeSans 896 90 0 0 user_clock2
port 306 nsew signal input
flabel metal2 s 580664 -960 580888 480 0 FreeSans 896 90 0 0 user_irq[0]
port 307 nsew signal tristate
flabel metal2 s 582568 -960 582792 480 0 FreeSans 896 90 0 0 user_irq[1]
port 308 nsew signal tristate
flabel metal2 s 584472 -960 584696 480 0 FreeSans 896 90 0 0 user_irq[2]
port 309 nsew signal tristate
flabel metal4 s -956 -684 -336 597308 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -956 -684 597020 -64 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -956 596688 597020 597308 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 596400 -684 597020 597308 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 5418 -1644 6038 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 36138 -1644 36758 114770 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 36138 129486 36758 256610 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 36138 267966 36758 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 66858 -1644 67478 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 97578 -1644 98198 44578 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 97578 50558 98198 399122 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 97578 406894 98198 473234 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 97578 480894 98198 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 128298 -1644 128918 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 159018 -1644 159638 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 189738 -1644 190358 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 220458 -1644 221078 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 251178 -1644 251798 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 281898 -1644 282518 68098 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 281898 567214 282518 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 312618 -1644 313238 68098 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 312618 567214 313238 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 343338 -1644 343958 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 374058 -1644 374678 115218 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 374058 121870 374678 399570 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 374058 404318 374678 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 404778 -1644 405398 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 435498 -1644 436118 45698 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 435498 53694 436118 114322 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 435498 119854 436118 404498 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 435498 409918 436118 472114 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 435498 478094 436118 540962 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 435498 551870 436118 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 466218 -1644 466838 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 496938 -1644 497558 115106 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 496938 125454 497558 262994 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 496938 268414 497558 330274 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 496938 338718 497558 470322 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 496938 476414 497558 551602 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 496938 557694 497558 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 527658 -1644 528278 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 558378 -1644 558998 42338 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 558378 52910 558998 468754 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 558378 482014 558998 545554 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 558378 550974 558998 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s 589098 -1644 589718 598268 0 FreeSans 2560 90 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 3826 597980 4446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 21826 597980 22446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 39826 597980 40446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 57826 597980 58446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 75826 597980 76446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 93826 597980 94446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 111826 597980 112446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 129826 597980 130446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 147826 597980 148446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 165826 597980 166446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 183826 597980 184446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 201826 597980 202446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 219826 597980 220446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 237826 597980 238446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 255826 597980 256446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 273826 597980 274446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 291826 597980 292446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 309826 597980 310446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 327826 597980 328446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 345826 597980 346446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 363826 597980 364446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 381826 597980 382446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 399826 597980 400446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 417826 597980 418446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 435826 597980 436446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 453826 597980 454446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 471826 597980 472446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 489826 597980 490446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 507826 597980 508446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 525826 597980 526446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 543826 597980 544446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 561826 597980 562446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal5 s -1916 579826 597980 580446 0 FreeSans 4608 0 0 0 vdd
port 310 nsew power bidirectional
flabel metal4 s -1916 -1644 -1296 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 -1644 597980 -1024 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 597648 597980 598268 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 597360 -1644 597980 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 9138 -1644 9758 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 39858 -1644 40478 30164 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 39858 69788 40478 101364 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 39858 140988 40478 172564 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 39858 568188 40478 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 70578 -1644 71198 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 101298 -1644 101918 30164 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 101298 69788 101918 101364 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 101298 140988 101918 172564 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 101298 568188 101918 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 132018 -1644 132638 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 162738 -1644 163358 48274 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 162738 53358 163358 120034 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 162738 125678 163358 184626 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 162738 193966 163358 262098 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 162738 266958 163358 329602 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 162738 342190 163358 542754 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 162738 553886 163358 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 193458 -1644 194078 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 224178 -1644 224798 473122 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 224178 483918 224798 543986 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 224178 551870 224798 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 254898 -1644 255518 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 285618 -1644 286238 68098 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 285618 567214 286238 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 316338 -1644 316958 68098 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 316338 567214 316958 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 347058 -1644 347678 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 377778 -1644 378398 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 408498 -1644 409118 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 439218 -1644 439838 404498 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 439218 409918 439838 540962 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 439218 551870 439838 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 469938 -1644 470558 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 500658 -1644 501278 262994 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 500658 268414 501278 403714 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 500658 409246 501278 551602 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 500658 557694 501278 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 531378 -1644 531998 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 562098 -1644 562718 332178 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 562098 338830 562718 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal4 s 592818 -1644 593438 598268 0 FreeSans 2560 90 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 9826 597980 10446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 27826 597980 28446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 45826 597980 46446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 63826 597980 64446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 81826 597980 82446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 99826 597980 100446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 117826 597980 118446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 135826 597980 136446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 153826 597980 154446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 171826 597980 172446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 189826 597980 190446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 207826 597980 208446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 225826 597980 226446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 243826 597980 244446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 261826 597980 262446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 279826 597980 280446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 297826 597980 298446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 315826 597980 316446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 333826 597980 334446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 351826 597980 352446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 369826 597980 370446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 387826 597980 388446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 405826 597980 406446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 423826 597980 424446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 441826 597980 442446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 459826 597980 460446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 477826 597980 478446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 495826 597980 496446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 513826 597980 514446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 531826 597980 532446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 549826 597980 550446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 567826 597980 568446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal5 s -1916 585826 597980 586446 0 FreeSans 4608 0 0 0 vss
port 311 nsew ground bidirectional
flabel metal2 s 11368 -960 11592 480 0 FreeSans 896 90 0 0 wb_clk_i
port 312 nsew signal input
flabel metal2 s 13272 -960 13496 480 0 FreeSans 896 90 0 0 wb_rst_i
port 313 nsew signal input
flabel metal2 s 15176 -960 15400 480 0 FreeSans 896 90 0 0 wbs_ack_o
port 314 nsew signal tristate
flabel metal2 s 22792 -960 23016 480 0 FreeSans 896 90 0 0 wbs_adr_i[0]
port 315 nsew signal input
flabel metal2 s 87528 -960 87752 480 0 FreeSans 896 90 0 0 wbs_adr_i[10]
port 316 nsew signal input
flabel metal2 s 93240 -960 93464 480 0 FreeSans 896 90 0 0 wbs_adr_i[11]
port 317 nsew signal input
flabel metal2 s 98952 -960 99176 480 0 FreeSans 896 90 0 0 wbs_adr_i[12]
port 318 nsew signal input
flabel metal2 s 104664 -960 104888 480 0 FreeSans 896 90 0 0 wbs_adr_i[13]
port 319 nsew signal input
flabel metal2 s 110376 -960 110600 480 0 FreeSans 896 90 0 0 wbs_adr_i[14]
port 320 nsew signal input
flabel metal2 s 116088 -960 116312 480 0 FreeSans 896 90 0 0 wbs_adr_i[15]
port 321 nsew signal input
flabel metal2 s 121800 -960 122024 480 0 FreeSans 896 90 0 0 wbs_adr_i[16]
port 322 nsew signal input
flabel metal2 s 127512 -960 127736 480 0 FreeSans 896 90 0 0 wbs_adr_i[17]
port 323 nsew signal input
flabel metal2 s 133224 -960 133448 480 0 FreeSans 896 90 0 0 wbs_adr_i[18]
port 324 nsew signal input
flabel metal2 s 138936 -960 139160 480 0 FreeSans 896 90 0 0 wbs_adr_i[19]
port 325 nsew signal input
flabel metal2 s 30408 -960 30632 480 0 FreeSans 896 90 0 0 wbs_adr_i[1]
port 326 nsew signal input
flabel metal2 s 144648 -960 144872 480 0 FreeSans 896 90 0 0 wbs_adr_i[20]
port 327 nsew signal input
flabel metal2 s 150360 -960 150584 480 0 FreeSans 896 90 0 0 wbs_adr_i[21]
port 328 nsew signal input
flabel metal2 s 156072 -960 156296 480 0 FreeSans 896 90 0 0 wbs_adr_i[22]
port 329 nsew signal input
flabel metal2 s 161784 -960 162008 480 0 FreeSans 896 90 0 0 wbs_adr_i[23]
port 330 nsew signal input
flabel metal2 s 167496 -960 167720 480 0 FreeSans 896 90 0 0 wbs_adr_i[24]
port 331 nsew signal input
flabel metal2 s 173208 -960 173432 480 0 FreeSans 896 90 0 0 wbs_adr_i[25]
port 332 nsew signal input
flabel metal2 s 178920 -960 179144 480 0 FreeSans 896 90 0 0 wbs_adr_i[26]
port 333 nsew signal input
flabel metal2 s 184632 -960 184856 480 0 FreeSans 896 90 0 0 wbs_adr_i[27]
port 334 nsew signal input
flabel metal2 s 190344 -960 190568 480 0 FreeSans 896 90 0 0 wbs_adr_i[28]
port 335 nsew signal input
flabel metal2 s 196056 -960 196280 480 0 FreeSans 896 90 0 0 wbs_adr_i[29]
port 336 nsew signal input
flabel metal2 s 38024 -960 38248 480 0 FreeSans 896 90 0 0 wbs_adr_i[2]
port 337 nsew signal input
flabel metal2 s 201768 -960 201992 480 0 FreeSans 896 90 0 0 wbs_adr_i[30]
port 338 nsew signal input
flabel metal2 s 207480 -960 207704 480 0 FreeSans 896 90 0 0 wbs_adr_i[31]
port 339 nsew signal input
flabel metal2 s 45640 -960 45864 480 0 FreeSans 896 90 0 0 wbs_adr_i[3]
port 340 nsew signal input
flabel metal2 s 53256 -960 53480 480 0 FreeSans 896 90 0 0 wbs_adr_i[4]
port 341 nsew signal input
flabel metal2 s 58968 -960 59192 480 0 FreeSans 896 90 0 0 wbs_adr_i[5]
port 342 nsew signal input
flabel metal2 s 64680 -960 64904 480 0 FreeSans 896 90 0 0 wbs_adr_i[6]
port 343 nsew signal input
flabel metal2 s 70392 -960 70616 480 0 FreeSans 896 90 0 0 wbs_adr_i[7]
port 344 nsew signal input
flabel metal2 s 76104 -960 76328 480 0 FreeSans 896 90 0 0 wbs_adr_i[8]
port 345 nsew signal input
flabel metal2 s 81816 -960 82040 480 0 FreeSans 896 90 0 0 wbs_adr_i[9]
port 346 nsew signal input
flabel metal2 s 17080 -960 17304 480 0 FreeSans 896 90 0 0 wbs_cyc_i
port 347 nsew signal input
flabel metal2 s 24696 -960 24920 480 0 FreeSans 896 90 0 0 wbs_dat_i[0]
port 348 nsew signal input
flabel metal2 s 89432 -960 89656 480 0 FreeSans 896 90 0 0 wbs_dat_i[10]
port 349 nsew signal input
flabel metal2 s 95144 -960 95368 480 0 FreeSans 896 90 0 0 wbs_dat_i[11]
port 350 nsew signal input
flabel metal2 s 100856 -960 101080 480 0 FreeSans 896 90 0 0 wbs_dat_i[12]
port 351 nsew signal input
flabel metal2 s 106568 -960 106792 480 0 FreeSans 896 90 0 0 wbs_dat_i[13]
port 352 nsew signal input
flabel metal2 s 112280 -960 112504 480 0 FreeSans 896 90 0 0 wbs_dat_i[14]
port 353 nsew signal input
flabel metal2 s 117992 -960 118216 480 0 FreeSans 896 90 0 0 wbs_dat_i[15]
port 354 nsew signal input
flabel metal2 s 123704 -960 123928 480 0 FreeSans 896 90 0 0 wbs_dat_i[16]
port 355 nsew signal input
flabel metal2 s 129416 -960 129640 480 0 FreeSans 896 90 0 0 wbs_dat_i[17]
port 356 nsew signal input
flabel metal2 s 135128 -960 135352 480 0 FreeSans 896 90 0 0 wbs_dat_i[18]
port 357 nsew signal input
flabel metal2 s 140840 -960 141064 480 0 FreeSans 896 90 0 0 wbs_dat_i[19]
port 358 nsew signal input
flabel metal2 s 32312 -960 32536 480 0 FreeSans 896 90 0 0 wbs_dat_i[1]
port 359 nsew signal input
flabel metal2 s 146552 -960 146776 480 0 FreeSans 896 90 0 0 wbs_dat_i[20]
port 360 nsew signal input
flabel metal2 s 152264 -960 152488 480 0 FreeSans 896 90 0 0 wbs_dat_i[21]
port 361 nsew signal input
flabel metal2 s 157976 -960 158200 480 0 FreeSans 896 90 0 0 wbs_dat_i[22]
port 362 nsew signal input
flabel metal2 s 163688 -960 163912 480 0 FreeSans 896 90 0 0 wbs_dat_i[23]
port 363 nsew signal input
flabel metal2 s 169400 -960 169624 480 0 FreeSans 896 90 0 0 wbs_dat_i[24]
port 364 nsew signal input
flabel metal2 s 175112 -960 175336 480 0 FreeSans 896 90 0 0 wbs_dat_i[25]
port 365 nsew signal input
flabel metal2 s 180824 -960 181048 480 0 FreeSans 896 90 0 0 wbs_dat_i[26]
port 366 nsew signal input
flabel metal2 s 186536 -960 186760 480 0 FreeSans 896 90 0 0 wbs_dat_i[27]
port 367 nsew signal input
flabel metal2 s 192248 -960 192472 480 0 FreeSans 896 90 0 0 wbs_dat_i[28]
port 368 nsew signal input
flabel metal2 s 197960 -960 198184 480 0 FreeSans 896 90 0 0 wbs_dat_i[29]
port 369 nsew signal input
flabel metal2 s 39928 -960 40152 480 0 FreeSans 896 90 0 0 wbs_dat_i[2]
port 370 nsew signal input
flabel metal2 s 203672 -960 203896 480 0 FreeSans 896 90 0 0 wbs_dat_i[30]
port 371 nsew signal input
flabel metal2 s 209384 -960 209608 480 0 FreeSans 896 90 0 0 wbs_dat_i[31]
port 372 nsew signal input
flabel metal2 s 47544 -960 47768 480 0 FreeSans 896 90 0 0 wbs_dat_i[3]
port 373 nsew signal input
flabel metal2 s 55160 -960 55384 480 0 FreeSans 896 90 0 0 wbs_dat_i[4]
port 374 nsew signal input
flabel metal2 s 60872 -960 61096 480 0 FreeSans 896 90 0 0 wbs_dat_i[5]
port 375 nsew signal input
flabel metal2 s 66584 -960 66808 480 0 FreeSans 896 90 0 0 wbs_dat_i[6]
port 376 nsew signal input
flabel metal2 s 72296 -960 72520 480 0 FreeSans 896 90 0 0 wbs_dat_i[7]
port 377 nsew signal input
flabel metal2 s 78008 -960 78232 480 0 FreeSans 896 90 0 0 wbs_dat_i[8]
port 378 nsew signal input
flabel metal2 s 83720 -960 83944 480 0 FreeSans 896 90 0 0 wbs_dat_i[9]
port 379 nsew signal input
flabel metal2 s 26600 -960 26824 480 0 FreeSans 896 90 0 0 wbs_dat_o[0]
port 380 nsew signal tristate
flabel metal2 s 91336 -960 91560 480 0 FreeSans 896 90 0 0 wbs_dat_o[10]
port 381 nsew signal tristate
flabel metal2 s 97048 -960 97272 480 0 FreeSans 896 90 0 0 wbs_dat_o[11]
port 382 nsew signal tristate
flabel metal2 s 102760 -960 102984 480 0 FreeSans 896 90 0 0 wbs_dat_o[12]
port 383 nsew signal tristate
flabel metal2 s 108472 -960 108696 480 0 FreeSans 896 90 0 0 wbs_dat_o[13]
port 384 nsew signal tristate
flabel metal2 s 114184 -960 114408 480 0 FreeSans 896 90 0 0 wbs_dat_o[14]
port 385 nsew signal tristate
flabel metal2 s 119896 -960 120120 480 0 FreeSans 896 90 0 0 wbs_dat_o[15]
port 386 nsew signal tristate
flabel metal2 s 125608 -960 125832 480 0 FreeSans 896 90 0 0 wbs_dat_o[16]
port 387 nsew signal tristate
flabel metal2 s 131320 -960 131544 480 0 FreeSans 896 90 0 0 wbs_dat_o[17]
port 388 nsew signal tristate
flabel metal2 s 137032 -960 137256 480 0 FreeSans 896 90 0 0 wbs_dat_o[18]
port 389 nsew signal tristate
flabel metal2 s 142744 -960 142968 480 0 FreeSans 896 90 0 0 wbs_dat_o[19]
port 390 nsew signal tristate
flabel metal2 s 34216 -960 34440 480 0 FreeSans 896 90 0 0 wbs_dat_o[1]
port 391 nsew signal tristate
flabel metal2 s 148456 -960 148680 480 0 FreeSans 896 90 0 0 wbs_dat_o[20]
port 392 nsew signal tristate
flabel metal2 s 154168 -960 154392 480 0 FreeSans 896 90 0 0 wbs_dat_o[21]
port 393 nsew signal tristate
flabel metal2 s 159880 -960 160104 480 0 FreeSans 896 90 0 0 wbs_dat_o[22]
port 394 nsew signal tristate
flabel metal2 s 165592 -960 165816 480 0 FreeSans 896 90 0 0 wbs_dat_o[23]
port 395 nsew signal tristate
flabel metal2 s 171304 -960 171528 480 0 FreeSans 896 90 0 0 wbs_dat_o[24]
port 396 nsew signal tristate
flabel metal2 s 177016 -960 177240 480 0 FreeSans 896 90 0 0 wbs_dat_o[25]
port 397 nsew signal tristate
flabel metal2 s 182728 -960 182952 480 0 FreeSans 896 90 0 0 wbs_dat_o[26]
port 398 nsew signal tristate
flabel metal2 s 188440 -960 188664 480 0 FreeSans 896 90 0 0 wbs_dat_o[27]
port 399 nsew signal tristate
flabel metal2 s 194152 -960 194376 480 0 FreeSans 896 90 0 0 wbs_dat_o[28]
port 400 nsew signal tristate
flabel metal2 s 199864 -960 200088 480 0 FreeSans 896 90 0 0 wbs_dat_o[29]
port 401 nsew signal tristate
flabel metal2 s 41832 -960 42056 480 0 FreeSans 896 90 0 0 wbs_dat_o[2]
port 402 nsew signal tristate
flabel metal2 s 205576 -960 205800 480 0 FreeSans 896 90 0 0 wbs_dat_o[30]
port 403 nsew signal tristate
flabel metal2 s 211288 -960 211512 480 0 FreeSans 896 90 0 0 wbs_dat_o[31]
port 404 nsew signal tristate
flabel metal2 s 49448 -960 49672 480 0 FreeSans 896 90 0 0 wbs_dat_o[3]
port 405 nsew signal tristate
flabel metal2 s 57064 -960 57288 480 0 FreeSans 896 90 0 0 wbs_dat_o[4]
port 406 nsew signal tristate
flabel metal2 s 62776 -960 63000 480 0 FreeSans 896 90 0 0 wbs_dat_o[5]
port 407 nsew signal tristate
flabel metal2 s 68488 -960 68712 480 0 FreeSans 896 90 0 0 wbs_dat_o[6]
port 408 nsew signal tristate
flabel metal2 s 74200 -960 74424 480 0 FreeSans 896 90 0 0 wbs_dat_o[7]
port 409 nsew signal tristate
flabel metal2 s 79912 -960 80136 480 0 FreeSans 896 90 0 0 wbs_dat_o[8]
port 410 nsew signal tristate
flabel metal2 s 85624 -960 85848 480 0 FreeSans 896 90 0 0 wbs_dat_o[9]
port 411 nsew signal tristate
flabel metal2 s 28504 -960 28728 480 0 FreeSans 896 90 0 0 wbs_sel_i[0]
port 412 nsew signal input
flabel metal2 s 36120 -960 36344 480 0 FreeSans 896 90 0 0 wbs_sel_i[1]
port 413 nsew signal input
flabel metal2 s 43736 -960 43960 480 0 FreeSans 896 90 0 0 wbs_sel_i[2]
port 414 nsew signal input
flabel metal2 s 51352 -960 51576 480 0 FreeSans 896 90 0 0 wbs_sel_i[3]
port 415 nsew signal input
flabel metal2 s 18984 -960 19208 480 0 FreeSans 896 90 0 0 wbs_stb_i
port 416 nsew signal input
flabel metal2 s 20888 -960 21112 480 0 FreeSans 896 90 0 0 wbs_we_i
port 417 nsew signal input
rlabel via4 55390 130322 55390 130322 0 vdd
rlabel via4 40354 100322 40354 100322 0 vss
rlabel metal2 273672 570038 273672 570038 0 io_in[10]
rlabel metal2 274792 569870 274792 569870 0 io_in[11]
rlabel metal2 269192 569814 269192 569814 0 io_in[6]
rlabel metal4 270312 568344 270312 568344 0 io_in[7]
rlabel metal3 591458 324520 591458 324520 0 io_in[8]
rlabel metal4 272552 568232 272552 568232 0 io_in[9]
rlabel metal4 289352 567907 289352 567907 0 io_oeb[0]
rlabel metal2 400680 498904 400680 498904 0 io_oeb[10]
rlabel metal3 590562 469896 590562 469896 0 io_oeb[11]
rlabel metal3 302792 568624 302792 568624 0 io_oeb[12]
rlabel metal4 303688 568512 303688 568512 0 io_oeb[13]
rlabel metal2 305032 579054 305032 579054 0 io_oeb[14]
rlabel metal2 306152 571662 306152 571662 0 io_oeb[15]
rlabel metal2 307272 576646 307272 576646 0 io_oeb[16]
rlabel metal2 308392 573342 308392 573342 0 io_oeb[17]
rlabel metal2 309512 574182 309512 574182 0 io_oeb[18]
rlabel metal2 310632 571774 310632 571774 0 io_oeb[19]
rlabel metal2 290472 569646 290472 569646 0 io_oeb[1]
rlabel metal2 209608 588938 209608 588938 0 io_oeb[20]
rlabel metal2 143416 584794 143416 584794 0 io_oeb[21]
rlabel metal2 77336 584682 77336 584682 0 io_oeb[22]
rlabel metal2 11032 587202 11032 587202 0 io_oeb[23]
rlabel metal3 2310 559160 2310 559160 0 io_oeb[24]
rlabel metal3 134302 516600 134302 516600 0 io_oeb[25]
rlabel metal3 2478 474488 2478 474488 0 io_oeb[26]
rlabel metal2 266392 500304 266392 500304 0 io_oeb[27]
rlabel metal3 168336 569128 168336 569128 0 io_oeb[28]
rlabel metal3 4046 347480 4046 347480 0 io_oeb[29]
rlabel metal3 591402 113064 591402 113064 0 io_oeb[2]
rlabel metal2 266616 437192 266616 437192 0 io_oeb[30]
rlabel metal3 2422 262808 2422 262808 0 io_oeb[31]
rlabel metal3 2366 220472 2366 220472 0 io_oeb[32]
rlabel metal2 326312 570486 326312 570486 0 io_oeb[33]
rlabel metal2 327432 570598 327432 570598 0 io_oeb[34]
rlabel metal2 328552 570934 328552 570934 0 io_oeb[35]
rlabel metal3 2310 51128 2310 51128 0 io_oeb[36]
rlabel metal2 330792 570374 330792 570374 0 io_oeb[37]
rlabel metal2 292712 569926 292712 569926 0 io_oeb[3]
rlabel metal2 293832 569646 293832 569646 0 io_oeb[4]
rlabel metal2 294952 569982 294952 569982 0 io_oeb[5]
rlabel metal2 296072 569702 296072 569702 0 io_oeb[6]
rlabel metal2 474600 440384 474600 440384 0 io_oeb[7]
rlabel metal3 593082 350952 593082 350952 0 io_oeb[8]
rlabel metal3 593138 390600 593138 390600 0 io_oeb[9]
rlabel metal3 593194 496328 593194 496328 0 io_out[12]
rlabel metal3 593138 535864 593138 535864 0 io_out[13]
rlabel metal2 278152 572446 278152 572446 0 io_out[14]
rlabel metal2 562632 593082 562632 593082 0 io_out[15]
rlabel metal2 496440 593082 496440 593082 0 io_out[16]
rlabel metal2 430248 593082 430248 593082 0 io_out[17]
rlabel metal3 285376 574392 285376 574392 0 io_out[18]
rlabel metal3 286776 576184 286776 576184 0 io_out[19]
rlabel metal2 284872 573342 284872 573342 0 io_out[20]
rlabel metal2 165704 593138 165704 593138 0 io_out[21]
rlabel metal2 99512 593082 99512 593082 0 io_out[22]
rlabel metal2 46200 587160 46200 587160 0 io_out[23]
rlabel metal2 76440 301392 76440 301392 0 io_out[24]
rlabel metal3 145600 29624 145600 29624 0 io_out[25]
rlabel metal3 148568 29512 148568 29512 0 io_out[26]
rlabel metal2 287112 28826 287112 28826 0 io_out[27]
rlabel metal3 3990 403704 3990 403704 0 io_out[28]
rlabel metal2 266392 195216 266392 195216 0 io_out[29]
rlabel metal2 299880 28882 299880 28882 0 io_out[30]
rlabel metal2 304136 29162 304136 29162 0 io_out[31]
rlabel metal2 308392 28770 308392 28770 0 io_out[32]
rlabel metal3 2534 192024 2534 192024 0 io_out[33]
rlabel metal3 2422 149688 2422 149688 0 io_out[34]
rlabel metal2 265496 28896 265496 28896 0 io_out[35]
rlabel metal3 2422 65016 2422 65016 0 io_out[36]
rlabel metal3 2310 22904 2310 22904 0 io_out[37]
rlabel metal2 50344 79646 50344 79646 0 itasegm1\[0\]
rlabel metal3 337078 117768 337078 117768 0 itasegm1\[100\]
rlabel metal3 335342 118328 335342 118328 0 itasegm1\[101\]
rlabel metal3 338646 118888 338646 118888 0 itasegm1\[102\]
rlabel metal3 340326 119448 340326 119448 0 itasegm1\[103\]
rlabel metal3 334446 120008 334446 120008 0 itasegm1\[104\]
rlabel metal3 336910 120568 336910 120568 0 itasegm1\[105\]
rlabel metal4 350280 96320 350280 96320 0 itasegm1\[106\]
rlabel metal4 351848 117964 351848 117964 0 itasegm1\[107\]
rlabel metal3 334502 122248 334502 122248 0 itasegm1\[108\]
rlabel metal4 352296 100520 352296 100520 0 itasegm1\[109\]
rlabel metal4 263816 95200 263816 95200 0 itasegm1\[10\]
rlabel metal3 334390 123368 334390 123368 0 itasegm1\[110\]
rlabel metal3 338646 123928 338646 123928 0 itasegm1\[111\]
rlabel metal4 263816 150920 263816 150920 0 itasegm1\[112\]
rlabel metal2 38920 99666 38920 99666 0 itasegm1\[113\]
rlabel metal2 42280 147406 42280 147406 0 itasegm1\[114\]
rlabel metal4 69720 135800 69720 135800 0 itasegm1\[115\]
rlabel metal2 73080 125496 73080 125496 0 itasegm1\[116\]
rlabel metal3 88928 100968 88928 100968 0 itasegm1\[117\]
rlabel metal3 63294 117880 63294 117880 0 itasegm1\[118\]
rlabel metal2 74760 128464 74760 128464 0 itasegm1\[119\]
rlabel metal4 74760 69664 74760 69664 0 itasegm1\[11\]
rlabel metal2 69720 128352 69720 128352 0 itasegm1\[120\]
rlabel metal3 19138 121240 19138 121240 0 itasegm1\[121\]
rlabel metal3 63350 121912 63350 121912 0 itasegm1\[122\]
rlabel metal3 63462 121240 63462 121240 0 itasegm1\[123\]
rlabel metal3 63560 101080 63560 101080 0 itasegm1\[124\]
rlabel metal3 63406 126616 63406 126616 0 itasegm1\[125\]
rlabel metal2 88088 150766 88088 150766 0 itasegm1\[126\]
rlabel metal3 125510 119896 125510 119896 0 itasegm1\[127\]
rlabel metal2 125272 129528 125272 129528 0 itasegm1\[128\]
rlabel metal3 125734 136696 125734 136696 0 itasegm1\[129\]
rlabel metal4 69832 67312 69832 67312 0 itasegm1\[12\]
rlabel metal3 125398 119224 125398 119224 0 itasegm1\[130\]
rlabel metal2 104216 99666 104216 99666 0 itasegm1\[131\]
rlabel metal3 197666 162568 197666 162568 0 itasegm1\[132\]
rlabel metal3 125678 125944 125678 125944 0 itasegm1\[133\]
rlabel metal3 125454 122584 125454 122584 0 itasegm1\[134\]
rlabel metal3 125566 121912 125566 121912 0 itasegm1\[135\]
rlabel metal2 263032 132832 263032 132832 0 itasegm1\[136\]
rlabel metal2 261576 157976 261576 157976 0 itasegm1\[137\]
rlabel metal3 118552 100632 118552 100632 0 itasegm1\[138\]
rlabel metal2 125160 134064 125160 134064 0 itasegm1\[139\]
rlabel metal2 42952 27986 42952 27986 0 itasegm1\[13\]
rlabel metal3 233562 167048 233562 167048 0 itasegm1\[140\]
rlabel metal3 185864 118902 185864 118902 0 itasegm1\[141\]
rlabel metal3 190806 125944 190806 125944 0 itasegm1\[142\]
rlabel metal3 189126 125272 189126 125272 0 itasegm1\[143\]
rlabel metal2 168952 99666 168952 99666 0 itasegm1\[144\]
rlabel metal3 187446 124600 187446 124600 0 itasegm1\[145\]
rlabel metal2 187320 135576 187320 135576 0 itasegm1\[146\]
rlabel metal2 166264 99610 166264 99610 0 itasegm1\[147\]
rlabel metal2 263816 171024 263816 171024 0 itasegm1\[148\]
rlabel metal2 161560 144718 161560 144718 0 itasegm1\[149\]
rlabel metal2 89432 27874 89432 27874 0 itasegm1\[14\]
rlabel metal2 162904 146510 162904 146510 0 itasegm1\[150\]
rlabel metal2 164248 144774 164248 144774 0 itasegm1\[151\]
rlabel metal3 142450 124600 142450 124600 0 itasegm1\[152\]
rlabel metal2 168350 142296 168350 142296 0 itasegm1\[153\]
rlabel metal2 256312 167664 256312 167664 0 itasegm1\[154\]
rlabel metal3 241248 100744 241248 100744 0 itasegm1\[155\]
rlabel metal4 263816 175000 263816 175000 0 itasegm1\[156\]
rlabel metal2 257992 167664 257992 167664 0 itasegm1\[157\]
rlabel metal3 242200 100632 242200 100632 0 itasegm1\[158\]
rlabel metal4 264712 174944 264712 174944 0 itasegm1\[159\]
rlabel metal3 123928 56238 123928 56238 0 itasegm1\[15\]
rlabel metal3 252182 121912 252182 121912 0 itasegm1\[160\]
rlabel metal3 252910 126616 252910 126616 0 itasegm1\[161\]
rlabel metal4 262920 146944 262920 146944 0 itasegm1\[162\]
rlabel metal3 250390 125272 250390 125272 0 itasegm1\[163\]
rlabel metal4 230216 101248 230216 101248 0 itasegm1\[164\]
rlabel metal2 259784 169064 259784 169064 0 itasegm1\[165\]
rlabel metal4 264600 155064 264600 155064 0 itasegm1\[166\]
rlabel metal3 247912 117278 247912 117278 0 itasegm1\[167\]
rlabel metal4 396536 143360 396536 143360 0 itasegm1\[168\]
rlabel metal4 368872 101248 368872 101248 0 itasegm1\[169\]
rlabel metal3 267736 101136 267736 101136 0 itasegm1\[16\]
rlabel metal2 374248 144718 374248 144718 0 itasegm1\[170\]
rlabel metal2 376936 147238 376936 147238 0 itasegm1\[171\]
rlabel metal4 368200 101304 368200 101304 0 itasegm1\[172\]
rlabel metal3 333998 154168 333998 154168 0 itasegm1\[173\]
rlabel metal4 396984 129248 396984 129248 0 itasegm1\[174\]
rlabel metal4 397096 124880 397096 124880 0 itasegm1\[175\]
rlabel metal4 357224 149800 357224 149800 0 itasegm1\[176\]
rlabel metal3 349930 120568 349930 120568 0 itasegm1\[177\]
rlabel metal3 393960 118902 393960 118902 0 itasegm1\[178\]
rlabel metal4 396760 133336 396760 133336 0 itasegm1\[179\]
rlabel metal2 100856 72982 100856 72982 0 itasegm1\[17\]
rlabel metal4 396536 118328 396536 118328 0 itasegm1\[180\]
rlabel metal4 352072 149744 352072 149744 0 itasegm1\[181\]
rlabel metal4 422072 101360 422072 101360 0 itasegm1\[182\]
rlabel metal2 428792 100394 428792 100394 0 itasegm1\[183\]
rlabel metal3 457478 118552 457478 118552 0 itasegm1\[184\]
rlabel metal2 407400 130872 407400 130872 0 itasegm1\[185\]
rlabel metal4 429464 101304 429464 101304 0 itasegm1\[186\]
rlabel metal3 456022 119224 456022 119224 0 itasegm1\[187\]
rlabel metal3 457310 117208 457310 117208 0 itasegm1\[188\]
rlabel metal4 452760 152600 452760 152600 0 itasegm1\[189\]
rlabel metal4 141960 71568 141960 71568 0 itasegm1\[18\]
rlabel metal3 371350 163688 371350 163688 0 itasegm1\[190\]
rlabel metal2 399000 133000 399000 133000 0 itasegm1\[191\]
rlabel metal3 335286 164808 335286 164808 0 itasegm1\[192\]
rlabel metal3 393638 165368 393638 165368 0 itasegm1\[193\]
rlabel metal3 373030 165928 373030 165928 0 itasegm1\[194\]
rlabel metal4 357000 161056 357000 161056 0 itasegm1\[195\]
rlabel metal2 494200 150598 494200 150598 0 itasegm1\[196\]
rlabel metal3 518574 115864 518574 115864 0 itasegm1\[197\]
rlabel metal3 334446 168168 334446 168168 0 itasegm1\[198\]
rlabel metal3 333214 168728 333214 168728 0 itasegm1\[199\]
rlabel metal4 138600 83104 138600 83104 0 itasegm1\[19\]
rlabel metal3 247394 93688 247394 93688 0 itasegm1\[1\]
rlabel metal3 519470 117208 519470 117208 0 itasegm1\[200\]
rlabel metal2 472920 135352 472920 135352 0 itasegm1\[201\]
rlabel metal3 468706 119896 468706 119896 0 itasegm1\[202\]
rlabel metal4 380520 161560 380520 161560 0 itasegm1\[203\]
rlabel metal3 333998 171528 333998 171528 0 itasegm1\[204\]
rlabel metal3 519526 119896 519526 119896 0 itasegm1\[205\]
rlabel metal3 474474 117208 474474 117208 0 itasegm1\[206\]
rlabel metal4 517496 149912 517496 149912 0 itasegm1\[207\]
rlabel metal4 472136 119000 472136 119000 0 itasegm1\[208\]
rlabel metal2 474600 137480 474600 137480 0 itasegm1\[209\]
rlabel metal4 263928 102984 263928 102984 0 itasegm1\[20\]
rlabel metal4 351960 165144 351960 165144 0 itasegm1\[210\]
rlabel metal3 462448 163800 462448 163800 0 itasegm1\[211\]
rlabel metal3 581574 124600 581574 124600 0 itasegm1\[212\]
rlabel metal3 333214 176568 333214 176568 0 itasegm1\[213\]
rlabel metal4 350280 159544 350280 159544 0 itasegm1\[214\]
rlabel metal3 333662 177688 333662 177688 0 itasegm1\[215\]
rlabel metal3 449400 162120 449400 162120 0 itasegm1\[216\]
rlabel metal2 351960 165424 351960 165424 0 itasegm1\[217\]
rlabel metal3 333662 179368 333662 179368 0 itasegm1\[218\]
rlabel metal3 581630 122584 581630 122584 0 itasegm1\[219\]
rlabel metal4 263816 104104 263816 104104 0 itasegm1\[21\]
rlabel metal2 564312 99778 564312 99778 0 itasegm1\[220\]
rlabel metal3 536578 117208 536578 117208 0 itasegm1\[221\]
rlabel metal2 558936 99722 558936 99722 0 itasegm1\[222\]
rlabel metal3 336182 182168 336182 182168 0 itasegm1\[223\]
rlabel metal4 263816 210000 263816 210000 0 itasegm1\[224\]
rlabel metal2 46662 213528 46662 213528 0 itasegm1\[225\]
rlabel metal3 61768 194614 61768 194614 0 itasegm1\[226\]
rlabel metal2 125160 190344 125160 190344 0 itasegm1\[227\]
rlabel metal2 44968 214326 44968 214326 0 itasegm1\[228\]
rlabel metal2 259672 190960 259672 190960 0 itasegm1\[229\]
rlabel metal2 258216 98616 258216 98616 0 itasegm1\[22\]
rlabel metal2 69720 192136 69720 192136 0 itasegm1\[230\]
rlabel metal4 263816 212800 263816 212800 0 itasegm1\[231\]
rlabel metal3 63294 187096 63294 187096 0 itasegm1\[232\]
rlabel metal4 74760 201544 74760 201544 0 itasegm1\[233\]
rlabel metal2 264712 194544 264712 194544 0 itasegm1\[234\]
rlabel metal4 263928 214536 263928 214536 0 itasegm1\[235\]
rlabel metal4 263816 215264 263816 215264 0 itasegm1\[236\]
rlabel metal2 44968 171472 44968 171472 0 itasegm1\[237\]
rlabel metal2 104216 215502 104216 215502 0 itasegm1\[238\]
rlabel metal2 106232 215782 106232 215782 0 itasegm1\[239\]
rlabel metal3 125454 54152 125454 54152 0 itasegm1\[23\]
rlabel metal4 263816 218064 263816 218064 0 itasegm1\[240\]
rlabel metal2 102200 216342 102200 216342 0 itasegm1\[241\]
rlabel metal2 105560 216622 105560 216622 0 itasegm1\[242\]
rlabel metal4 263816 219744 263816 219744 0 itasegm1\[243\]
rlabel metal3 81130 193816 81130 193816 0 itasegm1\[244\]
rlabel metal3 81018 194488 81018 194488 0 itasegm1\[245\]
rlabel metal3 125454 192472 125454 192472 0 itasegm1\[246\]
rlabel metal3 81242 195160 81242 195160 0 itasegm1\[247\]
rlabel metal3 81074 190456 81074 190456 0 itasegm1\[248\]
rlabel metal3 125398 189112 125398 189112 0 itasegm1\[249\]
rlabel metal2 256424 96600 256424 96600 0 itasegm1\[24\]
rlabel metal2 100184 171402 100184 171402 0 itasegm1\[250\]
rlabel metal3 81186 197848 81186 197848 0 itasegm1\[251\]
rlabel metal4 144088 216440 144088 216440 0 itasegm1\[252\]
rlabel metal3 189126 193816 189126 193816 0 itasegm1\[253\]
rlabel metal3 191646 197176 191646 197176 0 itasegm1\[254\]
rlabel metal3 213458 226968 213458 226968 0 itasegm1\[255\]
rlabel metal3 187446 193144 187446 193144 0 itasegm1\[256\]
rlabel metal3 187558 195160 187558 195160 0 itasegm1\[257\]
rlabel metal3 215810 228648 215810 228648 0 itasegm1\[258\]
rlabel metal3 217154 229208 217154 229208 0 itasegm1\[259\]
rlabel metal4 259784 95984 259784 95984 0 itasegm1\[25\]
rlabel metal3 142506 188440 142506 188440 0 itasegm1\[260\]
rlabel metal3 142450 192472 142450 192472 0 itasegm1\[261\]
rlabel metal2 166936 171458 166936 171458 0 itasegm1\[262\]
rlabel metal3 142394 198520 142394 198520 0 itasegm1\[263\]
rlabel metal3 182000 171752 182000 171752 0 itasegm1\[264\]
rlabel metal3 142338 187768 142338 187768 0 itasegm1\[265\]
rlabel metal3 246778 233128 246778 233128 0 itasegm1\[266\]
rlabel metal3 260904 233464 260904 233464 0 itasegm1\[267\]
rlabel metal4 256200 213024 256200 213024 0 itasegm1\[268\]
rlabel metal4 261240 220360 261240 220360 0 itasegm1\[269\]
rlabel metal2 98840 74606 98840 74606 0 itasegm1\[26\]
rlabel metal3 263368 235144 263368 235144 0 itasegm1\[270\]
rlabel metal4 264936 225904 264936 225904 0 itasegm1\[271\]
rlabel metal3 204666 187096 204666 187096 0 itasegm1\[272\]
rlabel metal2 259560 204176 259560 204176 0 itasegm1\[273\]
rlabel metal2 261240 204680 261240 204680 0 itasegm1\[274\]
rlabel metal2 262920 204680 262920 204680 0 itasegm1\[275\]
rlabel metal3 260904 235368 260904 235368 0 itasegm1\[276\]
rlabel metal4 263816 237664 263816 237664 0 itasegm1\[277\]
rlabel metal3 204610 187768 204610 187768 0 itasegm1\[278\]
rlabel metal2 263816 239904 263816 239904 0 itasegm1\[279\]
rlabel metal3 263984 105336 263984 105336 0 itasegm1\[27\]
rlabel metal2 339304 211624 339304 211624 0 itasegm1\[280\]
rlabel metal3 346178 192472 346178 192472 0 itasegm1\[281\]
rlabel metal4 396872 199584 396872 199584 0 itasegm1\[282\]
rlabel metal4 396536 199556 396536 199556 0 itasegm1\[283\]
rlabel metal3 345282 191128 345282 191128 0 itasegm1\[284\]
rlabel metal3 331912 212478 331912 212478 0 itasegm1\[285\]
rlabel metal3 331912 212898 331912 212898 0 itasegm1\[286\]
rlabel metal3 346122 194488 346122 194488 0 itasegm1\[287\]
rlabel metal3 346346 195832 346346 195832 0 itasegm1\[288\]
rlabel metal3 346234 195160 346234 195160 0 itasegm1\[289\]
rlabel metal4 265160 103544 265160 103544 0 itasegm1\[28\]
rlabel metal3 334502 215208 334502 215208 0 itasegm1\[290\]
rlabel metal3 334390 215768 334390 215768 0 itasegm1\[291\]
rlabel metal3 333998 216328 333998 216328 0 itasegm1\[292\]
rlabel metal2 372904 215222 372904 215222 0 itasegm1\[293\]
rlabel metal2 436184 215502 436184 215502 0 itasegm1\[294\]
rlabel metal4 356216 216216 356216 216216 0 itasegm1\[295\]
rlabel metal3 372190 218568 372190 218568 0 itasegm1\[296\]
rlabel metal4 339304 216160 339304 216160 0 itasegm1\[297\]
rlabel metal4 407400 205408 407400 205408 0 itasegm1\[298\]
rlabel metal2 399000 195720 399000 195720 0 itasegm1\[299\]
rlabel metal3 190806 55496 190806 55496 0 itasegm1\[29\]
rlabel metal2 263816 93800 263816 93800 0 itasegm1\[2\]
rlabel metal3 333942 220808 333942 220808 0 itasegm1\[300\]
rlabel metal4 351960 216272 351960 216272 0 itasegm1\[301\]
rlabel metal2 429240 219856 429240 219856 0 itasegm1\[302\]
rlabel metal3 455336 196546 455336 196546 0 itasegm1\[303\]
rlabel metal2 406616 221200 406616 221200 0 itasegm1\[304\]
rlabel metal3 457422 191800 457422 191800 0 itasegm1\[305\]
rlabel metal3 423136 171640 423136 171640 0 itasegm1\[306\]
rlabel metal2 427560 221424 427560 221424 0 itasegm1\[307\]
rlabel metal4 472136 211400 472136 211400 0 itasegm1\[308\]
rlabel metal2 496216 171402 496216 171402 0 itasegm1\[309\]
rlabel metal3 187670 65576 187670 65576 0 itasegm1\[30\]
rlabel metal2 495544 171346 495544 171346 0 itasegm1\[310\]
rlabel metal3 518126 176344 518126 176344 0 itasegm1\[311\]
rlabel metal2 494872 171234 494872 171234 0 itasegm1\[312\]
rlabel metal3 519582 181720 519582 181720 0 itasegm1\[313\]
rlabel metal3 517944 196070 517944 196070 0 itasegm1\[314\]
rlabel metal3 519470 196504 519470 196504 0 itasegm1\[315\]
rlabel metal3 518966 193144 518966 193144 0 itasegm1\[316\]
rlabel metal2 501592 215670 501592 215670 0 itasegm1\[317\]
rlabel metal2 494200 171290 494200 171290 0 itasegm1\[318\]
rlabel metal3 517944 190806 517944 190806 0 itasegm1\[319\]
rlabel metal2 165592 80598 165592 80598 0 itasegm1\[31\]
rlabel metal3 519526 192472 519526 192472 0 itasegm1\[320\]
rlabel metal2 500920 215614 500920 215614 0 itasegm1\[321\]
rlabel metal2 350280 227864 350280 227864 0 itasegm1\[322\]
rlabel metal3 581686 189784 581686 189784 0 itasegm1\[323\]
rlabel metal3 395710 234248 395710 234248 0 itasegm1\[324\]
rlabel metal2 571704 171472 571704 171472 0 itasegm1\[325\]
rlabel metal3 580622 189112 580622 189112 0 itasegm1\[326\]
rlabel metal2 562296 215110 562296 215110 0 itasegm1\[327\]
rlabel metal4 400680 223720 400680 223720 0 itasegm1\[328\]
rlabel metal3 333550 237048 333550 237048 0 itasegm1\[329\]
rlabel metal2 162904 75446 162904 75446 0 itasegm1\[32\]
rlabel metal3 335230 237608 335230 237608 0 itasegm1\[330\]
rlabel metal3 333214 238168 333214 238168 0 itasegm1\[331\]
rlabel metal3 333830 238728 333830 238728 0 itasegm1\[332\]
rlabel metal3 333158 239288 333158 239288 0 itasegm1\[333\]
rlabel metal3 333942 239848 333942 239848 0 itasegm1\[334\]
rlabel metal3 417550 240408 417550 240408 0 itasegm1\[335\]
rlabel metal4 124376 272070 124376 272070 0 itasegm1\[336\]
rlabel metal2 264936 276304 264936 276304 0 itasegm1\[337\]
rlabel metal3 258440 285768 258440 285768 0 itasegm1\[338\]
rlabel metal4 263816 269179 263816 269179 0 itasegm1\[339\]
rlabel metal3 143402 65576 143402 65576 0 itasegm1\[33\]
rlabel metal2 26824 241514 26824 241514 0 itasegm1\[340\]
rlabel metal2 143640 285376 143640 285376 0 itasegm1\[341\]
rlabel metal2 167160 241304 167160 241304 0 itasegm1\[342\]
rlabel metal4 263928 271289 263928 271289 0 itasegm1\[343\]
rlabel metal4 194936 270810 194936 270810 0 itasegm1\[344\]
rlabel metal4 262136 271579 262136 271579 0 itasegm1\[345\]
rlabel metal2 44296 242354 44296 242354 0 itasegm1\[346\]
rlabel metal3 260064 273784 260064 273784 0 itasegm1\[347\]
rlabel metal2 262920 257040 262920 257040 0 itasegm1\[348\]
rlabel metal3 63070 267736 63070 267736 0 itasegm1\[349\]
rlabel metal2 169624 27818 169624 27818 0 itasegm1\[34\]
rlabel metal4 262248 274329 262248 274329 0 itasegm1\[350\]
rlabel metal3 176232 284536 176232 284536 0 itasegm1\[351\]
rlabel metal4 263816 276239 263816 276239 0 itasegm1\[352\]
rlabel metal4 262136 276879 262136 276879 0 itasegm1\[353\]
rlabel metal2 102200 285334 102200 285334 0 itasegm1\[354\]
rlabel metal2 257992 260680 257992 260680 0 itasegm1\[355\]
rlabel metal4 263368 278529 263368 278529 0 itasegm1\[356\]
rlabel metal4 195720 272610 195720 272610 0 itasegm1\[357\]
rlabel metal2 258664 283920 258664 283920 0 itasegm1\[358\]
rlabel metal3 255360 281288 255360 281288 0 itasegm1\[359\]
rlabel metal2 167608 27762 167608 27762 0 itasegm1\[35\]
rlabel metal3 127134 266392 127134 266392 0 itasegm1\[360\]
rlabel metal3 130438 264376 130438 264376 0 itasegm1\[361\]
rlabel metal3 81186 263032 81186 263032 0 itasegm1\[362\]
rlabel metal4 138600 271656 138600 271656 0 itasegm1\[363\]
rlabel metal3 195006 263032 195006 263032 0 itasegm1\[364\]
rlabel metal4 261240 284648 261240 284648 0 itasegm1\[365\]
rlabel metal3 263144 284704 263144 284704 0 itasegm1\[366\]
rlabel metal2 162232 241234 162232 241234 0 itasegm1\[367\]
rlabel metal3 143402 261016 143402 261016 0 itasegm1\[368\]
rlabel metal2 168952 285558 168952 285558 0 itasegm1\[369\]
rlabel metal3 187502 49448 187502 49448 0 itasegm1\[36\]
rlabel metal2 170646 284760 170646 284760 0 itasegm1\[370\]
rlabel metal2 169624 286118 169624 286118 0 itasegm1\[371\]
rlabel metal3 193326 260344 193326 260344 0 itasegm1\[372\]
rlabel metal2 165592 241066 165592 241066 0 itasegm1\[373\]
rlabel metal3 187446 259000 187446 259000 0 itasegm1\[374\]
rlabel metal2 170296 241514 170296 241514 0 itasegm1\[375\]
rlabel metal3 187558 263704 187558 263704 0 itasegm1\[376\]
rlabel metal3 142506 265048 142506 265048 0 itasegm1\[377\]
rlabel metal3 205506 266392 205506 266392 0 itasegm1\[378\]
rlabel metal2 232904 288358 232904 288358 0 itasegm1\[379\]
rlabel metal3 187614 54824 187614 54824 0 itasegm1\[37\]
rlabel metal3 250390 258328 250390 258328 0 itasegm1\[380\]
rlabel metal4 206136 279048 206136 279048 0 itasegm1\[381\]
rlabel metal3 205450 279160 205450 279160 0 itasegm1\[382\]
rlabel metal2 224168 289478 224168 289478 0 itasegm1\[383\]
rlabel metal3 204610 267064 204610 267064 0 itasegm1\[384\]
rlabel metal2 224840 290038 224840 290038 0 itasegm1\[385\]
rlabel metal3 204554 264376 204554 264376 0 itasegm1\[386\]
rlabel metal2 228872 290598 228872 290598 0 itasegm1\[387\]
rlabel metal2 257880 268296 257880 268296 0 itasegm1\[388\]
rlabel metal2 263816 297080 263816 297080 0 itasegm1\[389\]
rlabel metal3 187446 54152 187446 54152 0 itasegm1\[38\]
rlabel metal2 263928 296464 263928 296464 0 itasegm1\[390\]
rlabel metal3 262080 285656 262080 285656 0 itasegm1\[391\]
rlabel metal2 368872 285222 368872 285222 0 itasegm1\[392\]
rlabel metal3 333158 268408 333158 268408 0 itasegm1\[393\]
rlabel metal3 333830 268968 333830 268968 0 itasegm1\[394\]
rlabel metal2 352184 276976 352184 276976 0 itasegm1\[395\]
rlabel metal3 333214 270088 333214 270088 0 itasegm1\[396\]
rlabel metal2 375592 285390 375592 285390 0 itasegm1\[397\]
rlabel metal2 375592 242074 375592 242074 0 itasegm1\[398\]
rlabel metal3 356720 243320 356720 243320 0 itasegm1\[399\]
rlabel metal2 168280 79758 168280 79758 0 itasegm1\[39\]
rlabel metal2 38920 27874 38920 27874 0 itasegm1\[3\]
rlabel metal3 333214 272328 333214 272328 0 itasegm1\[400\]
rlabel metal4 351064 272299 351064 272299 0 itasegm1\[401\]
rlabel metal3 333158 273448 333158 273448 0 itasegm1\[402\]
rlabel metal3 333214 274008 333214 274008 0 itasegm1\[403\]
rlabel metal3 333270 274568 333270 274568 0 itasegm1\[404\]
rlabel metal3 334446 275128 334446 275128 0 itasegm1\[405\]
rlabel metal3 333158 275688 333158 275688 0 itasegm1\[406\]
rlabel metal3 390096 284312 390096 284312 0 itasegm1\[407\]
rlabel metal3 333214 276808 333214 276808 0 itasegm1\[408\]
rlabel metal3 395584 242984 395584 242984 0 itasegm1\[409\]
rlabel metal3 258874 115528 258874 115528 0 itasegm1\[40\]
rlabel metal2 433818 284760 433818 284760 0 itasegm1\[410\]
rlabel metal3 333214 278488 333214 278488 0 itasegm1\[411\]
rlabel metal3 333998 279048 333998 279048 0 itasegm1\[412\]
rlabel metal3 333214 279608 333214 279608 0 itasegm1\[413\]
rlabel metal3 340270 280168 340270 280168 0 itasegm1\[414\]
rlabel metal3 331912 280910 331912 280910 0 itasegm1\[415\]
rlabel metal3 338590 281288 338590 281288 0 itasegm1\[416\]
rlabel metal3 455896 258510 455896 258510 0 itasegm1\[417\]
rlabel metal3 393638 282408 393638 282408 0 itasegm1\[418\]
rlabel metal3 456470 265720 456470 265720 0 itasegm1\[419\]
rlabel metal3 187558 52136 187558 52136 0 itasegm1\[41\]
rlabel metal2 475496 284648 475496 284648 0 itasegm1\[420\]
rlabel metal3 474474 263704 474474 263704 0 itasegm1\[421\]
rlabel metal3 331912 284578 331912 284578 0 itasegm1\[422\]
rlabel metal2 499576 285222 499576 285222 0 itasegm1\[423\]
rlabel metal3 474530 264376 474530 264376 0 itasegm1\[424\]
rlabel metal2 500248 285558 500248 285558 0 itasegm1\[425\]
rlabel metal4 352744 284984 352744 284984 0 itasegm1\[426\]
rlabel metal3 331912 287630 331912 287630 0 itasegm1\[427\]
rlabel metal2 498904 286398 498904 286398 0 itasegm1\[428\]
rlabel metal2 494200 242298 494200 242298 0 itasegm1\[429\]
rlabel metal2 222152 28770 222152 28770 0 itasegm1\[42\]
rlabel metal3 518574 260344 518574 260344 0 itasegm1\[430\]
rlabel metal3 424774 289688 424774 289688 0 itasegm1\[431\]
rlabel metal4 449400 287560 449400 287560 0 itasegm1\[432\]
rlabel metal3 333942 290808 333942 290808 0 itasegm1\[433\]
rlabel metal3 542752 286440 542752 286440 0 itasegm1\[434\]
rlabel metal4 430136 288344 430136 288344 0 itasegm1\[435\]
rlabel metal3 579880 261870 579880 261870 0 itasegm1\[436\]
rlabel metal4 523320 288064 523320 288064 0 itasegm1\[437\]
rlabel metal3 580622 259672 580622 259672 0 itasegm1\[438\]
rlabel metal3 579880 263270 579880 263270 0 itasegm1\[439\]
rlabel metal2 256312 106120 256312 106120 0 itasegm1\[43\]
rlabel metal3 579880 265958 579880 265958 0 itasegm1\[440\]
rlabel metal3 581742 266392 581742 266392 0 itasegm1\[441\]
rlabel metal2 560350 284760 560350 284760 0 itasegm1\[442\]
rlabel metal2 518280 293104 518280 293104 0 itasegm1\[443\]
rlabel metal2 563710 284760 563710 284760 0 itasegm1\[444\]
rlabel metal2 562002 284760 562002 284760 0 itasegm1\[445\]
rlabel metal3 333214 298088 333214 298088 0 itasegm1\[446\]
rlabel metal2 562296 242354 562296 242354 0 itasegm1\[447\]
rlabel metal2 261352 320040 261352 320040 0 itasegm1\[448\]
rlabel metal2 264600 341096 264600 341096 0 itasegm1\[449\]
rlabel metal2 232232 78022 232232 78022 0 itasegm1\[44\]
rlabel metal2 258104 320656 258104 320656 0 itasegm1\[450\]
rlabel metal4 263816 327639 263816 327639 0 itasegm1\[451\]
rlabel metal2 264712 340984 264712 340984 0 itasegm1\[452\]
rlabel metal3 20664 336658 20664 336658 0 itasegm1\[453\]
rlabel metal2 44296 356062 44296 356062 0 itasegm1\[454\]
rlabel metal2 256312 342664 256312 342664 0 itasegm1\[455\]
rlabel metal4 162568 331200 162568 331200 0 itasegm1\[456\]
rlabel metal4 263816 331029 263816 331029 0 itasegm1\[457\]
rlabel metal4 166264 330750 166264 330750 0 itasegm1\[458\]
rlabel metal2 45640 357070 45640 357070 0 itasegm1\[459\]
rlabel metal3 262962 118328 262962 118328 0 itasegm1\[45\]
rlabel metal4 263816 332139 263816 332139 0 itasegm1\[460\]
rlabel metal4 264712 338089 264712 338089 0 itasegm1\[461\]
rlabel metal4 264936 329909 264936 329909 0 itasegm1\[462\]
rlabel metal2 258104 345464 258104 345464 0 itasegm1\[463\]
rlabel metal4 260344 337669 260344 337669 0 itasegm1\[464\]
rlabel metal4 264040 333179 264040 333179 0 itasegm1\[465\]
rlabel metal3 178696 355656 178696 355656 0 itasegm1\[466\]
rlabel metal4 264600 331219 264600 331219 0 itasegm1\[467\]
rlabel metal2 99512 356118 99512 356118 0 itasegm1\[468\]
rlabel metal2 97496 357014 97496 357014 0 itasegm1\[469\]
rlabel metal2 264824 113624 264824 113624 0 itasegm1\[46\]
rlabel metal2 259672 346920 259672 346920 0 itasegm1\[470\]
rlabel metal2 261688 348432 261688 348432 0 itasegm1\[471\]
rlabel metal4 122696 339480 122696 339480 0 itasegm1\[472\]
rlabel metal2 100184 313978 100184 313978 0 itasegm1\[473\]
rlabel metal4 263928 341099 263928 341099 0 itasegm1\[474\]
rlabel metal4 263816 341289 263816 341289 0 itasegm1\[475\]
rlabel metal2 166264 356958 166264 356958 0 itasegm1\[476\]
rlabel metal3 189126 332920 189126 332920 0 itasegm1\[477\]
rlabel metal2 167608 313250 167608 313250 0 itasegm1\[478\]
rlabel metal2 186424 356104 186424 356104 0 itasegm1\[479\]
rlabel metal2 264936 116424 264936 116424 0 itasegm1\[47\]
rlabel metal3 190862 336280 190862 336280 0 itasegm1\[480\]
rlabel metal2 158200 356230 158200 356230 0 itasegm1\[481\]
rlabel metal3 189182 337624 189182 337624 0 itasegm1\[482\]
rlabel metal3 190806 335608 190806 335608 0 itasegm1\[483\]
rlabel metal3 187502 333592 187502 333592 0 itasegm1\[484\]
rlabel metal2 164248 313194 164248 313194 0 itasegm1\[485\]
rlabel metal3 187670 331576 187670 331576 0 itasegm1\[486\]
rlabel metal4 263816 347889 263816 347889 0 itasegm1\[487\]
rlabel metal2 262920 331576 262920 331576 0 itasegm1\[488\]
rlabel metal3 208656 355880 208656 355880 0 itasegm1\[489\]
rlabel metal3 204610 53480 204610 53480 0 itasegm1\[48\]
rlabel metal2 225512 357070 225512 357070 0 itasegm1\[490\]
rlabel metal4 263816 349819 263816 349819 0 itasegm1\[491\]
rlabel metal3 247912 350014 247912 350014 0 itasegm1\[492\]
rlabel metal2 261240 331632 261240 331632 0 itasegm1\[493\]
rlabel metal4 263368 350209 263368 350209 0 itasegm1\[494\]
rlabel metal4 264600 346360 264600 346360 0 itasegm1\[495\]
rlabel metal4 265160 344960 265160 344960 0 itasegm1\[496\]
rlabel metal2 263816 355096 263816 355096 0 itasegm1\[497\]
rlabel metal3 205450 332920 205450 332920 0 itasegm1\[498\]
rlabel metal3 263816 354368 263816 354368 0 itasegm1\[499\]
rlabel metal3 204554 52808 204554 52808 0 itasegm1\[49\]
rlabel metal2 167384 90160 167384 90160 0 itasegm1\[4\]
rlabel metal4 264824 345744 264824 345744 0 itasegm1\[500\]
rlabel metal3 204554 333592 204554 333592 0 itasegm1\[501\]
rlabel metal2 259560 335384 259560 335384 0 itasegm1\[502\]
rlabel metal3 204498 329560 204498 329560 0 itasegm1\[503\]
rlabel metal3 333158 326088 333158 326088 0 itasegm1\[504\]
rlabel metal4 350280 337699 350280 337699 0 itasegm1\[505\]
rlabel metal3 333214 327208 333214 327208 0 itasegm1\[506\]
rlabel metal3 333214 327768 333214 327768 0 itasegm1\[507\]
rlabel metal3 355040 314104 355040 314104 0 itasegm1\[508\]
rlabel metal3 335286 328888 335286 328888 0 itasegm1\[509\]
rlabel metal3 252070 53480 252070 53480 0 itasegm1\[50\]
rlabel metal4 344456 330729 344456 330729 0 itasegm1\[510\]
rlabel metal3 333214 330008 333214 330008 0 itasegm1\[511\]
rlabel metal2 378280 356286 378280 356286 0 itasegm1\[512\]
rlabel metal3 338646 331128 338646 331128 0 itasegm1\[513\]
rlabel metal3 333214 331688 333214 331688 0 itasegm1\[514\]
rlabel metal2 374248 356062 374248 356062 0 itasegm1\[515\]
rlabel metal2 374248 313754 374248 313754 0 itasegm1\[516\]
rlabel metal3 333214 333368 333214 333368 0 itasegm1\[517\]
rlabel metal2 444248 313922 444248 313922 0 itasegm1\[518\]
rlabel metal3 333214 334488 333214 334488 0 itasegm1\[519\]
rlabel metal3 253750 52808 253750 52808 0 itasegm1\[51\]
rlabel metal3 333214 335048 333214 335048 0 itasegm1\[520\]
rlabel metal4 351176 337589 351176 337589 0 itasegm1\[521\]
rlabel metal3 333214 336168 333214 336168 0 itasegm1\[522\]
rlabel metal3 333214 336728 333214 336728 0 itasegm1\[523\]
rlabel metal3 333158 337288 333158 337288 0 itasegm1\[524\]
rlabel metal3 333214 337848 333214 337848 0 itasegm1\[525\]
rlabel metal4 455336 331085 455336 331085 0 itasegm1\[526\]
rlabel metal3 333158 338968 333158 338968 0 itasegm1\[527\]
rlabel metal2 434840 313866 434840 313866 0 itasegm1\[528\]
rlabel metal3 333214 340088 333214 340088 0 itasegm1\[529\]
rlabel metal3 238168 29848 238168 29848 0 itasegm1\[52\]
rlabel metal3 333158 340648 333158 340648 0 itasegm1\[530\]
rlabel metal3 333214 341208 333214 341208 0 itasegm1\[531\]
rlabel metal2 500920 356230 500920 356230 0 itasegm1\[532\]
rlabel metal3 333158 342328 333158 342328 0 itasegm1\[533\]
rlabel metal2 496216 313978 496216 313978 0 itasegm1\[534\]
rlabel metal3 474642 349720 474642 349720 0 itasegm1\[535\]
rlabel metal3 419104 355544 419104 355544 0 itasegm1\[536\]
rlabel metal2 497560 356174 497560 356174 0 itasegm1\[537\]
rlabel metal3 519526 332920 519526 332920 0 itasegm1\[538\]
rlabel metal3 519470 332248 519470 332248 0 itasegm1\[539\]
rlabel metal3 249942 49448 249942 49448 0 itasegm1\[53\]
rlabel metal2 501354 355656 501354 355656 0 itasegm1\[540\]
rlabel metal2 351960 330680 351960 330680 0 itasegm1\[541\]
rlabel metal3 338590 347368 338590 347368 0 itasegm1\[542\]
rlabel metal2 500010 314104 500010 314104 0 itasegm1\[543\]
rlabel metal2 475496 355824 475496 355824 0 itasegm1\[544\]
rlabel metal2 495922 355880 495922 355880 0 itasegm1\[545\]
rlabel metal3 333214 349608 333214 349608 0 itasegm1\[546\]
rlabel metal3 333662 350168 333662 350168 0 itasegm1\[547\]
rlabel metal3 333214 350728 333214 350728 0 itasegm1\[548\]
rlabel metal4 352632 352072 352632 352072 0 itasegm1\[549\]
rlabel metal2 261464 109144 261464 109144 0 itasegm1\[54\]
rlabel metal3 335230 351848 335230 351848 0 itasegm1\[550\]
rlabel metal4 351064 352744 351064 352744 0 itasegm1\[551\]
rlabel metal3 455798 352968 455798 352968 0 itasegm1\[552\]
rlabel metal3 333158 353528 333158 353528 0 itasegm1\[553\]
rlabel metal3 456190 354088 456190 354088 0 itasegm1\[554\]
rlabel metal3 331912 354830 331912 354830 0 itasegm1\[555\]
rlabel metal3 331912 355334 331912 355334 0 itasegm1\[556\]
rlabel metal3 581518 337624 581518 337624 0 itasegm1\[557\]
rlabel metal3 580622 336952 580622 336952 0 itasegm1\[558\]
rlabel metal2 352744 357504 352744 357504 0 itasegm1\[559\]
rlabel metal2 264712 114464 264712 114464 0 itasegm1\[55\]
rlabel metal4 74872 389816 74872 389816 0 itasegm1\[560\]
rlabel metal3 20104 411866 20104 411866 0 itasegm1\[561\]
rlabel metal3 71694 406728 71694 406728 0 itasegm1\[562\]
rlabel metal2 69720 408072 69720 408072 0 itasegm1\[563\]
rlabel metal3 19978 410760 19978 410760 0 itasegm1\[564\]
rlabel metal4 73080 396256 73080 396256 0 itasegm1\[565\]
rlabel metal4 74760 398888 74760 398888 0 itasegm1\[566\]
rlabel metal2 264824 407904 264824 407904 0 itasegm1\[567\]
rlabel metal2 261352 407792 261352 407792 0 itasegm1\[568\]
rlabel metal2 171416 429184 171416 429184 0 itasegm1\[569\]
rlabel metal3 335342 93128 335342 93128 0 itasegm1\[56\]
rlabel metal4 263816 388920 263816 388920 0 itasegm1\[570\]
rlabel metal4 263928 389256 263928 389256 0 itasegm1\[571\]
rlabel metal3 20664 407050 20664 407050 0 itasegm1\[572\]
rlabel metal2 256200 410032 256200 410032 0 itasegm1\[573\]
rlabel metal2 257992 409248 257992 409248 0 itasegm1\[574\]
rlabel metal4 263816 392879 263816 392879 0 itasegm1\[575\]
rlabel metal2 256312 388976 256312 388976 0 itasegm1\[576\]
rlabel metal3 177968 384552 177968 384552 0 itasegm1\[577\]
rlabel metal2 102872 427854 102872 427854 0 itasegm1\[578\]
rlabel metal4 263928 395619 263928 395619 0 itasegm1\[579\]
rlabel metal4 396536 48384 396536 48384 0 itasegm1\[57\]
rlabel metal4 125160 401580 125160 401580 0 itasegm1\[580\]
rlabel metal3 176176 427000 176176 427000 0 itasegm1\[581\]
rlabel metal3 258762 396648 258762 396648 0 itasegm1\[582\]
rlabel metal2 264936 411936 264936 411936 0 itasegm1\[583\]
rlabel metal4 263816 397919 263816 397919 0 itasegm1\[584\]
rlabel metal4 263816 399009 263816 399009 0 itasegm1\[585\]
rlabel metal2 98168 428694 98168 428694 0 itasegm1\[586\]
rlabel metal2 258216 413168 258216 413168 0 itasegm1\[587\]
rlabel metal3 144424 407666 144424 407666 0 itasegm1\[588\]
rlabel metal3 187726 402024 187726 402024 0 itasegm1\[589\]
rlabel metal3 335230 94248 335230 94248 0 itasegm1\[58\]
rlabel metal3 257922 401128 257922 401128 0 itasegm1\[590\]
rlabel metal3 144312 406658 144312 406658 0 itasegm1\[591\]
rlabel metal3 258874 402248 258874 402248 0 itasegm1\[592\]
rlabel metal4 263816 402959 263816 402959 0 itasegm1\[593\]
rlabel metal3 144312 409654 144312 409654 0 itasegm1\[594\]
rlabel metal3 144312 408562 144312 408562 0 itasegm1\[595\]
rlabel metal3 187670 404712 187670 404712 0 itasegm1\[596\]
rlabel metal4 263928 406059 263928 406059 0 itasegm1\[597\]
rlabel metal2 164248 427910 164248 427910 0 itasegm1\[598\]
rlabel metal3 187614 403368 187614 403368 0 itasegm1\[599\]
rlabel metal2 355320 87416 355320 87416 0 itasegm1\[59\]
rlabel metal2 74760 61376 74760 61376 0 itasegm1\[5\]
rlabel metal3 187726 404040 187726 404040 0 itasegm1\[600\]
rlabel metal3 188734 406056 188734 406056 0 itasegm1\[601\]
rlabel metal2 263144 416976 263144 416976 0 itasegm1\[602\]
rlabel metal2 256312 417760 256312 417760 0 itasegm1\[603\]
rlabel metal4 260344 411979 260344 411979 0 itasegm1\[604\]
rlabel metal2 222152 428806 222152 428806 0 itasegm1\[605\]
rlabel metal2 240296 427966 240296 427966 0 itasegm1\[606\]
rlabel metal4 262136 411376 262136 411376 0 itasegm1\[607\]
rlabel metal2 261464 398384 261464 398384 0 itasegm1\[608\]
rlabel metal2 258104 398104 258104 398104 0 itasegm1\[609\]
rlabel metal4 396648 59136 396648 59136 0 itasegm1\[60\]
rlabel metal4 232232 426216 232232 426216 0 itasegm1\[610\]
rlabel metal4 263816 412319 263816 412319 0 itasegm1\[611\]
rlabel metal4 263368 410760 263368 410760 0 itasegm1\[612\]
rlabel metal4 262920 408688 262920 408688 0 itasegm1\[613\]
rlabel metal2 229278 427112 229278 427112 0 itasegm1\[614\]
rlabel metal4 263928 412664 263928 412664 0 itasegm1\[615\]
rlabel metal3 331912 384454 331912 384454 0 itasegm1\[616\]
rlabel metal2 352744 383432 352744 383432 0 itasegm1\[617\]
rlabel metal3 331912 385518 331912 385518 0 itasegm1\[618\]
rlabel metal3 331912 385938 331912 385938 0 itasegm1\[619\]
rlabel metal3 336126 95928 336126 95928 0 itasegm1\[61\]
rlabel metal3 334390 386568 334390 386568 0 itasegm1\[620\]
rlabel metal2 351176 385616 351176 385616 0 itasegm1\[621\]
rlabel metal3 335286 387688 335286 387688 0 itasegm1\[622\]
rlabel metal3 344176 403256 344176 403256 0 itasegm1\[623\]
rlabel metal3 333998 388808 333998 388808 0 itasegm1\[624\]
rlabel metal2 352632 387240 352632 387240 0 itasegm1\[625\]
rlabel metal3 355376 384216 355376 384216 0 itasegm1\[626\]
rlabel metal2 350616 387408 350616 387408 0 itasegm1\[627\]
rlabel metal2 347816 388416 347816 388416 0 itasegm1\[628\]
rlabel metal2 352520 388416 352520 388416 0 itasegm1\[629\]
rlabel metal2 350280 63112 350280 63112 0 itasegm1\[62\]
rlabel metal3 333214 392168 333214 392168 0 itasegm1\[630\]
rlabel metal3 333158 392728 333158 392728 0 itasegm1\[631\]
rlabel metal4 436856 426608 436856 426608 0 itasegm1\[632\]
rlabel metal3 333158 393848 333158 393848 0 itasegm1\[633\]
rlabel metal3 333214 394408 333214 394408 0 itasegm1\[634\]
rlabel metal2 435512 427910 435512 427910 0 itasegm1\[635\]
rlabel metal3 333158 395528 333158 395528 0 itasegm1\[636\]
rlabel metal3 333214 396088 333214 396088 0 itasegm1\[637\]
rlabel metal3 333158 396648 333158 396648 0 itasegm1\[638\]
rlabel metal3 333214 397208 333214 397208 0 itasegm1\[639\]
rlabel metal3 348642 47432 348642 47432 0 itasegm1\[63\]
rlabel metal2 350392 391104 350392 391104 0 itasegm1\[640\]
rlabel metal4 351064 400359 351064 400359 0 itasegm1\[641\]
rlabel metal3 333214 398888 333214 398888 0 itasegm1\[642\]
rlabel metal3 334110 399448 334110 399448 0 itasegm1\[643\]
rlabel metal3 335230 400008 335230 400008 0 itasegm1\[644\]
rlabel metal3 338702 400568 338702 400568 0 itasegm1\[645\]
rlabel metal3 333158 401128 333158 401128 0 itasegm1\[646\]
rlabel metal4 472136 420771 472136 420771 0 itasegm1\[647\]
rlabel metal2 352072 393288 352072 393288 0 itasegm1\[648\]
rlabel metal3 333214 402808 333214 402808 0 itasegm1\[649\]
rlabel metal3 346122 49448 346122 49448 0 itasegm1\[64\]
rlabel metal2 350280 394408 350280 394408 0 itasegm1\[650\]
rlabel metal3 333214 403928 333214 403928 0 itasegm1\[651\]
rlabel metal2 500920 427798 500920 427798 0 itasegm1\[652\]
rlabel metal2 352072 415688 352072 415688 0 itasegm1\[653\]
rlabel metal3 333998 405608 333998 405608 0 itasegm1\[654\]
rlabel metal3 337022 406168 337022 406168 0 itasegm1\[655\]
rlabel metal3 335342 406728 335342 406728 0 itasegm1\[656\]
rlabel metal3 334446 407288 334446 407288 0 itasegm1\[657\]
rlabel metal3 333214 407848 333214 407848 0 itasegm1\[658\]
rlabel metal3 333774 408408 333774 408408 0 itasegm1\[659\]
rlabel metal3 333214 98168 333214 98168 0 itasegm1\[65\]
rlabel metal3 454104 383992 454104 383992 0 itasegm1\[660\]
rlabel metal3 333214 409528 333214 409528 0 itasegm1\[661\]
rlabel metal3 333158 410088 333158 410088 0 itasegm1\[662\]
rlabel metal3 333662 410648 333662 410648 0 itasegm1\[663\]
rlabel metal3 333214 411208 333214 411208 0 itasegm1\[664\]
rlabel metal3 333214 411768 333214 411768 0 itasegm1\[665\]
rlabel metal3 333158 412328 333158 412328 0 itasegm1\[666\]
rlabel metal4 351064 411329 351064 411329 0 itasegm1\[667\]
rlabel metal3 333214 413448 333214 413448 0 itasegm1\[668\]
rlabel metal3 333550 414008 333550 414008 0 itasegm1\[669\]
rlabel metal3 347018 52136 347018 52136 0 itasegm1\[66\]
rlabel metal3 333214 414568 333214 414568 0 itasegm1\[670\]
rlabel metal3 333214 415128 333214 415128 0 itasegm1\[671\]
rlabel metal4 69720 475272 69720 475272 0 itasegm1\[672\]
rlabel metal4 264936 447104 264936 447104 0 itasegm1\[673\]
rlabel metal2 37576 498694 37576 498694 0 itasegm1\[674\]
rlabel metal3 174762 444248 174762 444248 0 itasegm1\[675\]
rlabel metal3 19082 475944 19082 475944 0 itasegm1\[676\]
rlabel metal2 36232 499646 36232 499646 0 itasegm1\[677\]
rlabel metal4 78344 461272 78344 461272 0 itasegm1\[678\]
rlabel metal4 73192 462560 73192 462560 0 itasegm1\[679\]
rlabel metal3 333326 99288 333326 99288 0 itasegm1\[67\]
rlabel metal3 121352 497784 121352 497784 0 itasegm1\[680\]
rlabel metal3 166474 447608 166474 447608 0 itasegm1\[681\]
rlabel metal3 143122 448168 143122 448168 0 itasegm1\[682\]
rlabel metal3 166586 448728 166586 448728 0 itasegm1\[683\]
rlabel metal3 166418 449288 166418 449288 0 itasegm1\[684\]
rlabel metal2 46984 498806 46984 498806 0 itasegm1\[685\]
rlabel metal4 143640 471912 143640 471912 0 itasegm1\[686\]
rlabel metal4 142184 456064 142184 456064 0 itasegm1\[687\]
rlabel metal3 175098 451528 175098 451528 0 itasegm1\[688\]
rlabel metal3 186130 452088 186130 452088 0 itasegm1\[689\]
rlabel metal3 333158 99848 333158 99848 0 itasegm1\[68\]
rlabel metal4 263816 454384 263816 454384 0 itasegm1\[690\]
rlabel metal3 185794 453208 185794 453208 0 itasegm1\[691\]
rlabel metal4 142072 469616 142072 469616 0 itasegm1\[692\]
rlabel metal4 138600 465304 138600 465304 0 itasegm1\[693\]
rlabel metal2 258104 476616 258104 476616 0 itasegm1\[694\]
rlabel metal3 124978 482664 124978 482664 0 itasegm1\[695\]
rlabel metal3 129598 476616 129598 476616 0 itasegm1\[696\]
rlabel metal2 98840 499758 98840 499758 0 itasegm1\[697\]
rlabel metal3 128758 479976 128758 479976 0 itasegm1\[698\]
rlabel metal4 127624 481208 127624 481208 0 itasegm1\[699\]
rlabel metal3 335286 100408 335286 100408 0 itasegm1\[69\]
rlabel metal4 69720 72576 69720 72576 0 itasegm1\[6\]
rlabel metal2 261576 478800 261576 478800 0 itasegm1\[700\]
rlabel metal3 195062 479304 195062 479304 0 itasegm1\[701\]
rlabel metal2 164248 498918 164248 498918 0 itasegm1\[702\]
rlabel metal3 142506 492744 142506 492744 0 itasegm1\[703\]
rlabel metal4 264152 465009 264152 465009 0 itasegm1\[704\]
rlabel metal2 256312 479472 256312 479472 0 itasegm1\[705\]
rlabel metal3 190414 477960 190414 477960 0 itasegm1\[706\]
rlabel metal3 142506 477288 142506 477288 0 itasegm1\[707\]
rlabel metal4 263816 463159 263816 463159 0 itasegm1\[708\]
rlabel metal3 187726 473928 187726 473928 0 itasegm1\[709\]
rlabel metal3 333606 100968 333606 100968 0 itasegm1\[70\]
rlabel metal3 187726 475944 187726 475944 0 itasegm1\[710\]
rlabel metal2 162582 498344 162582 498344 0 itasegm1\[711\]
rlabel metal3 144424 471562 144424 471562 0 itasegm1\[712\]
rlabel metal4 160888 457464 160888 457464 0 itasegm1\[713\]
rlabel metal4 259560 471352 259560 471352 0 itasegm1\[714\]
rlabel metal2 232232 498694 232232 498694 0 itasegm1\[715\]
rlabel metal3 237888 455224 237888 455224 0 itasegm1\[716\]
rlabel metal4 261352 474208 261352 474208 0 itasegm1\[717\]
rlabel metal2 258328 483784 258328 483784 0 itasegm1\[718\]
rlabel metal2 259560 462672 259560 462672 0 itasegm1\[719\]
rlabel metal3 333270 101528 333270 101528 0 itasegm1\[71\]
rlabel metal2 259896 485184 259896 485184 0 itasegm1\[720\]
rlabel metal4 262136 471968 262136 471968 0 itasegm1\[721\]
rlabel metal3 239680 455112 239680 455112 0 itasegm1\[722\]
rlabel metal2 256200 464632 256200 464632 0 itasegm1\[723\]
rlabel metal3 258034 471688 258034 471688 0 itasegm1\[724\]
rlabel metal3 260848 468664 260848 468664 0 itasegm1\[725\]
rlabel metal3 258090 472808 258090 472808 0 itasegm1\[726\]
rlabel metal4 263816 473519 263816 473519 0 itasegm1\[727\]
rlabel metal3 333886 442568 333886 442568 0 itasegm1\[728\]
rlabel metal3 333942 443128 333942 443128 0 itasegm1\[729\]
rlabel metal3 333214 102088 333214 102088 0 itasegm1\[72\]
rlabel metal3 335398 443688 335398 443688 0 itasegm1\[730\]
rlabel metal3 337022 444248 337022 444248 0 itasegm1\[731\]
rlabel metal4 396536 462616 396536 462616 0 itasegm1\[732\]
rlabel metal3 338646 445368 338646 445368 0 itasegm1\[733\]
rlabel metal2 374248 454034 374248 454034 0 itasegm1\[734\]
rlabel metal2 350504 472752 350504 472752 0 itasegm1\[735\]
rlabel metal4 396872 479360 396872 479360 0 itasegm1\[736\]
rlabel metal4 396760 469896 396760 469896 0 itasegm1\[737\]
rlabel metal2 352072 473032 352072 473032 0 itasegm1\[738\]
rlabel metal2 374248 498806 374248 498806 0 itasegm1\[739\]
rlabel metal2 351960 66080 351960 66080 0 itasegm1\[73\]
rlabel metal3 363510 449288 363510 449288 0 itasegm1\[740\]
rlabel metal3 338590 449848 338590 449848 0 itasegm1\[741\]
rlabel metal4 354424 453320 354424 453320 0 itasegm1\[742\]
rlabel metal4 399000 456904 399000 456904 0 itasegm1\[743\]
rlabel metal3 394870 451528 394870 451528 0 itasegm1\[744\]
rlabel metal3 333998 452088 333998 452088 0 itasegm1\[745\]
rlabel metal3 334054 452648 334054 452648 0 itasegm1\[746\]
rlabel metal3 334502 453208 334502 453208 0 itasegm1\[747\]
rlabel metal3 334838 453768 334838 453768 0 itasegm1\[748\]
rlabel metal3 394030 454328 394030 454328 0 itasegm1\[749\]
rlabel metal4 353640 87472 353640 87472 0 itasegm1\[74\]
rlabel metal3 394590 454888 394590 454888 0 itasegm1\[750\]
rlabel metal3 393750 455448 393750 455448 0 itasegm1\[751\]
rlabel metal2 430808 456218 430808 456218 0 itasegm1\[752\]
rlabel metal3 331912 456638 331912 456638 0 itasegm1\[753\]
rlabel metal3 331912 457058 331912 457058 0 itasegm1\[754\]
rlabel metal2 432824 498806 432824 498806 0 itasegm1\[755\]
rlabel metal2 474712 478072 474712 478072 0 itasegm1\[756\]
rlabel metal3 518238 477288 518238 477288 0 itasegm1\[757\]
rlabel metal3 517944 482258 517944 482258 0 itasegm1\[758\]
rlabel metal3 333662 459928 333662 459928 0 itasegm1\[759\]
rlabel metal4 350504 91840 350504 91840 0 itasegm1\[75\]
rlabel metal3 519526 473928 519526 473928 0 itasegm1\[760\]
rlabel metal3 333214 461048 333214 461048 0 itasegm1\[761\]
rlabel metal2 352632 459088 352632 459088 0 itasegm1\[762\]
rlabel metal2 351960 458696 351960 458696 0 itasegm1\[763\]
rlabel metal2 351064 460320 351064 460320 0 itasegm1\[764\]
rlabel metal2 352520 459872 352520 459872 0 itasegm1\[765\]
rlabel metal2 350280 459480 350280 459480 0 itasegm1\[766\]
rlabel metal3 333214 464408 333214 464408 0 itasegm1\[767\]
rlabel metal2 498904 454762 498904 454762 0 itasegm1\[768\]
rlabel metal3 419160 498120 419160 498120 0 itasegm1\[769\]
rlabel metal4 351176 102984 351176 102984 0 itasegm1\[76\]
rlabel metal3 495096 457856 495096 457856 0 itasegm1\[770\]
rlabel metal2 352184 482888 352184 482888 0 itasegm1\[771\]
rlabel metal3 336966 467208 336966 467208 0 itasegm1\[772\]
rlabel metal2 562968 498974 562968 498974 0 itasegm1\[773\]
rlabel metal3 336182 468328 336182 468328 0 itasegm1\[774\]
rlabel metal3 333214 468888 333214 468888 0 itasegm1\[775\]
rlabel metal3 336126 469448 336126 469448 0 itasegm1\[776\]
rlabel metal3 335230 470008 335230 470008 0 itasegm1\[777\]
rlabel metal3 333214 470568 333214 470568 0 itasegm1\[778\]
rlabel metal3 333158 471128 333158 471128 0 itasegm1\[779\]
rlabel metal3 412426 52136 412426 52136 0 itasegm1\[77\]
rlabel metal4 351064 470159 351064 470159 0 itasegm1\[780\]
rlabel metal3 333214 472248 333214 472248 0 itasegm1\[781\]
rlabel metal3 333550 472808 333550 472808 0 itasegm1\[782\]
rlabel metal3 333214 473368 333214 473368 0 itasegm1\[783\]
rlabel metal2 46984 570374 46984 570374 0 itasegm1\[784\]
rlabel metal3 99008 518504 99008 518504 0 itasegm1\[785\]
rlabel metal3 144074 501928 144074 501928 0 itasegm1\[786\]
rlabel metal3 63406 538440 63406 538440 0 itasegm1\[787\]
rlabel metal2 39592 515354 39592 515354 0 itasegm1\[788\]
rlabel metal2 46550 569464 46550 569464 0 itasegm1\[789\]
rlabel metal3 457310 54824 457310 54824 0 itasegm1\[78\]
rlabel metal3 19250 551880 19250 551880 0 itasegm1\[790\]
rlabel metal3 63462 544488 63462 544488 0 itasegm1\[791\]
rlabel metal3 63350 545832 63350 545832 0 itasegm1\[792\]
rlabel metal2 45640 570542 45640 570542 0 itasegm1\[793\]
rlabel metal3 63294 548520 63294 548520 0 itasegm1\[794\]
rlabel metal2 264600 538720 264600 538720 0 itasegm1\[795\]
rlabel metal4 261576 517888 261576 517888 0 itasegm1\[796\]
rlabel metal4 74872 529536 74872 529536 0 itasegm1\[797\]
rlabel metal4 143640 528584 143640 528584 0 itasegm1\[798\]
rlabel metal4 138600 527184 138600 527184 0 itasegm1\[799\]
rlabel metal3 457366 54152 457366 54152 0 itasegm1\[79\]
rlabel metal4 73080 74200 73080 74200 0 itasegm1\[7\]
rlabel metal2 192472 515816 192472 515816 0 itasegm1\[800\]
rlabel metal2 100184 525602 100184 525602 0 itasegm1\[801\]
rlabel metal3 125566 545832 125566 545832 0 itasegm1\[802\]
rlabel metal2 102872 519554 102872 519554 0 itasegm1\[803\]
rlabel metal2 99512 519834 99512 519834 0 itasegm1\[804\]
rlabel metal4 264936 515480 264936 515480 0 itasegm1\[805\]
rlabel metal3 125398 547848 125398 547848 0 itasegm1\[806\]
rlabel metal3 125510 547176 125510 547176 0 itasegm1\[807\]
rlabel metal4 263816 517104 263816 517104 0 itasegm1\[808\]
rlabel metal4 142072 530656 142072 530656 0 itasegm1\[809\]
rlabel metal3 333942 106568 333942 106568 0 itasegm1\[80\]
rlabel metal2 188104 518672 188104 518672 0 itasegm1\[810\]
rlabel metal3 175042 515928 175042 515928 0 itasegm1\[811\]
rlabel metal3 142562 563976 142562 563976 0 itasegm1\[812\]
rlabel metal2 168952 525658 168952 525658 0 itasegm1\[813\]
rlabel metal2 168952 569646 168952 569646 0 itasegm1\[814\]
rlabel metal2 169624 569758 169624 569758 0 itasegm1\[815\]
rlabel metal2 168280 523194 168280 523194 0 itasegm1\[816\]
rlabel metal2 162904 569702 162904 569702 0 itasegm1\[817\]
rlabel metal3 142408 546056 142408 546056 0 itasegm1\[818\]
rlabel metal3 143402 543144 143402 543144 0 itasegm1\[819\]
rlabel metal2 352520 92792 352520 92792 0 itasegm1\[81\]
rlabel metal3 142450 545160 142450 545160 0 itasegm1\[820\]
rlabel metal3 187670 545160 187670 545160 0 itasegm1\[821\]
rlabel metal3 187558 548520 187558 548520 0 itasegm1\[822\]
rlabel metal3 191646 545832 191646 545832 0 itasegm1\[823\]
rlabel metal3 143528 529144 143528 529144 0 itasegm1\[824\]
rlabel metal2 162904 525714 162904 525714 0 itasegm1\[825\]
rlabel metal3 249942 547176 249942 547176 0 itasegm1\[826\]
rlabel metal4 256312 534688 256312 534688 0 itasegm1\[827\]
rlabel metal2 224168 570374 224168 570374 0 itasegm1\[828\]
rlabel metal2 224728 526848 224728 526848 0 itasegm1\[829\]
rlabel metal2 350504 102312 350504 102312 0 itasegm1\[82\]
rlabel metal4 260008 535864 260008 535864 0 itasegm1\[830\]
rlabel metal2 259784 548576 259784 548576 0 itasegm1\[831\]
rlabel metal3 246442 527688 246442 527688 0 itasegm1\[832\]
rlabel metal2 227206 527912 227206 527912 0 itasegm1\[833\]
rlabel metal4 261352 540680 261352 540680 0 itasegm1\[834\]
rlabel metal4 263928 531384 263928 531384 0 itasegm1\[835\]
rlabel metal3 205968 549976 205968 549976 0 itasegm1\[836\]
rlabel metal2 263816 529144 263816 529144 0 itasegm1\[837\]
rlabel metal4 263816 532239 263816 532239 0 itasegm1\[838\]
rlabel metal3 251230 545832 251230 545832 0 itasegm1\[839\]
rlabel metal3 389368 29288 389368 29288 0 itasegm1\[83\]
rlabel metal2 376264 515410 376264 515410 0 itasegm1\[840\]
rlabel metal4 396648 523936 396648 523936 0 itasegm1\[841\]
rlabel metal3 333942 501928 333942 501928 0 itasegm1\[842\]
rlabel metal2 380296 569814 380296 569814 0 itasegm1\[843\]
rlabel metal3 393960 543522 393960 543522 0 itasegm1\[844\]
rlabel metal3 345282 549192 345282 549192 0 itasegm1\[845\]
rlabel metal2 352072 536592 352072 536592 0 itasegm1\[846\]
rlabel metal3 336126 504728 336126 504728 0 itasegm1\[847\]
rlabel metal2 377608 525546 377608 525546 0 itasegm1\[848\]
rlabel metal2 376936 525602 376936 525602 0 itasegm1\[849\]
rlabel metal3 519470 51464 519470 51464 0 itasegm1\[84\]
rlabel metal2 375242 569464 375242 569464 0 itasegm1\[850\]
rlabel metal3 361480 568904 361480 568904 0 itasegm1\[851\]
rlabel metal3 333158 507528 333158 507528 0 itasegm1\[852\]
rlabel metal3 336966 508088 336966 508088 0 itasegm1\[853\]
rlabel metal2 339304 510216 339304 510216 0 itasegm1\[854\]
rlabel metal2 435946 569464 435946 569464 0 itasegm1\[855\]
rlabel metal3 333214 509768 333214 509768 0 itasegm1\[856\]
rlabel metal4 354424 511000 354424 511000 0 itasegm1\[857\]
rlabel metal2 435512 569814 435512 569814 0 itasegm1\[858\]
rlabel metal2 428120 522242 428120 522242 0 itasegm1\[859\]
rlabel metal3 519638 43400 519638 43400 0 itasegm1\[85\]
rlabel metal4 355320 516096 355320 516096 0 itasegm1\[860\]
rlabel metal3 458304 546056 458304 546056 0 itasegm1\[861\]
rlabel metal3 457408 547736 457408 547736 0 itasegm1\[862\]
rlabel metal4 380520 516880 380520 516880 0 itasegm1\[863\]
rlabel metal3 333214 514248 333214 514248 0 itasegm1\[864\]
rlabel metal3 394478 514808 394478 514808 0 itasegm1\[865\]
rlabel metal2 381416 516152 381416 516152 0 itasegm1\[866\]
rlabel metal4 399000 529872 399000 529872 0 itasegm1\[867\]
rlabel metal2 356216 519120 356216 519120 0 itasegm1\[868\]
rlabel metal3 474754 553896 474754 553896 0 itasegm1\[869\]
rlabel metal3 519582 53480 519582 53480 0 itasegm1\[86\]
rlabel metal2 495194 569464 495194 569464 0 itasegm1\[870\]
rlabel metal3 517944 545426 517944 545426 0 itasegm1\[871\]
rlabel metal3 474642 552552 474642 552552 0 itasegm1\[872\]
rlabel metal3 518630 546504 518630 546504 0 itasegm1\[873\]
rlabel metal2 475496 521584 475496 521584 0 itasegm1\[874\]
rlabel metal2 379736 521920 379736 521920 0 itasegm1\[875\]
rlabel metal2 492562 569464 492562 569464 0 itasegm1\[876\]
rlabel metal2 501592 570654 501592 570654 0 itasegm1\[877\]
rlabel metal3 519414 543144 519414 543144 0 itasegm1\[878\]
rlabel metal3 517944 551138 517944 551138 0 itasegm1\[879\]
rlabel metal3 518574 50792 518574 50792 0 itasegm1\[87\]
rlabel metal2 500920 569758 500920 569758 0 itasegm1\[880\]
rlabel metal3 519582 541800 519582 541800 0 itasegm1\[881\]
rlabel metal2 564312 525994 564312 525994 0 itasegm1\[882\]
rlabel metal2 554232 570374 554232 570374 0 itasegm1\[883\]
rlabel metal2 562296 526554 562296 526554 0 itasegm1\[884\]
rlabel metal4 354424 527016 354424 527016 0 itasegm1\[885\]
rlabel metal3 581574 563976 581574 563976 0 itasegm1\[886\]
rlabel metal2 558264 570542 558264 570542 0 itasegm1\[887\]
rlabel metal3 445774 527688 445774 527688 0 itasegm1\[888\]
rlabel metal3 331912 528122 331912 528122 0 itasegm1\[889\]
rlabel metal3 422408 94920 422408 94920 0 itasegm1\[88\]
rlabel metal3 331912 528570 331912 528570 0 itasegm1\[890\]
rlabel metal2 539224 528584 539224 528584 0 itasegm1\[891\]
rlabel metal3 579880 551586 579880 551586 0 itasegm1\[892\]
rlabel metal4 523320 539504 523320 539504 0 itasegm1\[893\]
rlabel metal2 555576 570430 555576 570430 0 itasegm1\[894\]
rlabel metal2 554904 526722 554904 526722 0 itasegm1\[895\]
rlabel metal3 519526 52808 519526 52808 0 itasegm1\[89\]
rlabel metal3 201754 97608 201754 97608 0 itasegm1\[8\]
rlabel metal3 333718 112168 333718 112168 0 itasegm1\[90\]
rlabel metal3 518742 44072 518742 44072 0 itasegm1\[91\]
rlabel metal3 474474 44744 474474 44744 0 itasegm1\[92\]
rlabel metal2 494200 28042 494200 28042 0 itasegm1\[93\]
rlabel metal2 352072 101304 352072 101304 0 itasegm1\[94\]
rlabel metal2 498232 78806 498232 78806 0 itasegm1\[95\]
rlabel metal2 495544 28882 495544 28882 0 itasegm1\[96\]
rlabel metal3 333830 116088 333830 116088 0 itasegm1\[97\]
rlabel metal3 335286 116648 335286 116648 0 itasegm1\[98\]
rlabel metal3 333606 117208 333606 117208 0 itasegm1\[99\]
rlabel metal4 78120 74704 78120 74704 0 itasegm1\[9\]
rlabel metal2 264936 48720 264936 48720 0 itasel1\[0\]
rlabel metal4 73864 123329 73864 123329 0 itasel1\[100\]
rlabel metal2 263928 125384 263928 125384 0 itasel1\[101\]
rlabel metal5 166264 120960 166264 120960 0 itasel1\[102\]
rlabel metal4 263872 127170 263872 127170 0 itasel1\[103\]
rlabel metal3 20664 126910 20664 126910 0 itasel1\[104\]
rlabel metal4 263928 130419 263928 130419 0 itasel1\[105\]
rlabel metal4 263816 129349 263816 129349 0 itasel1\[106\]
rlabel metal4 260008 119177 260008 119177 0 itasel1\[107\]
rlabel metal2 102326 142296 102326 142296 0 itasel1\[108\]
rlabel metal3 260960 127624 260960 127624 0 itasel1\[109\]
rlabel metal2 45640 72590 45640 72590 0 itasel1\[10\]
rlabel metal2 99190 142072 99190 142072 0 itasel1\[110\]
rlabel metal3 178024 100520 178024 100520 0 itasel1\[111\]
rlabel metal4 138600 129420 138600 129420 0 itasel1\[112\]
rlabel metal4 263928 133379 263928 133379 0 itasel1\[113\]
rlabel metal3 81200 123928 81200 123928 0 itasel1\[114\]
rlabel metal2 98406 141960 98406 141960 0 itasel1\[115\]
rlabel metal2 102872 142702 102872 142702 0 itasel1\[116\]
rlabel metal4 143640 128520 143640 128520 0 itasel1\[117\]
rlabel metal4 263928 138264 263928 138264 0 itasel1\[118\]
rlabel metal2 106904 143598 106904 143598 0 itasel1\[119\]
rlabel metal2 45150 71064 45150 71064 0 itasel1\[11\]
rlabel metal3 143024 118440 143024 118440 0 itasel1\[120\]
rlabel metal3 192598 120568 192598 120568 0 itasel1\[121\]
rlabel metal3 190862 117208 190862 117208 0 itasel1\[122\]
rlabel metal3 141568 122696 141568 122696 0 itasel1\[123\]
rlabel metal3 195846 123256 195846 123256 0 itasel1\[124\]
rlabel metal3 183232 100968 183232 100968 0 itasel1\[125\]
rlabel metal3 187726 117880 187726 117880 0 itasel1\[126\]
rlabel metal2 187432 121800 187432 121800 0 itasel1\[127\]
rlabel metal2 192360 121520 192360 121520 0 itasel1\[128\]
rlabel metal3 187502 121240 187502 121240 0 itasel1\[129\]
rlabel metal3 81802 50120 81802 50120 0 itasel1\[12\]
rlabel metal3 187838 122584 187838 122584 0 itasel1\[130\]
rlabel metal3 142506 123928 142506 123928 0 itasel1\[131\]
rlabel metal3 205128 119224 205128 119224 0 itasel1\[132\]
rlabel metal3 204666 119896 204666 119896 0 itasel1\[133\]
rlabel metal2 224840 144046 224840 144046 0 itasel1\[134\]
rlabel metal3 261744 146104 261744 146104 0 itasel1\[135\]
rlabel metal3 254590 119896 254590 119896 0 itasel1\[136\]
rlabel metal3 204610 123928 204610 123928 0 itasel1\[137\]
rlabel metal2 232232 99610 232232 99610 0 itasel1\[138\]
rlabel metal2 226184 145446 226184 145446 0 itasel1\[139\]
rlabel metal2 102872 72310 102872 72310 0 itasel1\[13\]
rlabel metal2 237720 148176 237720 148176 0 itasel1\[140\]
rlabel metal3 253862 121240 253862 121240 0 itasel1\[141\]
rlabel metal3 253974 122584 253974 122584 0 itasel1\[142\]
rlabel metal3 254646 125944 254646 125944 0 itasel1\[143\]
rlabel metal2 373576 142702 373576 142702 0 itasel1\[144\]
rlabel metal3 338590 125048 338590 125048 0 itasel1\[145\]
rlabel metal3 333214 125608 333214 125608 0 itasel1\[146\]
rlabel metal2 350616 134680 350616 134680 0 itasel1\[147\]
rlabel metal3 333214 126728 333214 126728 0 itasel1\[148\]
rlabel metal3 347018 117208 347018 117208 0 itasel1\[149\]
rlabel metal3 124978 46760 124978 46760 0 itasel1\[14\]
rlabel metal3 347354 117880 347354 117880 0 itasel1\[150\]
rlabel metal2 352072 135464 352072 135464 0 itasel1\[151\]
rlabel metal2 372232 142590 372232 142590 0 itasel1\[152\]
rlabel metal3 334390 129528 334390 129528 0 itasel1\[153\]
rlabel metal3 347130 119896 347130 119896 0 itasel1\[154\]
rlabel metal3 359464 100632 359464 100632 0 itasel1\[155\]
rlabel metal5 396900 124290 396900 124290 0 itasel1\[156\]
rlabel metal3 333158 131768 333158 131768 0 itasel1\[157\]
rlabel metal3 333214 132328 333214 132328 0 itasel1\[158\]
rlabel metal4 351960 126879 351960 126879 0 itasel1\[159\]
rlabel metal2 105560 72870 105560 72870 0 itasel1\[15\]
rlabel metal4 411208 121865 411208 121865 0 itasel1\[160\]
rlabel metal2 430136 99554 430136 99554 0 itasel1\[161\]
rlabel metal3 333214 134568 333214 134568 0 itasel1\[162\]
rlabel metal3 333886 135128 333886 135128 0 itasel1\[163\]
rlabel metal2 352184 139328 352184 139328 0 itasel1\[164\]
rlabel metal2 432824 143542 432824 143542 0 itasel1\[165\]
rlabel metal2 437528 143430 437528 143430 0 itasel1\[166\]
rlabel metal2 352744 144312 352744 144312 0 itasel1\[167\]
rlabel metal2 420280 100520 420280 100520 0 itasel1\[168\]
rlabel metal2 351064 140112 351064 140112 0 itasel1\[169\]
rlabel metal3 81242 46760 81242 46760 0 itasel1\[16\]
rlabel metal3 333214 139048 333214 139048 0 itasel1\[170\]
rlabel metal2 498232 142590 498232 142590 0 itasel1\[171\]
rlabel metal3 518686 125944 518686 125944 0 itasel1\[172\]
rlabel metal3 333550 140728 333550 140728 0 itasel1\[173\]
rlabel metal3 331912 141470 331912 141470 0 itasel1\[174\]
rlabel metal4 517608 129192 517608 129192 0 itasel1\[175\]
rlabel metal2 500920 142702 500920 142702 0 itasel1\[176\]
rlabel metal3 333158 142968 333158 142968 0 itasel1\[177\]
rlabel metal2 492856 99666 492856 99666 0 itasel1\[178\]
rlabel metal3 518630 122584 518630 122584 0 itasel1\[179\]
rlabel metal4 263816 74424 263816 74424 0 itasel1\[17\]
rlabel metal3 579880 118230 579880 118230 0 itasel1\[180\]
rlabel metal3 456806 145208 456806 145208 0 itasel1\[181\]
rlabel metal2 561624 144046 561624 144046 0 itasel1\[182\]
rlabel metal3 580678 121912 580678 121912 0 itasel1\[183\]
rlabel metal3 579768 119518 579768 119518 0 itasel1\[184\]
rlabel metal3 580734 125272 580734 125272 0 itasel1\[185\]
rlabel metal3 333214 148008 333214 148008 0 itasel1\[186\]
rlabel metal4 449400 146160 449400 146160 0 itasel1\[187\]
rlabel metal4 523320 136864 523320 136864 0 itasel1\[188\]
rlabel metal4 525000 137480 525000 137480 0 itasel1\[189\]
rlabel metal2 100184 72926 100184 72926 0 itasel1\[18\]
rlabel metal3 532378 123256 532378 123256 0 itasel1\[190\]
rlabel metal3 546840 101080 546840 101080 0 itasel1\[191\]
rlabel metal2 264824 196784 264824 196784 0 itasel1\[192\]
rlabel metal2 261464 198128 261464 198128 0 itasel1\[193\]
rlabel metal4 187320 192060 187320 192060 0 itasel1\[194\]
rlabel metal2 249592 198968 249592 198968 0 itasel1\[195\]
rlabel metal3 20328 195370 20328 195370 0 itasel1\[196\]
rlabel metal3 20664 196266 20664 196266 0 itasel1\[197\]
rlabel metal2 265048 198520 265048 198520 0 itasel1\[198\]
rlabel metal4 258664 186519 258664 186519 0 itasel1\[199\]
rlabel metal4 188104 74144 188104 74144 0 itasel1\[19\]
rlabel metal2 35560 72646 35560 72646 0 itasel1\[1\]
rlabel metal2 263144 200312 263144 200312 0 itasel1\[200\]
rlabel metal2 256312 201880 256312 201880 0 itasel1\[201\]
rlabel metal4 188104 192330 188104 192330 0 itasel1\[202\]
rlabel metal2 263256 178920 263256 178920 0 itasel1\[203\]
rlabel metal4 169736 191790 169736 191790 0 itasel1\[204\]
rlabel metal4 262136 191619 262136 191619 0 itasel1\[205\]
rlabel metal2 259784 203000 259784 203000 0 itasel1\[206\]
rlabel metal4 258440 188669 258440 188669 0 itasel1\[207\]
rlabel metal4 263816 191919 263816 191919 0 itasel1\[208\]
rlabel metal3 176288 171640 176288 171640 0 itasel1\[209\]
rlabel metal3 81130 46088 81130 46088 0 itasel1\[20\]
rlabel metal2 101528 214718 101528 214718 0 itasel1\[210\]
rlabel metal4 169736 186660 169736 186660 0 itasel1\[211\]
rlabel metal3 114240 212744 114240 212744 0 itasel1\[212\]
rlabel metal2 258216 204904 258216 204904 0 itasel1\[213\]
rlabel metal2 98840 213654 98840 213654 0 itasel1\[214\]
rlabel metal2 98168 214382 98168 214382 0 itasel1\[215\]
rlabel metal3 187726 189784 187726 189784 0 itasel1\[216\]
rlabel metal3 187726 195832 187726 195832 0 itasel1\[217\]
rlabel metal4 263816 197059 263816 197059 0 itasel1\[218\]
rlabel metal4 263928 197249 263928 197249 0 itasel1\[219\]
rlabel metal4 127624 48328 127624 48328 0 itasel1\[21\]
rlabel metal2 162904 170506 162904 170506 0 itasel1\[220\]
rlabel metal4 263816 198619 263816 198619 0 itasel1\[221\]
rlabel metal3 208656 215656 208656 215656 0 itasel1\[222\]
rlabel metal2 247912 206304 247912 206304 0 itasel1\[223\]
rlabel metal2 186424 213136 186424 213136 0 itasel1\[224\]
rlabel metal2 254520 207536 254520 207536 0 itasel1\[225\]
rlabel metal2 168280 170450 168280 170450 0 itasel1\[226\]
rlabel metal2 162232 170394 162232 170394 0 itasel1\[227\]
rlabel metal2 222824 214662 222824 214662 0 itasel1\[228\]
rlabel metal3 231560 212352 231560 212352 0 itasel1\[229\]
rlabel metal2 122696 28840 122696 28840 0 itasel1\[22\]
rlabel metal4 231784 212576 231784 212576 0 itasel1\[230\]
rlabel metal2 256536 210056 256536 210056 0 itasel1\[231\]
rlabel metal4 264600 198184 264600 198184 0 itasel1\[232\]
rlabel metal4 264824 199752 264824 199752 0 itasel1\[233\]
rlabel metal4 258104 197680 258104 197680 0 itasel1\[234\]
rlabel metal4 262136 206319 262136 206319 0 itasel1\[235\]
rlabel metal2 228872 214326 228872 214326 0 itasel1\[236\]
rlabel metal2 228200 171346 228200 171346 0 itasel1\[237\]
rlabel metal2 225512 170338 225512 170338 0 itasel1\[238\]
rlabel metal3 249942 187096 249942 187096 0 itasel1\[239\]
rlabel metal2 125160 52976 125160 52976 0 itasel1\[23\]
rlabel metal2 352184 177240 352184 177240 0 itasel1\[240\]
rlabel metal3 333550 183288 333550 183288 0 itasel1\[241\]
rlabel metal3 375816 212576 375816 212576 0 itasel1\[242\]
rlabel metal4 396536 190217 396536 190217 0 itasel1\[243\]
rlabel metal2 376264 213654 376264 213654 0 itasel1\[244\]
rlabel metal4 346136 186984 346136 186984 0 itasel1\[245\]
rlabel metal3 336910 186088 336910 186088 0 itasel1\[246\]
rlabel metal4 342664 186429 342664 186429 0 itasel1\[247\]
rlabel metal2 350616 179424 350616 179424 0 itasel1\[248\]
rlabel metal2 377608 170338 377608 170338 0 itasel1\[249\]
rlabel metal4 144088 52444 144088 52444 0 itasel1\[24\]
rlabel metal2 373576 170506 373576 170506 0 itasel1\[250\]
rlabel metal2 350392 201992 350392 201992 0 itasel1\[251\]
rlabel metal4 347816 190979 347816 190979 0 itasel1\[252\]
rlabel metal3 333998 190008 333998 190008 0 itasel1\[253\]
rlabel metal3 333158 190568 333158 190568 0 itasel1\[254\]
rlabel metal3 331912 191058 331912 191058 0 itasel1\[255\]
rlabel metal3 338758 191688 338758 191688 0 itasel1\[256\]
rlabel metal3 333214 192248 333214 192248 0 itasel1\[257\]
rlabel metal3 338646 192808 338646 192808 0 itasel1\[258\]
rlabel metal3 333214 193368 333214 193368 0 itasel1\[259\]
rlabel metal3 143346 52808 143346 52808 0 itasel1\[25\]
rlabel metal3 333158 193928 333158 193928 0 itasel1\[260\]
rlabel metal3 333214 194488 333214 194488 0 itasel1\[261\]
rlabel metal3 331912 195230 331912 195230 0 itasel1\[262\]
rlabel metal3 335230 195608 335230 195608 0 itasel1\[263\]
rlabel metal3 333214 196168 333214 196168 0 itasel1\[264\]
rlabel metal2 350504 205072 350504 205072 0 itasel1\[265\]
rlabel metal3 333214 197288 333214 197288 0 itasel1\[266\]
rlabel metal4 472136 191744 472136 191744 0 itasel1\[267\]
rlabel metal2 475496 213304 475496 213304 0 itasel1\[268\]
rlabel metal4 472136 194783 472136 194783 0 itasel1\[269\]
rlabel metal4 144312 64176 144312 64176 0 itasel1\[26\]
rlabel metal2 493528 171458 493528 171458 0 itasel1\[270\]
rlabel metal2 492184 214438 492184 214438 0 itasel1\[271\]
rlabel metal3 471954 196504 471954 196504 0 itasel1\[272\]
rlabel metal2 495544 214494 495544 214494 0 itasel1\[273\]
rlabel metal4 472136 187553 472136 187553 0 itasel1\[274\]
rlabel metal3 518574 189784 518574 189784 0 itasel1\[275\]
rlabel metal3 333606 202888 333606 202888 0 itasel1\[276\]
rlabel metal3 536802 195832 536802 195832 0 itasel1\[277\]
rlabel metal3 449848 212968 449848 212968 0 itasel1\[278\]
rlabel metal3 333214 204568 333214 204568 0 itasel1\[279\]
rlabel metal3 143080 49224 143080 49224 0 itasel1\[27\]
rlabel metal2 562856 170632 562856 170632 0 itasel1\[280\]
rlabel metal2 539224 213080 539224 213080 0 itasel1\[281\]
rlabel metal3 333214 206248 333214 206248 0 itasel1\[282\]
rlabel metal2 563640 214382 563640 214382 0 itasel1\[283\]
rlabel metal2 562968 214606 562968 214606 0 itasel1\[284\]
rlabel metal4 351176 209272 351176 209272 0 itasel1\[285\]
rlabel metal3 333550 208488 333550 208488 0 itasel1\[286\]
rlabel metal4 351064 209720 351064 209720 0 itasel1\[287\]
rlabel metal3 144074 240968 144074 240968 0 itasel1\[288\]
rlabel metal2 192360 262920 192360 262920 0 itasel1\[289\]
rlabel metal2 187320 55104 187320 55104 0 itasel1\[28\]
rlabel metal4 21000 243712 21000 243712 0 itasel1\[290\]
rlabel metal3 63070 263032 63070 263032 0 itasel1\[291\]
rlabel metal4 69720 254128 69720 254128 0 itasel1\[292\]
rlabel metal3 258216 285880 258216 285880 0 itasel1\[293\]
rlabel metal3 71750 258328 71750 258328 0 itasel1\[294\]
rlabel metal3 63350 261688 63350 261688 0 itasel1\[295\]
rlabel metal3 63294 260344 63294 260344 0 itasel1\[296\]
rlabel metal2 44702 284760 44702 284760 0 itasel1\[297\]
rlabel metal2 38248 242298 38248 242298 0 itasel1\[298\]
rlabel metal2 46312 241402 46312 241402 0 itasel1\[299\]
rlabel metal3 142394 53480 142394 53480 0 itasel1\[29\]
rlabel metal4 76440 54460 76440 54460 0 itasel1\[2\]
rlabel metal2 106232 242242 106232 242242 0 itasel1\[300\]
rlabel metal3 177184 284424 177184 284424 0 itasel1\[301\]
rlabel metal4 260344 251619 260344 251619 0 itasel1\[302\]
rlabel metal3 179368 242984 179368 242984 0 itasel1\[303\]
rlabel metal2 106232 285390 106232 285390 0 itasel1\[304\]
rlabel metal4 263816 250389 263816 250389 0 itasel1\[305\]
rlabel metal4 263816 251479 263816 251479 0 itasel1\[306\]
rlabel metal2 98840 286286 98840 286286 0 itasel1\[307\]
rlabel metal2 98168 286174 98168 286174 0 itasel1\[308\]
rlabel metal4 125160 256410 125160 256410 0 itasel1\[309\]
rlabel metal3 142450 54152 142450 54152 0 itasel1\[30\]
rlabel metal4 263816 253409 263816 253409 0 itasel1\[310\]
rlabel metal4 263816 254589 263816 254589 0 itasel1\[311\]
rlabel metal2 262920 281820 262920 281820 0 itasel1\[312\]
rlabel metal2 164248 285446 164248 285446 0 itasel1\[313\]
rlabel metal2 162904 286286 162904 286286 0 itasel1\[314\]
rlabel metal2 166936 286342 166936 286342 0 itasel1\[315\]
rlabel metal3 187726 266392 187726 266392 0 itasel1\[316\]
rlabel metal4 260008 260949 260008 260949 0 itasel1\[317\]
rlabel metal3 185864 262234 185864 262234 0 itasel1\[318\]
rlabel metal3 143346 266392 143346 266392 0 itasel1\[319\]
rlabel metal3 142506 45416 142506 45416 0 itasel1\[31\]
rlabel metal2 163576 241290 163576 241290 0 itasel1\[320\]
rlabel metal4 263928 259819 263928 259819 0 itasel1\[321\]
rlabel metal3 144312 263242 144312 263242 0 itasel1\[322\]
rlabel metal2 166264 242130 166264 242130 0 itasel1\[323\]
rlabel metal4 262472 264096 262472 264096 0 itasel1\[324\]
rlabel metal4 262248 263704 262248 263704 0 itasel1\[325\]
rlabel metal3 247912 262794 247912 262794 0 itasel1\[326\]
rlabel metal4 262136 261912 262136 261912 0 itasel1\[327\]
rlabel metal4 262360 261184 262360 261184 0 itasel1\[328\]
rlabel metal2 228200 286062 228200 286062 0 itasel1\[329\]
rlabel metal3 187726 46088 187726 46088 0 itasel1\[32\]
rlabel metal4 264040 261072 264040 261072 0 itasel1\[330\]
rlabel metal3 235872 243096 235872 243096 0 itasel1\[331\]
rlabel metal4 260344 263619 260344 263619 0 itasel1\[332\]
rlabel metal4 263816 266329 263816 266329 0 itasel1\[333\]
rlabel metal4 263816 266879 263816 266879 0 itasel1\[334\]
rlabel metal2 222824 241514 222824 241514 0 itasel1\[335\]
rlabel metal4 396648 252056 396648 252056 0 itasel1\[336\]
rlabel metal3 363454 241528 363454 241528 0 itasel1\[337\]
rlabel metal2 359576 241136 359576 241136 0 itasel1\[338\]
rlabel metal3 363510 242648 363510 242648 0 itasel1\[339\]
rlabel metal2 163576 72926 163576 72926 0 itasel1\[33\]
rlabel metal2 376264 286286 376264 286286 0 itasel1\[340\]
rlabel metal3 333998 243768 333998 243768 0 itasel1\[341\]
rlabel metal3 334390 244328 334390 244328 0 itasel1\[342\]
rlabel metal3 348642 267064 348642 267064 0 itasel1\[343\]
rlabel metal2 349496 243656 349496 243656 0 itasel1\[344\]
rlabel metal3 350434 261016 350434 261016 0 itasel1\[345\]
rlabel metal3 349482 259672 349482 259672 0 itasel1\[346\]
rlabel metal3 335230 247128 335230 247128 0 itasel1\[347\]
rlabel metal4 351064 246736 351064 246736 0 itasel1\[348\]
rlabel metal3 333214 248248 333214 248248 0 itasel1\[349\]
rlabel metal3 142338 46088 142338 46088 0 itasel1\[34\]
rlabel metal3 333214 248808 333214 248808 0 itasel1\[350\]
rlabel metal2 350280 268520 350280 268520 0 itasel1\[351\]
rlabel metal2 439138 284760 439138 284760 0 itasel1\[352\]
rlabel metal3 333158 250488 333158 250488 0 itasel1\[353\]
rlabel metal4 351064 250669 351064 250669 0 itasel1\[354\]
rlabel metal3 333214 251608 333214 251608 0 itasel1\[355\]
rlabel metal2 352184 247688 352184 247688 0 itasel1\[356\]
rlabel metal3 333214 252728 333214 252728 0 itasel1\[357\]
rlabel metal2 350392 247352 350392 247352 0 itasel1\[358\]
rlabel metal3 333158 253848 333158 253848 0 itasel1\[359\]
rlabel metal3 191646 47432 191646 47432 0 itasel1\[35\]
rlabel metal4 472136 265496 472136 265496 0 itasel1\[360\]
rlabel metal3 333214 254968 333214 254968 0 itasel1\[361\]
rlabel metal3 333270 255528 333270 255528 0 itasel1\[362\]
rlabel metal4 351064 257419 351064 257419 0 itasel1\[363\]
rlabel metal4 351960 261929 351960 261929 0 itasel1\[364\]
rlabel metal3 333550 257208 333550 257208 0 itasel1\[365\]
rlabel metal3 333158 257768 333158 257768 0 itasel1\[366\]
rlabel metal3 333214 258328 333214 258328 0 itasel1\[367\]
rlabel metal3 333214 258888 333214 258888 0 itasel1\[368\]
rlabel metal2 498232 286118 498232 286118 0 itasel1\[369\]
rlabel metal3 205968 45976 205968 45976 0 itasel1\[36\]
rlabel metal3 333214 260008 333214 260008 0 itasel1\[370\]
rlabel metal3 331912 260498 331912 260498 0 itasel1\[371\]
rlabel metal3 331912 260890 331912 260890 0 itasel1\[372\]
rlabel metal3 333214 261688 333214 261688 0 itasel1\[373\]
rlabel metal3 336182 262248 336182 262248 0 itasel1\[374\]
rlabel metal3 333214 262808 333214 262808 0 itasel1\[375\]
rlabel metal3 333662 263368 333662 263368 0 itasel1\[376\]
rlabel metal3 333214 263928 333214 263928 0 itasel1\[377\]
rlabel metal3 333214 264488 333214 264488 0 itasel1\[378\]
rlabel metal3 335286 265048 335286 265048 0 itasel1\[379\]
rlabel metal4 264600 80864 264600 80864 0 itasel1\[37\]
rlabel metal3 333718 265608 333718 265608 0 itasel1\[380\]
rlabel metal3 333214 266168 333214 266168 0 itasel1\[381\]
rlabel metal3 333606 266728 333606 266728 0 itasel1\[382\]
rlabel metal3 333214 267288 333214 267288 0 itasel1\[383\]
rlabel metal3 19250 334936 19250 334936 0 itasel1\[384\]
rlabel metal3 19138 332248 19138 332248 0 itasel1\[385\]
rlabel metal2 74760 329112 74760 329112 0 itasel1\[386\]
rlabel metal2 36904 307482 36904 307482 0 itasel1\[387\]
rlabel metal2 35560 356958 35560 356958 0 itasel1\[388\]
rlabel metal3 19194 336280 19194 336280 0 itasel1\[389\]
rlabel metal3 261576 77336 261576 77336 0 itasel1\[38\]
rlabel metal2 43624 308322 43624 308322 0 itasel1\[390\]
rlabel metal2 40936 356118 40936 356118 0 itasel1\[391\]
rlabel metal3 63294 332920 63294 332920 0 itasel1\[392\]
rlabel metal4 263816 306264 263816 306264 0 itasel1\[393\]
rlabel metal3 63350 335608 63350 335608 0 itasel1\[394\]
rlabel metal2 38920 309722 38920 309722 0 itasel1\[395\]
rlabel metal2 106232 310002 106232 310002 0 itasel1\[396\]
rlabel metal2 99512 310282 99512 310282 0 itasel1\[397\]
rlabel metal2 101528 310562 101528 310562 0 itasel1\[398\]
rlabel metal4 141960 322504 141960 322504 0 itasel1\[399\]
rlabel metal3 205506 56168 205506 56168 0 itasel1\[39\]
rlabel metal4 20104 61712 20104 61712 0 itasel1\[3\]
rlabel metal3 81032 331464 81032 331464 0 itasel1\[400\]
rlabel metal2 104216 311402 104216 311402 0 itasel1\[401\]
rlabel metal3 125398 330232 125398 330232 0 itasel1\[402\]
rlabel metal2 166264 310744 166264 310744 0 itasel1\[403\]
rlabel metal4 143640 324464 143640 324464 0 itasel1\[404\]
rlabel metal2 100856 356958 100856 356958 0 itasel1\[405\]
rlabel metal4 161336 313096 161336 313096 0 itasel1\[406\]
rlabel metal3 81312 329336 81312 329336 0 itasel1\[407\]
rlabel metal3 234514 312648 234514 312648 0 itasel1\[408\]
rlabel metal2 163576 357014 163576 357014 0 itasel1\[409\]
rlabel metal2 223496 72982 223496 72982 0 itasel1\[40\]
rlabel metal3 195846 332248 195846 332248 0 itasel1\[410\]
rlabel metal3 142562 340312 142562 340312 0 itasel1\[411\]
rlabel metal2 187544 334992 187544 334992 0 itasel1\[412\]
rlabel metal2 166936 356286 166936 356286 0 itasel1\[413\]
rlabel metal3 187726 340312 187726 340312 0 itasel1\[414\]
rlabel metal3 142506 337624 142506 337624 0 itasel1\[415\]
rlabel metal3 187446 336952 187446 336952 0 itasel1\[416\]
rlabel metal2 248584 316120 248584 316120 0 itasel1\[417\]
rlabel metal2 168952 313138 168952 313138 0 itasel1\[418\]
rlabel metal2 160216 313922 160216 313922 0 itasel1\[419\]
rlabel metal3 231840 29232 231840 29232 0 itasel1\[41\]
rlabel metal2 229544 357126 229544 357126 0 itasel1\[420\]
rlabel metal2 224168 312970 224168 312970 0 itasel1\[421\]
rlabel metal4 261352 326368 261352 326368 0 itasel1\[422\]
rlabel metal2 223118 355880 223118 355880 0 itasel1\[423\]
rlabel metal3 249942 330232 249942 330232 0 itasel1\[424\]
rlabel metal4 261240 329896 261240 329896 0 itasel1\[425\]
rlabel metal4 259560 326144 259560 326144 0 itasel1\[426\]
rlabel metal2 257992 340704 257992 340704 0 itasel1\[427\]
rlabel metal4 263816 323969 263816 323969 0 itasel1\[428\]
rlabel metal2 232232 356006 232232 356006 0 itasel1\[429\]
rlabel metal2 225512 80430 225512 80430 0 itasel1\[42\]
rlabel metal3 249494 334264 249494 334264 0 itasel1\[430\]
rlabel via4 263816 325529 263816 325529 0 itasel1\[431\]
rlabel metal4 396536 333648 396536 333648 0 itasel1\[432\]
rlabel metal3 345282 330232 345282 330232 0 itasel1\[433\]
rlabel metal3 333550 300328 333550 300328 0 itasel1\[434\]
rlabel metal3 336910 300888 336910 300888 0 itasel1\[435\]
rlabel metal2 370888 357126 370888 357126 0 itasel1\[436\]
rlabel metal3 352086 302008 352086 302008 0 itasel1\[437\]
rlabel metal4 396872 317632 396872 317632 0 itasel1\[438\]
rlabel metal2 370216 308602 370216 308602 0 itasel1\[439\]
rlabel metal2 224840 72926 224840 72926 0 itasel1\[43\]
rlabel metal2 373576 308882 373576 308882 0 itasel1\[440\]
rlabel metal2 376264 309162 376264 309162 0 itasel1\[441\]
rlabel metal3 334446 304808 334446 304808 0 itasel1\[442\]
rlabel metal3 338590 305368 338590 305368 0 itasel1\[443\]
rlabel metal3 394870 305928 394870 305928 0 itasel1\[444\]
rlabel metal2 430808 310282 430808 310282 0 itasel1\[445\]
rlabel metal2 430808 356062 430808 356062 0 itasel1\[446\]
rlabel metal3 362950 307608 362950 307608 0 itasel1\[447\]
rlabel metal3 371350 308168 371350 308168 0 itasel1\[448\]
rlabel metal2 433496 311402 433496 311402 0 itasel1\[449\]
rlabel metal2 231560 28714 231560 28714 0 itasel1\[44\]
rlabel metal2 430136 311682 430136 311682 0 itasel1\[450\]
rlabel metal2 402360 334152 402360 334152 0 itasel1\[451\]
rlabel metal2 400680 333536 400680 333536 0 itasel1\[452\]
rlabel metal2 399000 333872 399000 333872 0 itasel1\[453\]
rlabel metal2 437528 312802 437528 312802 0 itasel1\[454\]
rlabel metal2 436184 313082 436184 313082 0 itasel1\[455\]
rlabel metal3 333830 312648 333830 312648 0 itasel1\[456\]
rlabel metal3 474474 338968 474474 338968 0 itasel1\[457\]
rlabel metal3 334558 313768 334558 313768 0 itasel1\[458\]
rlabel metal4 517496 325976 517496 325976 0 itasel1\[459\]
rlabel metal3 260904 85736 260904 85736 0 itasel1\[45\]
rlabel metal3 474642 339640 474642 339640 0 itasel1\[460\]
rlabel metal3 474586 333592 474586 333592 0 itasel1\[461\]
rlabel metal2 498232 357126 498232 357126 0 itasel1\[462\]
rlabel metal3 518574 335608 518574 335608 0 itasel1\[463\]
rlabel metal3 519414 336952 519414 336952 0 itasel1\[464\]
rlabel metal2 496888 312914 496888 312914 0 itasel1\[465\]
rlabel metal2 499576 313810 499576 313810 0 itasel1\[466\]
rlabel metal3 333214 318808 333214 318808 0 itasel1\[467\]
rlabel metal2 562296 313138 562296 313138 0 itasel1\[468\]
rlabel metal3 333214 319928 333214 319928 0 itasel1\[469\]
rlabel metal3 254590 52136 254590 52136 0 itasel1\[46\]
rlabel metal4 562968 314057 562968 314057 0 itasel1\[470\]
rlabel metal3 333718 321048 333718 321048 0 itasel1\[471\]
rlabel metal3 333214 321608 333214 321608 0 itasel1\[472\]
rlabel metal2 553560 313026 553560 313026 0 itasel1\[473\]
rlabel metal3 333158 322728 333158 322728 0 itasel1\[474\]
rlabel metal2 558026 314104 558026 314104 0 itasel1\[475\]
rlabel metal3 333214 323848 333214 323848 0 itasel1\[476\]
rlabel metal3 333214 324408 333214 324408 0 itasel1\[477\]
rlabel metal2 557592 356958 557592 356958 0 itasel1\[478\]
rlabel metal3 333214 325528 333214 325528 0 itasel1\[479\]
rlabel metal3 204498 54152 204498 54152 0 itasel1\[47\]
rlabel metal4 264600 368144 264600 368144 0 itasel1\[480\]
rlabel metal2 261464 369264 261464 369264 0 itasel1\[481\]
rlabel metal4 264824 368816 264824 368816 0 itasel1\[482\]
rlabel metal3 145040 380632 145040 380632 0 itasel1\[483\]
rlabel metal3 63294 406056 63294 406056 0 itasel1\[484\]
rlabel metal3 63406 401352 63406 401352 0 itasel1\[485\]
rlabel metal2 73080 393680 73080 393680 0 itasel1\[486\]
rlabel metal4 69720 393960 69720 393960 0 itasel1\[487\]
rlabel metal3 19082 411432 19082 411432 0 itasel1\[488\]
rlabel metal3 19194 408072 19194 408072 0 itasel1\[489\]
rlabel metal3 331912 66318 331912 66318 0 itasel1\[48\]
rlabel metal4 76440 389760 76440 389760 0 itasel1\[490\]
rlabel metal4 257880 371280 257880 371280 0 itasel1\[491\]
rlabel metal4 143640 383432 143640 383432 0 itasel1\[492\]
rlabel metal3 125566 406056 125566 406056 0 itasel1\[493\]
rlabel metal3 125398 410088 125398 410088 0 itasel1\[494\]
rlabel metal2 100184 375578 100184 375578 0 itasel1\[495\]
rlabel metal3 125454 404040 125454 404040 0 itasel1\[496\]
rlabel metal2 107576 376138 107576 376138 0 itasel1\[497\]
rlabel metal2 100856 376418 100856 376418 0 itasel1\[498\]
rlabel metal3 125622 408744 125622 408744 0 itasel1\[499\]
rlabel metal2 376936 72646 376936 72646 0 itasel1\[49\]
rlabel metal3 20104 47838 20104 47838 0 itasel1\[4\]
rlabel metal2 103544 376978 103544 376978 0 itasel1\[500\]
rlabel metal3 125510 410760 125510 410760 0 itasel1\[501\]
rlabel metal2 263816 371784 263816 371784 0 itasel1\[502\]
rlabel metal4 264936 375536 264936 375536 0 itasel1\[503\]
rlabel metal2 162904 428862 162904 428862 0 itasel1\[504\]
rlabel metal3 187446 408072 187446 408072 0 itasel1\[505\]
rlabel metal3 189126 401352 189126 401352 0 itasel1\[506\]
rlabel metal2 161560 428638 161560 428638 0 itasel1\[507\]
rlabel metal2 187432 399560 187432 399560 0 itasel1\[508\]
rlabel metal2 189000 400400 189000 400400 0 itasel1\[509\]
rlabel metal3 331912 67550 331912 67550 0 itasel1\[50\]
rlabel metal3 143402 410088 143402 410088 0 itasel1\[510\]
rlabel metal2 165592 427966 165592 427966 0 itasel1\[511\]
rlabel metal2 168952 428806 168952 428806 0 itasel1\[512\]
rlabel metal2 189112 401016 189112 401016 0 itasel1\[513\]
rlabel metal2 167608 380898 167608 380898 0 itasel1\[514\]
rlabel metal3 142562 403368 142562 403368 0 itasel1\[515\]
rlabel metal3 248794 377608 248794 377608 0 itasel1\[516\]
rlabel metal3 260848 383096 260848 383096 0 itasel1\[517\]
rlabel metal4 256200 393064 256200 393064 0 itasel1\[518\]
rlabel metal2 259560 404824 259560 404824 0 itasel1\[519\]
rlabel metal3 349426 54152 349426 54152 0 itasel1\[51\]
rlabel metal2 261240 405048 261240 405048 0 itasel1\[520\]
rlabel metal3 205506 408072 205506 408072 0 itasel1\[521\]
rlabel metal2 263032 405552 263032 405552 0 itasel1\[522\]
rlabel metal3 237090 381528 237090 381528 0 itasel1\[523\]
rlabel metal4 265048 385504 265048 385504 0 itasel1\[524\]
rlabel metal3 261688 386344 261688 386344 0 itasel1\[525\]
rlabel metal4 259672 392952 259672 392952 0 itasel1\[526\]
rlabel metal3 235634 383768 235634 383768 0 itasel1\[527\]
rlabel metal3 333942 357448 333942 357448 0 itasel1\[528\]
rlabel metal3 335230 358008 335230 358008 0 itasel1\[529\]
rlabel metal2 352744 71288 352744 71288 0 itasel1\[52\]
rlabel metal2 377608 372834 377608 372834 0 itasel1\[530\]
rlabel metal3 333942 359128 333942 359128 0 itasel1\[531\]
rlabel metal3 352086 359688 352086 359688 0 itasel1\[532\]
rlabel metal3 336910 360248 336910 360248 0 itasel1\[533\]
rlabel metal3 338590 360808 338590 360808 0 itasel1\[534\]
rlabel metal2 376936 428638 376936 428638 0 itasel1\[535\]
rlabel metal4 396760 392336 396760 392336 0 itasel1\[536\]
rlabel metal3 333270 362488 333270 362488 0 itasel1\[537\]
rlabel metal3 333214 363048 333214 363048 0 itasel1\[538\]
rlabel metal3 333550 363608 333550 363608 0 itasel1\[539\]
rlabel metal2 373898 70616 373898 70616 0 itasel1\[53\]
rlabel metal3 457478 404712 457478 404712 0 itasel1\[540\]
rlabel metal3 333158 364728 333158 364728 0 itasel1\[541\]
rlabel metal3 394030 365288 394030 365288 0 itasel1\[542\]
rlabel metal2 436184 428806 436184 428806 0 itasel1\[543\]
rlabel metal3 456526 406728 456526 406728 0 itasel1\[544\]
rlabel metal4 399000 384664 399000 384664 0 itasel1\[545\]
rlabel metal3 394646 367528 394646 367528 0 itasel1\[546\]
rlabel metal2 404040 397096 404040 397096 0 itasel1\[547\]
rlabel metal3 393638 368648 393638 368648 0 itasel1\[548\]
rlabel metal3 456582 404040 456582 404040 0 itasel1\[549\]
rlabel metal3 334502 69608 334502 69608 0 itasel1\[54\]
rlabel metal3 333606 369768 333606 369768 0 itasel1\[550\]
rlabel metal3 334054 370328 334054 370328 0 itasel1\[551\]
rlabel metal2 407400 398776 407400 398776 0 itasel1\[552\]
rlabel metal3 519470 402696 519470 402696 0 itasel1\[553\]
rlabel metal3 398230 372008 398230 372008 0 itasel1\[554\]
rlabel metal3 471954 408744 471954 408744 0 itasel1\[555\]
rlabel metal2 498232 379218 498232 379218 0 itasel1\[556\]
rlabel metal4 517496 387856 517496 387856 0 itasel1\[557\]
rlabel metal2 493528 379778 493528 379778 0 itasel1\[558\]
rlabel metal3 474474 406056 474474 406056 0 itasel1\[559\]
rlabel metal4 396760 60704 396760 60704 0 itasel1\[55\]
rlabel metal3 396550 375368 396550 375368 0 itasel1\[560\]
rlabel metal3 517944 405706 517944 405706 0 itasel1\[561\]
rlabel metal3 518574 408072 518574 408072 0 itasel1\[562\]
rlabel metal4 476280 381304 476280 381304 0 itasel1\[563\]
rlabel metal3 432726 377608 432726 377608 0 itasel1\[564\]
rlabel metal3 397390 378168 397390 378168 0 itasel1\[565\]
rlabel metal3 446110 378728 446110 378728 0 itasel1\[566\]
rlabel metal3 430990 379288 430990 379288 0 itasel1\[567\]
rlabel metal3 432670 379848 432670 379848 0 itasel1\[568\]
rlabel metal2 474712 403704 474712 403704 0 itasel1\[569\]
rlabel metal2 359576 72352 359576 72352 0 itasel1\[56\]
rlabel metal3 455798 380968 455798 380968 0 itasel1\[570\]
rlabel metal3 351638 381528 351638 381528 0 itasel1\[571\]
rlabel metal2 399224 404320 399224 404320 0 itasel1\[572\]
rlabel metal2 561624 428806 561624 428806 0 itasel1\[573\]
rlabel metal3 339878 383208 339878 383208 0 itasel1\[574\]
rlabel metal3 456638 383768 456638 383768 0 itasel1\[575\]
rlabel metal2 74760 469336 74760 469336 0 itasel1\[576\]
rlabel metal4 69832 456400 69832 456400 0 itasel1\[577\]
rlabel metal2 261688 427280 261688 427280 0 itasel1\[578\]
rlabel metal2 44968 447930 44968 447930 0 itasel1\[579\]
rlabel metal3 393960 53046 393960 53046 0 itasel1\[57\]
rlabel metal2 262920 459312 262920 459312 0 itasel1\[580\]
rlabel metal4 73080 453432 73080 453432 0 itasel1\[581\]
rlabel metal4 256200 430080 256200 430080 0 itasel1\[582\]
rlabel metal3 19026 477288 19026 477288 0 itasel1\[583\]
rlabel metal4 261240 428904 261240 428904 0 itasel1\[584\]
rlabel metal4 259560 430864 259560 430864 0 itasel1\[585\]
rlabel metal3 144032 452760 144032 452760 0 itasel1\[586\]
rlabel metal3 260554 421848 260554 421848 0 itasel1\[587\]
rlabel metal2 100856 450394 100856 450394 0 itasel1\[588\]
rlabel metal3 176232 447720 176232 447720 0 itasel1\[589\]
rlabel metal3 349482 52808 349482 52808 0 itasel1\[58\]
rlabel metal4 261352 434784 261352 434784 0 itasel1\[590\]
rlabel metal3 125398 474600 125398 474600 0 itasel1\[591\]
rlabel metal2 104888 499590 104888 499590 0 itasel1\[592\]
rlabel metal4 258216 439040 258216 439040 0 itasel1\[593\]
rlabel metal4 263368 430080 263368 430080 0 itasel1\[594\]
rlabel metal3 268072 426454 268072 426454 0 itasel1\[595\]
rlabel metal2 100856 499646 100856 499646 0 itasel1\[596\]
rlabel metal2 259672 463288 259672 463288 0 itasel1\[597\]
rlabel metal2 100184 499702 100184 499702 0 itasel1\[598\]
rlabel metal4 255640 430584 255640 430584 0 itasel1\[599\]
rlabel metal3 333662 72408 333662 72408 0 itasel1\[59\]
rlabel metal4 76440 67704 76440 67704 0 itasel1\[5\]
rlabel metal3 142450 476616 142450 476616 0 itasel1\[600\]
rlabel metal2 166264 499702 166264 499702 0 itasel1\[601\]
rlabel metal2 170968 499646 170968 499646 0 itasel1\[602\]
rlabel metal2 192360 464408 192360 464408 0 itasel1\[603\]
rlabel metal2 187544 464800 187544 464800 0 itasel1\[604\]
rlabel metal2 166264 449554 166264 449554 0 itasel1\[605\]
rlabel metal3 166712 449512 166712 449512 0 itasel1\[606\]
rlabel metal3 141512 475496 141512 475496 0 itasel1\[607\]
rlabel metal3 187502 482664 187502 482664 0 itasel1\[608\]
rlabel metal2 166936 445298 166936 445298 0 itasel1\[609\]
rlabel metal3 455896 47166 455896 47166 0 itasel1\[60\]
rlabel metal3 187446 478632 187446 478632 0 itasel1\[610\]
rlabel metal2 168952 445858 168952 445858 0 itasel1\[611\]
rlabel metal2 261352 468328 261352 468328 0 itasel1\[612\]
rlabel metal4 264600 456344 264600 456344 0 itasel1\[613\]
rlabel metal2 261464 467376 261464 467376 0 itasel1\[614\]
rlabel metal4 262920 459760 262920 459760 0 itasel1\[615\]
rlabel metal4 259672 460376 259672 460376 0 itasel1\[616\]
rlabel metal3 224056 450296 224056 450296 0 itasel1\[617\]
rlabel metal4 257880 456232 257880 456232 0 itasel1\[618\]
rlabel metal3 250390 477288 250390 477288 0 itasel1\[619\]
rlabel metal3 333214 73528 333214 73528 0 itasel1\[61\]
rlabel metal2 222824 498974 222824 498974 0 itasel1\[620\]
rlabel metal4 256536 457856 256536 457856 0 itasel1\[621\]
rlabel metal3 262752 441896 262752 441896 0 itasel1\[622\]
rlabel metal3 204666 481320 204666 481320 0 itasel1\[623\]
rlabel metal3 333550 415688 333550 415688 0 itasel1\[624\]
rlabel metal4 351960 432992 351960 432992 0 itasel1\[625\]
rlabel metal3 333718 416808 333718 416808 0 itasel1\[626\]
rlabel metal2 350280 431704 350280 431704 0 itasel1\[627\]
rlabel metal3 333606 417928 333606 417928 0 itasel1\[628\]
rlabel metal2 372904 499590 372904 499590 0 itasel1\[629\]
rlabel metal3 333270 74088 333270 74088 0 itasel1\[62\]
rlabel metal3 333662 419048 333662 419048 0 itasel1\[630\]
rlabel metal4 396872 461440 396872 461440 0 itasel1\[631\]
rlabel metal3 336070 420168 336070 420168 0 itasel1\[632\]
rlabel metal3 333550 420728 333550 420728 0 itasel1\[633\]
rlabel metal3 340270 421288 340270 421288 0 itasel1\[634\]
rlabel metal2 377608 450674 377608 450674 0 itasel1\[635\]
rlabel metal3 333214 422408 333214 422408 0 itasel1\[636\]
rlabel metal2 350392 461944 350392 461944 0 itasel1\[637\]
rlabel metal3 333214 423528 333214 423528 0 itasel1\[638\]
rlabel metal3 334390 424088 334390 424088 0 itasel1\[639\]
rlabel metal4 398104 71456 398104 71456 0 itasel1\[63\]
rlabel metal3 394478 424648 394478 424648 0 itasel1\[640\]
rlabel metal3 337134 425208 337134 425208 0 itasel1\[641\]
rlabel metal4 353640 436072 353640 436072 0 itasel1\[642\]
rlabel metal3 331912 426510 331912 426510 0 itasel1\[643\]
rlabel metal3 333886 426888 333886 426888 0 itasel1\[644\]
rlabel metal3 394534 427448 394534 427448 0 itasel1\[645\]
rlabel metal4 402360 450968 402360 450968 0 itasel1\[646\]
rlabel metal4 404040 453264 404040 453264 0 itasel1\[647\]
rlabel metal3 474474 479976 474474 479976 0 itasel1\[648\]
rlabel metal3 519582 479304 519582 479304 0 itasel1\[649\]
rlabel metal3 333158 75208 333158 75208 0 itasel1\[64\]
rlabel metal3 331912 430430 331912 430430 0 itasel1\[650\]
rlabel metal4 472136 482048 472136 482048 0 itasel1\[651\]
rlabel metal2 493528 498806 493528 498806 0 itasel1\[652\]
rlabel metal3 471954 477960 471954 477960 0 itasel1\[653\]
rlabel metal4 517496 456232 517496 456232 0 itasel1\[654\]
rlabel metal3 518574 483336 518574 483336 0 itasel1\[655\]
rlabel metal3 518630 476616 518630 476616 0 itasel1\[656\]
rlabel metal2 494200 453810 494200 453810 0 itasel1\[657\]
rlabel metal2 499576 452186 499576 452186 0 itasel1\[658\]
rlabel metal2 498904 499646 498904 499646 0 itasel1\[659\]
rlabel metal3 333214 75768 333214 75768 0 itasel1\[65\]
rlabel metal4 355320 441784 355320 441784 0 itasel1\[660\]
rlabel metal2 375480 443744 375480 443744 0 itasel1\[661\]
rlabel metal3 333886 436968 333886 436968 0 itasel1\[662\]
rlabel metal3 544488 497896 544488 497896 0 itasel1\[663\]
rlabel metal4 523320 458864 523320 458864 0 itasel1\[664\]
rlabel metal2 407512 469728 407512 469728 0 itasel1\[665\]
rlabel metal3 456694 439208 456694 439208 0 itasel1\[666\]
rlabel metal3 463736 449512 463736 449512 0 itasel1\[667\]
rlabel metal3 487368 446040 487368 446040 0 itasel1\[668\]
rlabel metal2 562296 499646 562296 499646 0 itasel1\[669\]
rlabel metal2 402360 75544 402360 75544 0 itasel1\[66\]
rlabel metal3 456638 441448 456638 441448 0 itasel1\[670\]
rlabel metal3 465472 444472 465472 444472 0 itasel1\[671\]
rlabel metal2 73080 539056 73080 539056 0 itasel1\[672\]
rlabel metal3 260904 480424 260904 480424 0 itasel1\[673\]
rlabel metal4 256312 498344 256312 498344 0 itasel1\[674\]
rlabel metal2 78120 537264 78120 537264 0 itasel1\[675\]
rlabel metal2 36582 569464 36582 569464 0 itasel1\[676\]
rlabel metal3 144984 523432 144984 523432 0 itasel1\[677\]
rlabel metal2 261688 494424 261688 494424 0 itasel1\[678\]
rlabel metal4 256200 503944 256200 503944 0 itasel1\[679\]
rlabel metal3 455896 52374 455896 52374 0 itasel1\[67\]
rlabel metal2 263816 479024 263816 479024 0 itasel1\[680\]
rlabel metal4 74760 527352 74760 527352 0 itasel1\[681\]
rlabel metal4 259560 504840 259560 504840 0 itasel1\[682\]
rlabel metal2 44296 570598 44296 570598 0 itasel1\[683\]
rlabel metal2 264712 496944 264712 496944 0 itasel1\[684\]
rlabel metal2 98840 526386 98840 526386 0 itasel1\[685\]
rlabel metal4 263144 500024 263144 500024 0 itasel1\[686\]
rlabel metal2 261240 526848 261240 526848 0 itasel1\[687\]
rlabel metal2 102200 518826 102200 518826 0 itasel1\[688\]
rlabel metal3 81130 544488 81130 544488 0 itasel1\[689\]
rlabel metal3 333550 77448 333550 77448 0 itasel1\[68\]
rlabel metal2 259784 500360 259784 500360 0 itasel1\[690\]
rlabel metal3 125622 552552 125622 552552 0 itasel1\[691\]
rlabel metal4 256536 503440 256536 503440 0 itasel1\[692\]
rlabel metal2 100184 570486 100184 570486 0 itasel1\[693\]
rlabel metal4 257992 500584 257992 500584 0 itasel1\[694\]
rlabel metal3 164136 520072 164136 520072 0 itasel1\[695\]
rlabel metal3 187446 549864 187446 549864 0 itasel1\[696\]
rlabel metal2 263032 529704 263032 529704 0 itasel1\[697\]
rlabel metal2 187320 534968 187320 534968 0 itasel1\[698\]
rlabel metal2 164248 570542 164248 570542 0 itasel1\[699\]
rlabel metal2 404040 53816 404040 53816 0 itasel1\[69\]
rlabel metal2 43848 70840 43848 70840 0 itasel1\[6\]
rlabel metal2 170296 570598 170296 570598 0 itasel1\[700\]
rlabel metal2 169624 516306 169624 516306 0 itasel1\[701\]
rlabel metal3 187502 551208 187502 551208 0 itasel1\[702\]
rlabel metal2 166390 569464 166390 569464 0 itasel1\[703\]
rlabel metal2 164248 526442 164248 526442 0 itasel1\[704\]
rlabel metal2 167608 517930 167608 517930 0 itasel1\[705\]
rlabel metal3 142562 544488 142562 544488 0 itasel1\[706\]
rlabel metal3 258818 493528 258818 493528 0 itasel1\[707\]
rlabel metal2 257992 532000 257992 532000 0 itasel1\[708\]
rlabel metal2 256200 533232 256200 533232 0 itasel1\[709\]
rlabel metal2 352072 52584 352072 52584 0 itasel1\[70\]
rlabel metal3 204610 543816 204610 543816 0 itasel1\[710\]
rlabel metal3 242704 568904 242704 568904 0 itasel1\[711\]
rlabel metal2 263144 533064 263144 533064 0 itasel1\[712\]
rlabel metal3 203672 544376 203672 544376 0 itasel1\[713\]
rlabel metal4 203168 544050 203168 544050 0 itasel1\[714\]
rlabel metal3 263424 500136 263424 500136 0 itasel1\[715\]
rlabel metal3 237328 525336 237328 525336 0 itasel1\[716\]
rlabel metal4 261240 521472 261240 521472 0 itasel1\[717\]
rlabel metal4 264600 523768 264600 523768 0 itasel1\[718\]
rlabel metal4 257880 524384 257880 524384 0 itasel1\[719\]
rlabel metal3 333942 79128 333942 79128 0 itasel1\[71\]
rlabel metal3 333886 473928 333886 473928 0 itasel1\[720\]
rlabel metal3 333774 474488 333774 474488 0 itasel1\[721\]
rlabel metal4 351960 498512 351960 498512 0 itasel1\[722\]
rlabel metal3 333774 475608 333774 475608 0 itasel1\[723\]
rlabel metal3 333550 476168 333550 476168 0 itasel1\[724\]
rlabel metal2 374248 570486 374248 570486 0 itasel1\[725\]
rlabel metal3 333662 477288 333662 477288 0 itasel1\[726\]
rlabel metal3 334614 477848 334614 477848 0 itasel1\[727\]
rlabel metal3 336910 478408 336910 478408 0 itasel1\[728\]
rlabel metal3 337022 478968 337022 478968 0 itasel1\[729\]
rlabel metal3 517944 47670 517944 47670 0 itasel1\[72\]
rlabel metal3 340270 479528 340270 479528 0 itasel1\[730\]
rlabel metal4 396872 527688 396872 527688 0 itasel1\[731\]
rlabel metal3 336126 480648 336126 480648 0 itasel1\[732\]
rlabel metal3 457366 545160 457366 545160 0 itasel1\[733\]
rlabel metal4 352184 494256 352184 494256 0 itasel1\[734\]
rlabel metal3 338758 482328 338758 482328 0 itasel1\[735\]
rlabel metal2 430808 570374 430808 570374 0 itasel1\[736\]
rlabel metal3 333718 483448 333718 483448 0 itasel1\[737\]
rlabel metal3 337078 484008 337078 484008 0 itasel1\[738\]
rlabel metal4 350616 495712 350616 495712 0 itasel1\[739\]
rlabel metal3 518686 48776 518686 48776 0 itasel1\[73\]
rlabel metal3 334446 485128 334446 485128 0 itasel1\[740\]
rlabel metal3 340438 485688 340438 485688 0 itasel1\[741\]
rlabel metal3 334558 486248 334558 486248 0 itasel1\[742\]
rlabel metal2 430136 515522 430136 515522 0 itasel1\[743\]
rlabel metal3 519638 551880 519638 551880 0 itasel1\[744\]
rlabel metal3 519470 549864 519470 549864 0 itasel1\[745\]
rlabel metal3 518574 544488 518574 544488 0 itasel1\[746\]
rlabel metal2 496216 570542 496216 570542 0 itasel1\[747\]
rlabel metal3 474474 553224 474474 553224 0 itasel1\[748\]
rlabel metal3 474656 547848 474656 547848 0 itasel1\[749\]
rlabel metal2 494200 74718 494200 74718 0 itasel1\[74\]
rlabel metal3 333606 490728 333606 490728 0 itasel1\[750\]
rlabel metal3 474530 546504 474530 546504 0 itasel1\[751\]
rlabel metal3 474586 550536 474586 550536 0 itasel1\[752\]
rlabel metal2 350616 500304 350616 500304 0 itasel1\[753\]
rlabel metal3 334390 492968 334390 492968 0 itasel1\[754\]
rlabel metal3 474698 545832 474698 545832 0 itasel1\[755\]
rlabel metal3 331912 494270 331912 494270 0 itasel1\[756\]
rlabel metal3 335342 494648 335342 494648 0 itasel1\[757\]
rlabel metal2 407400 533344 407400 533344 0 itasel1\[758\]
rlabel metal3 362950 495768 362950 495768 0 itasel1\[759\]
rlabel metal2 492562 71064 492562 71064 0 itasel1\[75\]
rlabel metal2 563640 516250 563640 516250 0 itasel1\[760\]
rlabel metal4 402360 501760 402360 501760 0 itasel1\[761\]
rlabel metal4 353752 507080 353752 507080 0 itasel1\[762\]
rlabel metal3 455798 498008 455798 498008 0 itasel1\[763\]
rlabel metal3 456638 498568 456638 498568 0 itasel1\[764\]
rlabel metal3 338758 499128 338758 499128 0 itasel1\[765\]
rlabel metal4 353864 504784 353864 504784 0 itasel1\[766\]
rlabel metal3 456694 500248 456694 500248 0 itasel1\[767\]
rlabel metal2 407400 55664 407400 55664 0 itasel1\[76\]
rlabel metal4 517608 67312 517608 67312 0 itasel1\[77\]
rlabel metal3 518630 48104 518630 48104 0 itasel1\[78\]
rlabel metal3 480368 29288 480368 29288 0 itasel1\[79\]
rlabel metal4 20664 68712 20664 68712 0 itasel1\[7\]
rlabel metal3 469434 52808 469434 52808 0 itasel1\[80\]
rlabel metal2 501592 72982 501592 72982 0 itasel1\[81\]
rlabel metal2 500920 72870 500920 72870 0 itasel1\[82\]
rlabel metal2 497560 73038 497560 73038 0 itasel1\[83\]
rlabel metal3 455854 86408 455854 86408 0 itasel1\[84\]
rlabel metal3 580734 54824 580734 54824 0 itasel1\[85\]
rlabel metal2 403256 84504 403256 84504 0 itasel1\[86\]
rlabel metal3 579880 46438 579880 46438 0 itasel1\[87\]
rlabel metal3 580678 55496 580678 55496 0 itasel1\[88\]
rlabel metal2 562296 72926 562296 72926 0 itasel1\[89\]
rlabel metal3 63294 51464 63294 51464 0 itasel1\[8\]
rlabel metal3 580622 47432 580622 47432 0 itasel1\[90\]
rlabel metal2 562296 27930 562296 27930 0 itasel1\[91\]
rlabel metal3 455798 90888 455798 90888 0 itasel1\[92\]
rlabel metal3 396942 91448 396942 91448 0 itasel1\[93\]
rlabel metal4 523320 72408 523320 72408 0 itasel1\[94\]
rlabel metal4 525000 71680 525000 71680 0 itasel1\[95\]
rlabel metal4 264824 127809 264824 127809 0 itasel1\[96\]
rlabel metal2 263816 125944 263816 125944 0 itasel1\[97\]
rlabel metal2 42952 143486 42952 143486 0 itasel1\[98\]
rlabel metal2 40936 142590 40936 142590 0 itasel1\[99\]
rlabel metal2 43624 28826 43624 28826 0 itasel1\[9\]
rlabel metal3 142562 56168 142562 56168 0 wb_clk_i
<< properties >>
string FIXED_BBOX 0 0 596040 596040
<< end >>
