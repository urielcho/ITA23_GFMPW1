magic
tech gf180mcuD
magscale 1 5
timestamp 1699641779
<< metal1 >>
rect 672 19221 20328 19238
rect 672 19195 2239 19221
rect 2265 19195 2291 19221
rect 2317 19195 2343 19221
rect 2369 19195 17599 19221
rect 17625 19195 17651 19221
rect 17677 19195 17703 19221
rect 17729 19195 20328 19221
rect 672 19178 20328 19195
rect 13119 19137 13145 19143
rect 13119 19105 13145 19111
rect 9081 19055 9087 19081
rect 9113 19055 9119 19081
rect 11097 19055 11103 19081
rect 11129 19055 11135 19081
rect 9865 18999 9871 19025
rect 9897 18999 9903 19025
rect 11769 18999 11775 19025
rect 11801 18999 11807 19025
rect 12833 18999 12839 19025
rect 12865 18999 12871 19025
rect 672 18829 20328 18846
rect 672 18803 9919 18829
rect 9945 18803 9971 18829
rect 9997 18803 10023 18829
rect 10049 18803 20328 18829
rect 672 18786 20328 18803
rect 9199 18745 9225 18751
rect 9199 18713 9225 18719
rect 11383 18745 11409 18751
rect 11383 18713 11409 18719
rect 8801 18607 8807 18633
rect 8833 18607 8839 18633
rect 10929 18607 10935 18633
rect 10961 18607 10967 18633
rect 672 18437 20328 18454
rect 672 18411 2239 18437
rect 2265 18411 2291 18437
rect 2317 18411 2343 18437
rect 2369 18411 17599 18437
rect 17625 18411 17651 18437
rect 17677 18411 17703 18437
rect 17729 18411 20328 18437
rect 672 18394 20328 18411
rect 672 18045 20328 18062
rect 672 18019 9919 18045
rect 9945 18019 9971 18045
rect 9997 18019 10023 18045
rect 10049 18019 20328 18045
rect 672 18002 20328 18019
rect 672 17653 20328 17670
rect 672 17627 2239 17653
rect 2265 17627 2291 17653
rect 2317 17627 2343 17653
rect 2369 17627 17599 17653
rect 17625 17627 17651 17653
rect 17677 17627 17703 17653
rect 17729 17627 20328 17653
rect 672 17610 20328 17627
rect 672 17261 20328 17278
rect 672 17235 9919 17261
rect 9945 17235 9971 17261
rect 9997 17235 10023 17261
rect 10049 17235 20328 17261
rect 672 17218 20328 17235
rect 672 16869 20328 16886
rect 672 16843 2239 16869
rect 2265 16843 2291 16869
rect 2317 16843 2343 16869
rect 2369 16843 17599 16869
rect 17625 16843 17651 16869
rect 17677 16843 17703 16869
rect 17729 16843 20328 16869
rect 672 16826 20328 16843
rect 672 16477 20328 16494
rect 672 16451 9919 16477
rect 9945 16451 9971 16477
rect 9997 16451 10023 16477
rect 10049 16451 20328 16477
rect 672 16434 20328 16451
rect 672 16085 20328 16102
rect 672 16059 2239 16085
rect 2265 16059 2291 16085
rect 2317 16059 2343 16085
rect 2369 16059 17599 16085
rect 17625 16059 17651 16085
rect 17677 16059 17703 16085
rect 17729 16059 20328 16085
rect 672 16042 20328 16059
rect 672 15693 20328 15710
rect 672 15667 9919 15693
rect 9945 15667 9971 15693
rect 9997 15667 10023 15693
rect 10049 15667 20328 15693
rect 672 15650 20328 15667
rect 672 15301 20328 15318
rect 672 15275 2239 15301
rect 2265 15275 2291 15301
rect 2317 15275 2343 15301
rect 2369 15275 17599 15301
rect 17625 15275 17651 15301
rect 17677 15275 17703 15301
rect 17729 15275 20328 15301
rect 672 15258 20328 15275
rect 672 14909 20328 14926
rect 672 14883 9919 14909
rect 9945 14883 9971 14909
rect 9997 14883 10023 14909
rect 10049 14883 20328 14909
rect 672 14866 20328 14883
rect 672 14517 20328 14534
rect 672 14491 2239 14517
rect 2265 14491 2291 14517
rect 2317 14491 2343 14517
rect 2369 14491 17599 14517
rect 17625 14491 17651 14517
rect 17677 14491 17703 14517
rect 17729 14491 20328 14517
rect 672 14474 20328 14491
rect 672 14125 20328 14142
rect 672 14099 9919 14125
rect 9945 14099 9971 14125
rect 9997 14099 10023 14125
rect 10049 14099 20328 14125
rect 672 14082 20328 14099
rect 18825 13903 18831 13929
rect 18857 13903 18863 13929
rect 19945 13847 19951 13873
rect 19977 13847 19983 13873
rect 672 13733 20328 13750
rect 672 13707 2239 13733
rect 2265 13707 2291 13733
rect 2317 13707 2343 13733
rect 2369 13707 17599 13733
rect 17625 13707 17651 13733
rect 17677 13707 17703 13733
rect 17729 13707 20328 13733
rect 672 13690 20328 13707
rect 20007 13593 20033 13599
rect 8577 13567 8583 13593
rect 8609 13567 8615 13593
rect 20007 13561 20033 13567
rect 10655 13537 10681 13543
rect 7177 13511 7183 13537
rect 7209 13511 7215 13537
rect 10655 13505 10681 13511
rect 10991 13537 11017 13543
rect 13449 13511 13455 13537
rect 13481 13511 13487 13537
rect 18937 13511 18943 13537
rect 18969 13511 18975 13537
rect 10991 13505 11017 13511
rect 8695 13481 8721 13487
rect 7513 13455 7519 13481
rect 7545 13455 7551 13481
rect 8695 13449 8721 13455
rect 8807 13481 8833 13487
rect 8807 13449 8833 13455
rect 8863 13481 8889 13487
rect 8863 13449 8889 13455
rect 9087 13481 9113 13487
rect 9087 13449 9113 13455
rect 12559 13481 12585 13487
rect 12559 13449 12585 13455
rect 12615 13481 12641 13487
rect 13561 13455 13567 13481
rect 13593 13455 13599 13481
rect 12615 13449 12641 13455
rect 10711 13425 10737 13431
rect 10711 13393 10737 13399
rect 10767 13425 10793 13431
rect 10767 13393 10793 13399
rect 12727 13425 12753 13431
rect 12727 13393 12753 13399
rect 672 13341 20328 13358
rect 672 13315 9919 13341
rect 9945 13315 9971 13341
rect 9997 13315 10023 13341
rect 10049 13315 20328 13341
rect 672 13298 20328 13315
rect 8079 13257 8105 13263
rect 11383 13257 11409 13263
rect 9305 13231 9311 13257
rect 9337 13231 9343 13257
rect 8079 13225 8105 13231
rect 11383 13225 11409 13231
rect 11495 13257 11521 13263
rect 11495 13225 11521 13231
rect 11551 13201 11577 13207
rect 10201 13175 10207 13201
rect 10233 13175 10239 13201
rect 11551 13169 11577 13175
rect 12279 13201 12305 13207
rect 12279 13169 12305 13175
rect 12335 13201 12361 13207
rect 12335 13169 12361 13175
rect 8023 13145 8049 13151
rect 8023 13113 8049 13119
rect 8191 13145 8217 13151
rect 8191 13113 8217 13119
rect 9479 13145 9505 13151
rect 11831 13145 11857 13151
rect 9865 13119 9871 13145
rect 9897 13119 9903 13145
rect 9479 13113 9505 13119
rect 11831 13113 11857 13119
rect 12167 13145 12193 13151
rect 12609 13119 12615 13145
rect 12641 13119 12647 13145
rect 18825 13119 18831 13145
rect 18857 13119 18863 13145
rect 12167 13113 12193 13119
rect 14463 13089 14489 13095
rect 11265 13063 11271 13089
rect 11297 13063 11303 13089
rect 13001 13063 13007 13089
rect 13033 13063 13039 13089
rect 14121 13063 14127 13089
rect 14153 13063 14159 13089
rect 14463 13057 14489 13063
rect 20007 13033 20033 13039
rect 20007 13001 20033 13007
rect 672 12949 20328 12966
rect 672 12923 2239 12949
rect 2265 12923 2291 12949
rect 2317 12923 2343 12949
rect 2369 12923 17599 12949
rect 17625 12923 17651 12949
rect 17677 12923 17703 12949
rect 17729 12923 20328 12949
rect 672 12906 20328 12923
rect 13175 12809 13201 12815
rect 9249 12783 9255 12809
rect 9281 12783 9287 12809
rect 12945 12783 12951 12809
rect 12977 12783 12983 12809
rect 13175 12777 13201 12783
rect 9535 12753 9561 12759
rect 7793 12727 7799 12753
rect 7825 12727 7831 12753
rect 9535 12721 9561 12727
rect 10431 12753 10457 12759
rect 10431 12721 10457 12727
rect 10599 12753 10625 12759
rect 11545 12727 11551 12753
rect 11577 12727 11583 12753
rect 13449 12727 13455 12753
rect 13481 12727 13487 12753
rect 10599 12721 10625 12727
rect 9479 12697 9505 12703
rect 8185 12671 8191 12697
rect 8217 12671 8223 12697
rect 9479 12665 9505 12671
rect 10263 12697 10289 12703
rect 10263 12665 10289 12671
rect 10319 12697 10345 12703
rect 11881 12671 11887 12697
rect 11913 12671 11919 12697
rect 13561 12671 13567 12697
rect 13593 12671 13599 12697
rect 10319 12665 10345 12671
rect 9367 12641 9393 12647
rect 9367 12609 9393 12615
rect 9759 12641 9785 12647
rect 9759 12609 9785 12615
rect 10823 12641 10849 12647
rect 10823 12609 10849 12615
rect 10879 12641 10905 12647
rect 10879 12609 10905 12615
rect 10935 12641 10961 12647
rect 10935 12609 10961 12615
rect 672 12557 20328 12574
rect 672 12531 9919 12557
rect 9945 12531 9971 12557
rect 9997 12531 10023 12557
rect 10049 12531 20328 12557
rect 672 12514 20328 12531
rect 6007 12473 6033 12479
rect 6007 12441 6033 12447
rect 8415 12473 8441 12479
rect 8415 12441 8441 12447
rect 8751 12473 8777 12479
rect 8751 12441 8777 12447
rect 9423 12473 9449 12479
rect 9423 12441 9449 12447
rect 11607 12473 11633 12479
rect 11607 12441 11633 12447
rect 11663 12473 11689 12479
rect 11663 12441 11689 12447
rect 12783 12473 12809 12479
rect 12783 12441 12809 12447
rect 7967 12417 7993 12423
rect 7967 12385 7993 12391
rect 9199 12417 9225 12423
rect 12615 12417 12641 12423
rect 9977 12391 9983 12417
rect 10009 12391 10015 12417
rect 9199 12385 9225 12391
rect 12615 12385 12641 12391
rect 12671 12417 12697 12423
rect 12671 12385 12697 12391
rect 20119 12417 20145 12423
rect 20119 12385 20145 12391
rect 8247 12361 8273 12367
rect 5889 12335 5895 12361
rect 5921 12335 5927 12361
rect 6169 12335 6175 12361
rect 6201 12335 6207 12361
rect 6561 12335 6567 12361
rect 6593 12335 6599 12361
rect 8073 12335 8079 12361
rect 8105 12335 8111 12361
rect 8247 12329 8273 12335
rect 9143 12361 9169 12367
rect 11719 12361 11745 12367
rect 9641 12335 9647 12361
rect 9673 12335 9679 12361
rect 9143 12329 9169 12335
rect 11719 12329 11745 12335
rect 11943 12361 11969 12367
rect 11943 12329 11969 12335
rect 8807 12305 8833 12311
rect 7625 12279 7631 12305
rect 7657 12279 7663 12305
rect 8017 12279 8023 12305
rect 8049 12279 8055 12305
rect 11041 12279 11047 12305
rect 11073 12279 11079 12305
rect 8807 12273 8833 12279
rect 8919 12249 8945 12255
rect 8919 12217 8945 12223
rect 672 12165 20328 12182
rect 672 12139 2239 12165
rect 2265 12139 2291 12165
rect 2317 12139 2343 12165
rect 2369 12139 17599 12165
rect 17625 12139 17651 12165
rect 17677 12139 17703 12165
rect 17729 12139 20328 12165
rect 672 12122 20328 12139
rect 10649 12055 10655 12081
rect 10681 12055 10687 12081
rect 7743 12025 7769 12031
rect 7905 11999 7911 12025
rect 7937 11999 7943 12025
rect 7743 11993 7769 11999
rect 10823 11969 10849 11975
rect 10823 11937 10849 11943
rect 10935 11969 10961 11975
rect 10935 11937 10961 11943
rect 672 11773 20328 11790
rect 672 11747 9919 11773
rect 9945 11747 9971 11773
rect 9997 11747 10023 11773
rect 10049 11747 20328 11773
rect 672 11730 20328 11747
rect 9087 11689 9113 11695
rect 9087 11657 9113 11663
rect 8079 11633 8105 11639
rect 8695 11633 8721 11639
rect 12895 11633 12921 11639
rect 6225 11607 6231 11633
rect 6257 11607 6263 11633
rect 8241 11607 8247 11633
rect 8273 11607 8279 11633
rect 10089 11607 10095 11633
rect 10121 11607 10127 11633
rect 8079 11601 8105 11607
rect 8695 11601 8721 11607
rect 12895 11601 12921 11607
rect 7911 11577 7937 11583
rect 12671 11577 12697 11583
rect 13735 11577 13761 11583
rect 5889 11551 5895 11577
rect 5921 11551 5927 11577
rect 8353 11551 8359 11577
rect 8385 11551 8391 11577
rect 8801 11551 8807 11577
rect 8833 11551 8839 11577
rect 8969 11551 8975 11577
rect 9001 11551 9007 11577
rect 10201 11551 10207 11577
rect 10233 11551 10239 11577
rect 10649 11551 10655 11577
rect 10681 11551 10687 11577
rect 12329 11551 12335 11577
rect 12361 11551 12367 11577
rect 13057 11551 13063 11577
rect 13089 11551 13095 11577
rect 13225 11551 13231 11577
rect 13257 11551 13263 11577
rect 7911 11545 7937 11551
rect 12671 11545 12697 11551
rect 13735 11545 13761 11551
rect 13847 11577 13873 11583
rect 13847 11545 13873 11551
rect 13959 11577 13985 11583
rect 13959 11545 13985 11551
rect 14015 11577 14041 11583
rect 14015 11545 14041 11551
rect 7519 11521 7545 11527
rect 13343 11521 13369 11527
rect 7289 11495 7295 11521
rect 7321 11495 7327 11521
rect 10481 11495 10487 11521
rect 10513 11495 10519 11521
rect 10873 11495 10879 11521
rect 10905 11495 10911 11521
rect 11937 11495 11943 11521
rect 11969 11495 11975 11521
rect 7519 11489 7545 11495
rect 13343 11489 13369 11495
rect 13063 11465 13089 11471
rect 8969 11439 8975 11465
rect 9001 11439 9007 11465
rect 13063 11433 13089 11439
rect 13399 11465 13425 11471
rect 13399 11433 13425 11439
rect 672 11381 20328 11398
rect 672 11355 2239 11381
rect 2265 11355 2291 11381
rect 2317 11355 2343 11381
rect 2369 11355 17599 11381
rect 17625 11355 17651 11381
rect 17677 11355 17703 11381
rect 17729 11355 20328 11381
rect 672 11338 20328 11355
rect 11831 11297 11857 11303
rect 10313 11271 10319 11297
rect 10345 11271 10351 11297
rect 11831 11265 11857 11271
rect 10767 11241 10793 11247
rect 10767 11209 10793 11215
rect 11551 11241 11577 11247
rect 14631 11241 14657 11247
rect 13225 11215 13231 11241
rect 13257 11215 13263 11241
rect 14289 11215 14295 11241
rect 14321 11215 14327 11241
rect 11551 11209 11577 11215
rect 14631 11209 14657 11215
rect 20007 11241 20033 11247
rect 20007 11209 20033 11215
rect 7463 11185 7489 11191
rect 7463 11153 7489 11159
rect 7743 11185 7769 11191
rect 7743 11153 7769 11159
rect 7855 11185 7881 11191
rect 7855 11153 7881 11159
rect 8079 11185 8105 11191
rect 8079 11153 8105 11159
rect 8135 11185 8161 11191
rect 9199 11185 9225 11191
rect 10655 11185 10681 11191
rect 8409 11159 8415 11185
rect 8441 11159 8447 11185
rect 8745 11159 8751 11185
rect 8777 11159 8783 11185
rect 9417 11159 9423 11185
rect 9449 11159 9455 11185
rect 10089 11159 10095 11185
rect 10121 11159 10127 11185
rect 10313 11159 10319 11185
rect 10345 11159 10351 11185
rect 8135 11153 8161 11159
rect 9199 11153 9225 11159
rect 10655 11153 10681 11159
rect 11103 11185 11129 11191
rect 11103 11153 11129 11159
rect 11607 11185 11633 11191
rect 12833 11159 12839 11185
rect 12865 11159 12871 11185
rect 18825 11159 18831 11185
rect 18857 11159 18863 11185
rect 11607 11153 11633 11159
rect 9143 11129 9169 11135
rect 9143 11097 9169 11103
rect 11159 11129 11185 11135
rect 11159 11097 11185 11103
rect 11775 11129 11801 11135
rect 11775 11097 11801 11103
rect 8023 11073 8049 11079
rect 8023 11041 8049 11047
rect 8527 11073 8553 11079
rect 11383 11073 11409 11079
rect 8857 11047 8863 11073
rect 8889 11047 8895 11073
rect 9529 11047 9535 11073
rect 9561 11047 9567 11073
rect 10929 11047 10935 11073
rect 10961 11047 10967 11073
rect 8527 11041 8553 11047
rect 11383 11041 11409 11047
rect 11495 11073 11521 11079
rect 11495 11041 11521 11047
rect 11831 11073 11857 11079
rect 11831 11041 11857 11047
rect 672 10989 20328 11006
rect 672 10963 9919 10989
rect 9945 10963 9971 10989
rect 9997 10963 10023 10989
rect 10049 10963 20328 10989
rect 672 10946 20328 10963
rect 7407 10905 7433 10911
rect 7407 10873 7433 10879
rect 8079 10905 8105 10911
rect 8079 10873 8105 10879
rect 10935 10905 10961 10911
rect 14631 10905 14657 10911
rect 11713 10879 11719 10905
rect 11745 10879 11751 10905
rect 10935 10873 10961 10879
rect 14631 10873 14657 10879
rect 8689 10823 8695 10849
rect 8721 10823 8727 10849
rect 9305 10823 9311 10849
rect 9337 10823 9343 10849
rect 9809 10823 9815 10849
rect 9841 10823 9847 10849
rect 13337 10823 13343 10849
rect 13369 10823 13375 10849
rect 8023 10793 8049 10799
rect 5777 10767 5783 10793
rect 5809 10767 5815 10793
rect 8023 10761 8049 10767
rect 8247 10793 8273 10799
rect 8247 10761 8273 10767
rect 8863 10793 8889 10799
rect 10599 10793 10625 10799
rect 9249 10767 9255 10793
rect 9281 10767 9287 10793
rect 8863 10761 8889 10767
rect 10599 10761 10625 10767
rect 10823 10793 10849 10799
rect 10823 10761 10849 10767
rect 11159 10793 11185 10799
rect 11159 10761 11185 10767
rect 11383 10793 11409 10799
rect 11383 10761 11409 10767
rect 11439 10793 11465 10799
rect 11439 10761 11465 10767
rect 11495 10793 11521 10799
rect 12945 10767 12951 10793
rect 12977 10767 12983 10793
rect 18825 10767 18831 10793
rect 18857 10767 18863 10793
rect 11495 10761 11521 10767
rect 10879 10737 10905 10743
rect 20007 10737 20033 10743
rect 6113 10711 6119 10737
rect 6145 10711 6151 10737
rect 7177 10711 7183 10737
rect 7209 10711 7215 10737
rect 10649 10711 10655 10737
rect 10681 10711 10687 10737
rect 14401 10711 14407 10737
rect 14433 10711 14439 10737
rect 10879 10705 10905 10711
rect 20007 10705 20033 10711
rect 672 10597 20328 10614
rect 672 10571 2239 10597
rect 2265 10571 2291 10597
rect 2317 10571 2343 10597
rect 2369 10571 17599 10597
rect 17625 10571 17651 10597
rect 17677 10571 17703 10597
rect 17729 10571 20328 10597
rect 672 10554 20328 10571
rect 9143 10513 9169 10519
rect 9143 10481 9169 10487
rect 9311 10513 9337 10519
rect 9311 10481 9337 10487
rect 10767 10513 10793 10519
rect 10767 10481 10793 10487
rect 967 10457 993 10463
rect 9031 10457 9057 10463
rect 8017 10431 8023 10457
rect 8049 10431 8055 10457
rect 967 10425 993 10431
rect 9031 10425 9057 10431
rect 9759 10457 9785 10463
rect 12945 10431 12951 10457
rect 12977 10431 12983 10457
rect 9759 10425 9785 10431
rect 9479 10401 9505 10407
rect 2137 10375 2143 10401
rect 2169 10375 2175 10401
rect 8129 10375 8135 10401
rect 8161 10375 8167 10401
rect 9479 10369 9505 10375
rect 10095 10401 10121 10407
rect 10095 10369 10121 10375
rect 10991 10401 11017 10407
rect 11769 10375 11775 10401
rect 11801 10375 11807 10401
rect 10991 10369 11017 10375
rect 7799 10345 7825 10351
rect 7799 10313 7825 10319
rect 10823 10345 10849 10351
rect 10823 10313 10849 10319
rect 11327 10345 11353 10351
rect 11327 10313 11353 10319
rect 10767 10289 10793 10295
rect 10257 10263 10263 10289
rect 10289 10263 10295 10289
rect 10767 10257 10793 10263
rect 11159 10289 11185 10295
rect 11159 10257 11185 10263
rect 11383 10289 11409 10295
rect 11383 10257 11409 10263
rect 11495 10289 11521 10295
rect 11495 10257 11521 10263
rect 672 10205 20328 10222
rect 672 10179 9919 10205
rect 9945 10179 9971 10205
rect 9997 10179 10023 10205
rect 10049 10179 20328 10205
rect 672 10162 20328 10179
rect 8751 10121 8777 10127
rect 8751 10089 8777 10095
rect 9087 10121 9113 10127
rect 9087 10089 9113 10095
rect 7519 10065 7545 10071
rect 7345 10039 7351 10065
rect 7377 10039 7383 10065
rect 7519 10033 7545 10039
rect 7799 10065 7825 10071
rect 7799 10033 7825 10039
rect 7911 10065 7937 10071
rect 7911 10033 7937 10039
rect 8359 10065 8385 10071
rect 8359 10033 8385 10039
rect 8863 10065 8889 10071
rect 13567 10065 13593 10071
rect 11713 10039 11719 10065
rect 11745 10039 11751 10065
rect 8863 10033 8889 10039
rect 13567 10033 13593 10039
rect 13791 10065 13817 10071
rect 13791 10033 13817 10039
rect 13903 10065 13929 10071
rect 13903 10033 13929 10039
rect 14015 10065 14041 10071
rect 14015 10033 14041 10039
rect 7239 10009 7265 10015
rect 6785 9983 6791 10009
rect 6817 9983 6823 10009
rect 7239 9977 7265 9983
rect 7967 10009 7993 10015
rect 7967 9977 7993 9983
rect 9031 10009 9057 10015
rect 9031 9977 9057 9983
rect 9199 10009 9225 10015
rect 13399 10009 13425 10015
rect 9697 9983 9703 10009
rect 9729 9983 9735 10009
rect 9199 9977 9225 9983
rect 13399 9977 13425 9983
rect 13679 10009 13705 10015
rect 13679 9977 13705 9983
rect 7015 9953 7041 9959
rect 9535 9953 9561 9959
rect 5329 9927 5335 9953
rect 5361 9927 5367 9953
rect 6393 9927 6399 9953
rect 6425 9927 6431 9953
rect 7177 9927 7183 9953
rect 7209 9927 7215 9953
rect 7015 9921 7041 9927
rect 9535 9921 9561 9927
rect 7631 9897 7657 9903
rect 7631 9865 7657 9871
rect 7687 9897 7713 9903
rect 7687 9865 7713 9871
rect 8415 9897 8441 9903
rect 8415 9865 8441 9871
rect 8695 9897 8721 9903
rect 8695 9865 8721 9871
rect 672 9813 20328 9830
rect 672 9787 2239 9813
rect 2265 9787 2291 9813
rect 2317 9787 2343 9813
rect 2369 9787 17599 9813
rect 17625 9787 17651 9813
rect 17677 9787 17703 9813
rect 17729 9787 20328 9813
rect 672 9770 20328 9787
rect 6175 9729 6201 9735
rect 6175 9697 6201 9703
rect 6791 9729 6817 9735
rect 6791 9697 6817 9703
rect 13735 9729 13761 9735
rect 13735 9697 13761 9703
rect 6231 9673 6257 9679
rect 6231 9641 6257 9647
rect 13119 9673 13145 9679
rect 13119 9641 13145 9647
rect 13959 9673 13985 9679
rect 13959 9641 13985 9647
rect 20007 9673 20033 9679
rect 20007 9641 20033 9647
rect 7575 9617 7601 9623
rect 11327 9617 11353 9623
rect 12615 9617 12641 9623
rect 10033 9591 10039 9617
rect 10065 9591 10071 9617
rect 11601 9591 11607 9617
rect 11633 9591 11639 9617
rect 7575 9585 7601 9591
rect 11327 9585 11353 9591
rect 12615 9585 12641 9591
rect 14127 9617 14153 9623
rect 18825 9591 18831 9617
rect 18857 9591 18863 9617
rect 14127 9585 14153 9591
rect 6847 9561 6873 9567
rect 11943 9561 11969 9567
rect 13007 9561 13033 9567
rect 8465 9535 8471 9561
rect 8497 9535 8503 9561
rect 10817 9535 10823 9561
rect 10849 9535 10855 9561
rect 12777 9535 12783 9561
rect 12809 9535 12815 9561
rect 6847 9529 6873 9535
rect 11943 9529 11969 9535
rect 13007 9529 13033 9535
rect 13903 9561 13929 9567
rect 13903 9529 13929 9535
rect 14071 9561 14097 9567
rect 14071 9529 14097 9535
rect 6791 9505 6817 9511
rect 10655 9505 10681 9511
rect 11775 9505 11801 9511
rect 7401 9479 7407 9505
rect 7433 9479 7439 9505
rect 11153 9479 11159 9505
rect 11185 9479 11191 9505
rect 11489 9479 11495 9505
rect 11521 9479 11527 9505
rect 6791 9473 6817 9479
rect 10655 9473 10681 9479
rect 11775 9473 11801 9479
rect 11887 9505 11913 9511
rect 11887 9473 11913 9479
rect 13063 9505 13089 9511
rect 13063 9473 13089 9479
rect 13623 9505 13649 9511
rect 13623 9473 13649 9479
rect 13679 9505 13705 9511
rect 13679 9473 13705 9479
rect 672 9421 20328 9438
rect 672 9395 9919 9421
rect 9945 9395 9971 9421
rect 9997 9395 10023 9421
rect 10049 9395 20328 9421
rect 672 9378 20328 9395
rect 7855 9337 7881 9343
rect 7855 9305 7881 9311
rect 7967 9337 7993 9343
rect 7967 9305 7993 9311
rect 8359 9337 8385 9343
rect 8359 9305 8385 9311
rect 9199 9337 9225 9343
rect 9199 9305 9225 9311
rect 9591 9337 9617 9343
rect 9591 9305 9617 9311
rect 9983 9337 10009 9343
rect 9983 9305 10009 9311
rect 8079 9281 8105 9287
rect 8079 9249 8105 9255
rect 8303 9281 8329 9287
rect 8303 9249 8329 9255
rect 9255 9281 9281 9287
rect 9927 9281 9953 9287
rect 9753 9255 9759 9281
rect 9785 9255 9791 9281
rect 9255 9249 9281 9255
rect 9927 9249 9953 9255
rect 10263 9281 10289 9287
rect 10263 9249 10289 9255
rect 10319 9281 10345 9287
rect 10319 9249 10345 9255
rect 11999 9281 12025 9287
rect 13729 9255 13735 9281
rect 13761 9255 13767 9281
rect 11999 9249 12025 9255
rect 6791 9225 6817 9231
rect 2137 9199 2143 9225
rect 2169 9199 2175 9225
rect 6225 9199 6231 9225
rect 6257 9199 6263 9225
rect 6617 9199 6623 9225
rect 6649 9199 6655 9225
rect 6791 9193 6817 9199
rect 6847 9225 6873 9231
rect 6847 9193 6873 9199
rect 6903 9225 6929 9231
rect 6903 9193 6929 9199
rect 7071 9225 7097 9231
rect 7071 9193 7097 9199
rect 7799 9225 7825 9231
rect 7799 9193 7825 9199
rect 8639 9225 8665 9231
rect 8639 9193 8665 9199
rect 8807 9225 8833 9231
rect 8807 9193 8833 9199
rect 8975 9225 9001 9231
rect 8975 9193 9001 9199
rect 10431 9225 10457 9231
rect 10431 9193 10457 9199
rect 10655 9225 10681 9231
rect 10655 9193 10681 9199
rect 10767 9225 10793 9231
rect 10767 9193 10793 9199
rect 11215 9225 11241 9231
rect 11215 9193 11241 9199
rect 11271 9225 11297 9231
rect 11271 9193 11297 9199
rect 11495 9225 11521 9231
rect 11495 9193 11521 9199
rect 11607 9225 11633 9231
rect 11607 9193 11633 9199
rect 11775 9225 11801 9231
rect 11775 9193 11801 9199
rect 12111 9225 12137 9231
rect 15023 9225 15049 9231
rect 13337 9199 13343 9225
rect 13369 9199 13375 9225
rect 18825 9199 18831 9225
rect 18857 9199 18863 9225
rect 12111 9193 12137 9199
rect 15023 9193 15049 9199
rect 7295 9169 7321 9175
rect 5161 9143 5167 9169
rect 5193 9143 5199 9169
rect 7295 9137 7321 9143
rect 8751 9169 8777 9175
rect 8751 9137 8777 9143
rect 11103 9169 11129 9175
rect 11103 9137 11129 9143
rect 11887 9169 11913 9175
rect 14793 9143 14799 9169
rect 14825 9143 14831 9169
rect 11887 9137 11913 9143
rect 967 9113 993 9119
rect 967 9081 993 9087
rect 8359 9113 8385 9119
rect 8359 9081 8385 9087
rect 9199 9113 9225 9119
rect 9199 9081 9225 9087
rect 9983 9113 10009 9119
rect 9983 9081 10009 9087
rect 10935 9113 10961 9119
rect 10935 9081 10961 9087
rect 20007 9113 20033 9119
rect 20007 9081 20033 9087
rect 672 9029 20328 9046
rect 672 9003 2239 9029
rect 2265 9003 2291 9029
rect 2317 9003 2343 9029
rect 2369 9003 17599 9029
rect 17625 9003 17651 9029
rect 17677 9003 17703 9029
rect 17729 9003 20328 9029
rect 672 8986 20328 9003
rect 6791 8945 6817 8951
rect 6791 8913 6817 8919
rect 9143 8945 9169 8951
rect 9143 8913 9169 8919
rect 13287 8945 13313 8951
rect 13287 8913 13313 8919
rect 14071 8945 14097 8951
rect 14071 8913 14097 8919
rect 9927 8889 9953 8895
rect 13175 8889 13201 8895
rect 11937 8863 11943 8889
rect 11969 8863 11975 8889
rect 13001 8863 13007 8889
rect 13033 8863 13039 8889
rect 9927 8857 9953 8863
rect 13175 8857 13201 8863
rect 20007 8889 20033 8895
rect 20007 8857 20033 8863
rect 8583 8833 8609 8839
rect 8583 8801 8609 8807
rect 9535 8833 9561 8839
rect 9535 8801 9561 8807
rect 9983 8833 10009 8839
rect 14239 8833 14265 8839
rect 11601 8807 11607 8833
rect 11633 8807 11639 8833
rect 13785 8807 13791 8833
rect 13817 8807 13823 8833
rect 9983 8801 10009 8807
rect 14239 8801 14265 8807
rect 14575 8833 14601 8839
rect 14575 8801 14601 8807
rect 14687 8833 14713 8839
rect 15129 8807 15135 8833
rect 15161 8807 15167 8833
rect 18825 8807 18831 8833
rect 18857 8807 18863 8833
rect 14687 8801 14713 8807
rect 6791 8777 6817 8783
rect 6791 8745 6817 8751
rect 6847 8777 6873 8783
rect 6847 8745 6873 8751
rect 8303 8777 8329 8783
rect 8303 8745 8329 8751
rect 9031 8777 9057 8783
rect 9759 8777 9785 8783
rect 9361 8751 9367 8777
rect 9393 8751 9399 8777
rect 13673 8751 13679 8777
rect 13705 8751 13711 8777
rect 14849 8751 14855 8777
rect 14881 8751 14887 8777
rect 9031 8745 9057 8751
rect 9759 8745 9785 8751
rect 8247 8721 8273 8727
rect 8247 8689 8273 8695
rect 8415 8721 8441 8727
rect 8415 8689 8441 8695
rect 9087 8721 9113 8727
rect 9087 8689 9113 8695
rect 9871 8721 9897 8727
rect 15023 8721 15049 8727
rect 13449 8695 13455 8721
rect 13481 8695 13487 8721
rect 9871 8689 9897 8695
rect 15023 8689 15049 8695
rect 672 8637 20328 8654
rect 672 8611 9919 8637
rect 9945 8611 9971 8637
rect 9997 8611 10023 8637
rect 10049 8611 20328 8637
rect 672 8594 20328 8611
rect 7015 8553 7041 8559
rect 7015 8521 7041 8527
rect 7351 8553 7377 8559
rect 7351 8521 7377 8527
rect 7743 8553 7769 8559
rect 7743 8521 7769 8527
rect 7855 8553 7881 8559
rect 7855 8521 7881 8527
rect 9647 8553 9673 8559
rect 9647 8521 9673 8527
rect 9759 8553 9785 8559
rect 9759 8521 9785 8527
rect 11215 8553 11241 8559
rect 11215 8521 11241 8527
rect 13119 8553 13145 8559
rect 13119 8521 13145 8527
rect 7127 8497 7153 8503
rect 7127 8465 7153 8471
rect 7463 8497 7489 8503
rect 7463 8465 7489 8471
rect 8247 8497 8273 8503
rect 8247 8465 8273 8471
rect 8303 8497 8329 8503
rect 14737 8471 14743 8497
rect 14769 8471 14775 8497
rect 8303 8465 8329 8471
rect 6847 8441 6873 8447
rect 2137 8415 2143 8441
rect 2169 8415 2175 8441
rect 6847 8409 6873 8415
rect 6903 8441 6929 8447
rect 6903 8409 6929 8415
rect 6959 8441 6985 8447
rect 6959 8409 6985 8415
rect 7295 8441 7321 8447
rect 7295 8409 7321 8415
rect 7687 8441 7713 8447
rect 8135 8441 8161 8447
rect 7961 8415 7967 8441
rect 7993 8415 7999 8441
rect 7687 8409 7713 8415
rect 8135 8409 8161 8415
rect 9983 8441 10009 8447
rect 9983 8409 10009 8415
rect 11271 8441 11297 8447
rect 11271 8409 11297 8415
rect 13511 8441 13537 8447
rect 15073 8415 15079 8441
rect 15105 8415 15111 8441
rect 13511 8409 13537 8415
rect 7799 8385 7825 8391
rect 7799 8353 7825 8359
rect 9703 8385 9729 8391
rect 13673 8359 13679 8385
rect 13705 8359 13711 8385
rect 9703 8353 9729 8359
rect 967 8329 993 8335
rect 967 8297 993 8303
rect 11215 8329 11241 8335
rect 11215 8297 11241 8303
rect 672 8245 20328 8262
rect 672 8219 2239 8245
rect 2265 8219 2291 8245
rect 2317 8219 2343 8245
rect 2369 8219 17599 8245
rect 17625 8219 17651 8245
rect 17677 8219 17703 8245
rect 17729 8219 20328 8245
rect 672 8202 20328 8219
rect 11999 8161 12025 8167
rect 11999 8129 12025 8135
rect 8415 8105 8441 8111
rect 7121 8079 7127 8105
rect 7153 8079 7159 8105
rect 8185 8079 8191 8105
rect 8217 8079 8223 8105
rect 8415 8073 8441 8079
rect 10711 8105 10737 8111
rect 10711 8073 10737 8079
rect 11439 8049 11465 8055
rect 6785 8023 6791 8049
rect 6817 8023 6823 8049
rect 10873 8023 10879 8049
rect 10905 8023 10911 8049
rect 11041 8023 11047 8049
rect 11073 8023 11079 8049
rect 11439 8017 11465 8023
rect 11551 8049 11577 8055
rect 11551 8017 11577 8023
rect 11943 8049 11969 8055
rect 11943 8017 11969 8023
rect 10655 7993 10681 7999
rect 11495 7993 11521 7999
rect 10655 7961 10681 7967
rect 10767 7965 10793 7971
rect 11495 7961 11521 7967
rect 10767 7933 10793 7939
rect 11999 7937 12025 7943
rect 11769 7911 11775 7937
rect 11801 7911 11807 7937
rect 11999 7905 12025 7911
rect 672 7853 20328 7870
rect 672 7827 9919 7853
rect 9945 7827 9971 7853
rect 9997 7827 10023 7853
rect 10049 7827 20328 7853
rect 672 7810 20328 7827
rect 13511 7769 13537 7775
rect 13511 7737 13537 7743
rect 13623 7769 13649 7775
rect 13623 7737 13649 7743
rect 11663 7713 11689 7719
rect 6561 7687 6567 7713
rect 6593 7687 6599 7713
rect 9585 7687 9591 7713
rect 9617 7687 9623 7713
rect 11663 7681 11689 7687
rect 13399 7657 13425 7663
rect 6953 7631 6959 7657
rect 6985 7631 6991 7657
rect 9193 7631 9199 7657
rect 9225 7631 9231 7657
rect 11545 7631 11551 7657
rect 11577 7631 11583 7657
rect 18825 7631 18831 7657
rect 18857 7631 18863 7657
rect 13399 7625 13425 7631
rect 7183 7601 7209 7607
rect 5497 7575 5503 7601
rect 5529 7575 5535 7601
rect 7183 7569 7209 7575
rect 9031 7601 9057 7607
rect 13455 7601 13481 7607
rect 10649 7575 10655 7601
rect 10681 7575 10687 7601
rect 9031 7569 9057 7575
rect 13455 7569 13481 7575
rect 20007 7601 20033 7607
rect 20007 7569 20033 7575
rect 672 7461 20328 7478
rect 672 7435 2239 7461
rect 2265 7435 2291 7461
rect 2317 7435 2343 7461
rect 2369 7435 17599 7461
rect 17625 7435 17651 7461
rect 17677 7435 17703 7461
rect 17729 7435 20328 7461
rect 672 7418 20328 7435
rect 7967 7377 7993 7383
rect 7967 7345 7993 7351
rect 8079 7377 8105 7383
rect 8079 7345 8105 7351
rect 10879 7377 10905 7383
rect 10879 7345 10905 7351
rect 13175 7377 13201 7383
rect 13175 7345 13201 7351
rect 13343 7377 13369 7383
rect 13343 7345 13369 7351
rect 8527 7321 8553 7327
rect 20007 7321 20033 7327
rect 8409 7295 8415 7321
rect 8441 7295 8447 7321
rect 8689 7295 8695 7321
rect 8721 7295 8727 7321
rect 11713 7295 11719 7321
rect 11745 7295 11751 7321
rect 12777 7295 12783 7321
rect 12809 7295 12815 7321
rect 8527 7289 8553 7295
rect 20007 7289 20033 7295
rect 9367 7265 9393 7271
rect 8185 7239 8191 7265
rect 8217 7239 8223 7265
rect 10201 7239 10207 7265
rect 10233 7239 10239 7265
rect 11041 7239 11047 7265
rect 11073 7239 11079 7265
rect 11321 7239 11327 7265
rect 11353 7239 11359 7265
rect 13337 7239 13343 7265
rect 13369 7239 13375 7265
rect 13897 7239 13903 7265
rect 13929 7239 13935 7265
rect 18825 7239 18831 7265
rect 18857 7239 18863 7265
rect 9367 7233 9393 7239
rect 7911 7209 7937 7215
rect 7911 7177 7937 7183
rect 8751 7209 8777 7215
rect 8751 7177 8777 7183
rect 8863 7209 8889 7215
rect 8863 7177 8889 7183
rect 9423 7209 9449 7215
rect 9423 7177 9449 7183
rect 9591 7209 9617 7215
rect 9591 7177 9617 7183
rect 10375 7209 10401 7215
rect 10375 7177 10401 7183
rect 10935 7209 10961 7215
rect 10935 7177 10961 7183
rect 8415 7153 8441 7159
rect 8415 7121 8441 7127
rect 9479 7153 9505 7159
rect 9479 7121 9505 7127
rect 10319 7153 10345 7159
rect 10319 7121 10345 7127
rect 13007 7153 13033 7159
rect 14009 7127 14015 7153
rect 14041 7127 14047 7153
rect 13007 7121 13033 7127
rect 672 7069 20328 7086
rect 672 7043 9919 7069
rect 9945 7043 9971 7069
rect 9997 7043 10023 7069
rect 10049 7043 20328 7069
rect 672 7026 20328 7043
rect 7345 6903 7351 6929
rect 7377 6903 7383 6929
rect 10537 6903 10543 6929
rect 10569 6903 10575 6929
rect 13169 6903 13175 6929
rect 13201 6903 13207 6929
rect 11831 6873 11857 6879
rect 14463 6873 14489 6879
rect 7009 6847 7015 6873
rect 7041 6847 7047 6873
rect 10201 6847 10207 6873
rect 10233 6847 10239 6873
rect 12777 6847 12783 6873
rect 12809 6847 12815 6873
rect 11831 6841 11857 6847
rect 14463 6841 14489 6847
rect 8751 6817 8777 6823
rect 8409 6791 8415 6817
rect 8441 6791 8447 6817
rect 11601 6791 11607 6817
rect 11633 6791 11639 6817
rect 14233 6791 14239 6817
rect 14265 6791 14271 6817
rect 8751 6785 8777 6791
rect 672 6677 20328 6694
rect 672 6651 2239 6677
rect 2265 6651 2291 6677
rect 2317 6651 2343 6677
rect 2369 6651 17599 6677
rect 17625 6651 17651 6677
rect 17677 6651 17703 6677
rect 17729 6651 20328 6677
rect 672 6634 20328 6651
rect 9927 6537 9953 6543
rect 8633 6511 8639 6537
rect 8665 6511 8671 6537
rect 9697 6511 9703 6537
rect 9729 6511 9735 6537
rect 9927 6505 9953 6511
rect 8297 6455 8303 6481
rect 8329 6455 8335 6481
rect 672 6285 20328 6302
rect 672 6259 9919 6285
rect 9945 6259 9971 6285
rect 9997 6259 10023 6285
rect 10049 6259 20328 6285
rect 672 6242 20328 6259
rect 672 5893 20328 5910
rect 672 5867 2239 5893
rect 2265 5867 2291 5893
rect 2317 5867 2343 5893
rect 2369 5867 17599 5893
rect 17625 5867 17651 5893
rect 17677 5867 17703 5893
rect 17729 5867 20328 5893
rect 672 5850 20328 5867
rect 672 5501 20328 5518
rect 672 5475 9919 5501
rect 9945 5475 9971 5501
rect 9997 5475 10023 5501
rect 10049 5475 20328 5501
rect 672 5458 20328 5475
rect 672 5109 20328 5126
rect 672 5083 2239 5109
rect 2265 5083 2291 5109
rect 2317 5083 2343 5109
rect 2369 5083 17599 5109
rect 17625 5083 17651 5109
rect 17677 5083 17703 5109
rect 17729 5083 20328 5109
rect 672 5066 20328 5083
rect 672 4717 20328 4734
rect 672 4691 9919 4717
rect 9945 4691 9971 4717
rect 9997 4691 10023 4717
rect 10049 4691 20328 4717
rect 672 4674 20328 4691
rect 672 4325 20328 4342
rect 672 4299 2239 4325
rect 2265 4299 2291 4325
rect 2317 4299 2343 4325
rect 2369 4299 17599 4325
rect 17625 4299 17651 4325
rect 17677 4299 17703 4325
rect 17729 4299 20328 4325
rect 672 4282 20328 4299
rect 672 3933 20328 3950
rect 672 3907 9919 3933
rect 9945 3907 9971 3933
rect 9997 3907 10023 3933
rect 10049 3907 20328 3933
rect 672 3890 20328 3907
rect 672 3541 20328 3558
rect 672 3515 2239 3541
rect 2265 3515 2291 3541
rect 2317 3515 2343 3541
rect 2369 3515 17599 3541
rect 17625 3515 17651 3541
rect 17677 3515 17703 3541
rect 17729 3515 20328 3541
rect 672 3498 20328 3515
rect 672 3149 20328 3166
rect 672 3123 9919 3149
rect 9945 3123 9971 3149
rect 9997 3123 10023 3149
rect 10049 3123 20328 3149
rect 672 3106 20328 3123
rect 672 2757 20328 2774
rect 672 2731 2239 2757
rect 2265 2731 2291 2757
rect 2317 2731 2343 2757
rect 2369 2731 17599 2757
rect 17625 2731 17651 2757
rect 17677 2731 17703 2757
rect 17729 2731 20328 2757
rect 672 2714 20328 2731
rect 8695 2617 8721 2623
rect 8695 2585 8721 2591
rect 8185 2535 8191 2561
rect 8217 2535 8223 2561
rect 672 2365 20328 2382
rect 672 2339 9919 2365
rect 9945 2339 9971 2365
rect 9997 2339 10023 2365
rect 10049 2339 20328 2365
rect 672 2322 20328 2339
rect 8689 2143 8695 2169
rect 8721 2143 8727 2169
rect 10537 2143 10543 2169
rect 10569 2143 10575 2169
rect 9199 2057 9225 2063
rect 9199 2025 9225 2031
rect 11047 2057 11073 2063
rect 11047 2025 11073 2031
rect 672 1973 20328 1990
rect 672 1947 2239 1973
rect 2265 1947 2291 1973
rect 2317 1947 2343 1973
rect 2369 1947 17599 1973
rect 17625 1947 17651 1973
rect 17677 1947 17703 1973
rect 17729 1947 20328 1973
rect 672 1930 20328 1947
rect 12783 1833 12809 1839
rect 12783 1801 12809 1807
rect 8801 1751 8807 1777
rect 8833 1751 8839 1777
rect 11937 1751 11943 1777
rect 11969 1751 11975 1777
rect 12273 1751 12279 1777
rect 12305 1751 12311 1777
rect 9697 1695 9703 1721
rect 9729 1695 9735 1721
rect 11097 1695 11103 1721
rect 11129 1695 11135 1721
rect 15247 1665 15273 1671
rect 15247 1633 15273 1639
rect 672 1581 20328 1598
rect 672 1555 9919 1581
rect 9945 1555 9971 1581
rect 9997 1555 10023 1581
rect 10049 1555 20328 1581
rect 672 1538 20328 1555
<< via1 >>
rect 2239 19195 2265 19221
rect 2291 19195 2317 19221
rect 2343 19195 2369 19221
rect 17599 19195 17625 19221
rect 17651 19195 17677 19221
rect 17703 19195 17729 19221
rect 13119 19111 13145 19137
rect 9087 19055 9113 19081
rect 11103 19055 11129 19081
rect 9871 18999 9897 19025
rect 11775 18999 11801 19025
rect 12839 18999 12865 19025
rect 9919 18803 9945 18829
rect 9971 18803 9997 18829
rect 10023 18803 10049 18829
rect 9199 18719 9225 18745
rect 11383 18719 11409 18745
rect 8807 18607 8833 18633
rect 10935 18607 10961 18633
rect 2239 18411 2265 18437
rect 2291 18411 2317 18437
rect 2343 18411 2369 18437
rect 17599 18411 17625 18437
rect 17651 18411 17677 18437
rect 17703 18411 17729 18437
rect 9919 18019 9945 18045
rect 9971 18019 9997 18045
rect 10023 18019 10049 18045
rect 2239 17627 2265 17653
rect 2291 17627 2317 17653
rect 2343 17627 2369 17653
rect 17599 17627 17625 17653
rect 17651 17627 17677 17653
rect 17703 17627 17729 17653
rect 9919 17235 9945 17261
rect 9971 17235 9997 17261
rect 10023 17235 10049 17261
rect 2239 16843 2265 16869
rect 2291 16843 2317 16869
rect 2343 16843 2369 16869
rect 17599 16843 17625 16869
rect 17651 16843 17677 16869
rect 17703 16843 17729 16869
rect 9919 16451 9945 16477
rect 9971 16451 9997 16477
rect 10023 16451 10049 16477
rect 2239 16059 2265 16085
rect 2291 16059 2317 16085
rect 2343 16059 2369 16085
rect 17599 16059 17625 16085
rect 17651 16059 17677 16085
rect 17703 16059 17729 16085
rect 9919 15667 9945 15693
rect 9971 15667 9997 15693
rect 10023 15667 10049 15693
rect 2239 15275 2265 15301
rect 2291 15275 2317 15301
rect 2343 15275 2369 15301
rect 17599 15275 17625 15301
rect 17651 15275 17677 15301
rect 17703 15275 17729 15301
rect 9919 14883 9945 14909
rect 9971 14883 9997 14909
rect 10023 14883 10049 14909
rect 2239 14491 2265 14517
rect 2291 14491 2317 14517
rect 2343 14491 2369 14517
rect 17599 14491 17625 14517
rect 17651 14491 17677 14517
rect 17703 14491 17729 14517
rect 9919 14099 9945 14125
rect 9971 14099 9997 14125
rect 10023 14099 10049 14125
rect 18831 13903 18857 13929
rect 19951 13847 19977 13873
rect 2239 13707 2265 13733
rect 2291 13707 2317 13733
rect 2343 13707 2369 13733
rect 17599 13707 17625 13733
rect 17651 13707 17677 13733
rect 17703 13707 17729 13733
rect 8583 13567 8609 13593
rect 20007 13567 20033 13593
rect 7183 13511 7209 13537
rect 10655 13511 10681 13537
rect 10991 13511 11017 13537
rect 13455 13511 13481 13537
rect 18943 13511 18969 13537
rect 7519 13455 7545 13481
rect 8695 13455 8721 13481
rect 8807 13455 8833 13481
rect 8863 13455 8889 13481
rect 9087 13455 9113 13481
rect 12559 13455 12585 13481
rect 12615 13455 12641 13481
rect 13567 13455 13593 13481
rect 10711 13399 10737 13425
rect 10767 13399 10793 13425
rect 12727 13399 12753 13425
rect 9919 13315 9945 13341
rect 9971 13315 9997 13341
rect 10023 13315 10049 13341
rect 8079 13231 8105 13257
rect 9311 13231 9337 13257
rect 11383 13231 11409 13257
rect 11495 13231 11521 13257
rect 10207 13175 10233 13201
rect 11551 13175 11577 13201
rect 12279 13175 12305 13201
rect 12335 13175 12361 13201
rect 8023 13119 8049 13145
rect 8191 13119 8217 13145
rect 9479 13119 9505 13145
rect 9871 13119 9897 13145
rect 11831 13119 11857 13145
rect 12167 13119 12193 13145
rect 12615 13119 12641 13145
rect 18831 13119 18857 13145
rect 11271 13063 11297 13089
rect 13007 13063 13033 13089
rect 14127 13063 14153 13089
rect 14463 13063 14489 13089
rect 20007 13007 20033 13033
rect 2239 12923 2265 12949
rect 2291 12923 2317 12949
rect 2343 12923 2369 12949
rect 17599 12923 17625 12949
rect 17651 12923 17677 12949
rect 17703 12923 17729 12949
rect 9255 12783 9281 12809
rect 12951 12783 12977 12809
rect 13175 12783 13201 12809
rect 7799 12727 7825 12753
rect 9535 12727 9561 12753
rect 10431 12727 10457 12753
rect 10599 12727 10625 12753
rect 11551 12727 11577 12753
rect 13455 12727 13481 12753
rect 8191 12671 8217 12697
rect 9479 12671 9505 12697
rect 10263 12671 10289 12697
rect 10319 12671 10345 12697
rect 11887 12671 11913 12697
rect 13567 12671 13593 12697
rect 9367 12615 9393 12641
rect 9759 12615 9785 12641
rect 10823 12615 10849 12641
rect 10879 12615 10905 12641
rect 10935 12615 10961 12641
rect 9919 12531 9945 12557
rect 9971 12531 9997 12557
rect 10023 12531 10049 12557
rect 6007 12447 6033 12473
rect 8415 12447 8441 12473
rect 8751 12447 8777 12473
rect 9423 12447 9449 12473
rect 11607 12447 11633 12473
rect 11663 12447 11689 12473
rect 12783 12447 12809 12473
rect 7967 12391 7993 12417
rect 9199 12391 9225 12417
rect 9983 12391 10009 12417
rect 12615 12391 12641 12417
rect 12671 12391 12697 12417
rect 20119 12391 20145 12417
rect 5895 12335 5921 12361
rect 6175 12335 6201 12361
rect 6567 12335 6593 12361
rect 8079 12335 8105 12361
rect 8247 12335 8273 12361
rect 9143 12335 9169 12361
rect 9647 12335 9673 12361
rect 11719 12335 11745 12361
rect 11943 12335 11969 12361
rect 7631 12279 7657 12305
rect 8023 12279 8049 12305
rect 8807 12279 8833 12305
rect 11047 12279 11073 12305
rect 8919 12223 8945 12249
rect 2239 12139 2265 12165
rect 2291 12139 2317 12165
rect 2343 12139 2369 12165
rect 17599 12139 17625 12165
rect 17651 12139 17677 12165
rect 17703 12139 17729 12165
rect 10655 12055 10681 12081
rect 7743 11999 7769 12025
rect 7911 11999 7937 12025
rect 10823 11943 10849 11969
rect 10935 11943 10961 11969
rect 9919 11747 9945 11773
rect 9971 11747 9997 11773
rect 10023 11747 10049 11773
rect 9087 11663 9113 11689
rect 6231 11607 6257 11633
rect 8079 11607 8105 11633
rect 8247 11607 8273 11633
rect 8695 11607 8721 11633
rect 10095 11607 10121 11633
rect 12895 11607 12921 11633
rect 5895 11551 5921 11577
rect 7911 11551 7937 11577
rect 8359 11551 8385 11577
rect 8807 11551 8833 11577
rect 8975 11551 9001 11577
rect 10207 11551 10233 11577
rect 10655 11551 10681 11577
rect 12335 11551 12361 11577
rect 12671 11551 12697 11577
rect 13063 11551 13089 11577
rect 13231 11551 13257 11577
rect 13735 11551 13761 11577
rect 13847 11551 13873 11577
rect 13959 11551 13985 11577
rect 14015 11551 14041 11577
rect 7295 11495 7321 11521
rect 7519 11495 7545 11521
rect 10487 11495 10513 11521
rect 10879 11495 10905 11521
rect 11943 11495 11969 11521
rect 13343 11495 13369 11521
rect 8975 11439 9001 11465
rect 13063 11439 13089 11465
rect 13399 11439 13425 11465
rect 2239 11355 2265 11381
rect 2291 11355 2317 11381
rect 2343 11355 2369 11381
rect 17599 11355 17625 11381
rect 17651 11355 17677 11381
rect 17703 11355 17729 11381
rect 10319 11271 10345 11297
rect 11831 11271 11857 11297
rect 10767 11215 10793 11241
rect 11551 11215 11577 11241
rect 13231 11215 13257 11241
rect 14295 11215 14321 11241
rect 14631 11215 14657 11241
rect 20007 11215 20033 11241
rect 7463 11159 7489 11185
rect 7743 11159 7769 11185
rect 7855 11159 7881 11185
rect 8079 11159 8105 11185
rect 8135 11159 8161 11185
rect 8415 11159 8441 11185
rect 8751 11159 8777 11185
rect 9199 11159 9225 11185
rect 9423 11159 9449 11185
rect 10095 11159 10121 11185
rect 10319 11159 10345 11185
rect 10655 11159 10681 11185
rect 11103 11159 11129 11185
rect 11607 11159 11633 11185
rect 12839 11159 12865 11185
rect 18831 11159 18857 11185
rect 9143 11103 9169 11129
rect 11159 11103 11185 11129
rect 11775 11103 11801 11129
rect 8023 11047 8049 11073
rect 8527 11047 8553 11073
rect 8863 11047 8889 11073
rect 9535 11047 9561 11073
rect 10935 11047 10961 11073
rect 11383 11047 11409 11073
rect 11495 11047 11521 11073
rect 11831 11047 11857 11073
rect 9919 10963 9945 10989
rect 9971 10963 9997 10989
rect 10023 10963 10049 10989
rect 7407 10879 7433 10905
rect 8079 10879 8105 10905
rect 10935 10879 10961 10905
rect 11719 10879 11745 10905
rect 14631 10879 14657 10905
rect 8695 10823 8721 10849
rect 9311 10823 9337 10849
rect 9815 10823 9841 10849
rect 13343 10823 13369 10849
rect 5783 10767 5809 10793
rect 8023 10767 8049 10793
rect 8247 10767 8273 10793
rect 8863 10767 8889 10793
rect 9255 10767 9281 10793
rect 10599 10767 10625 10793
rect 10823 10767 10849 10793
rect 11159 10767 11185 10793
rect 11383 10767 11409 10793
rect 11439 10767 11465 10793
rect 11495 10767 11521 10793
rect 12951 10767 12977 10793
rect 18831 10767 18857 10793
rect 6119 10711 6145 10737
rect 7183 10711 7209 10737
rect 10655 10711 10681 10737
rect 10879 10711 10905 10737
rect 14407 10711 14433 10737
rect 20007 10711 20033 10737
rect 2239 10571 2265 10597
rect 2291 10571 2317 10597
rect 2343 10571 2369 10597
rect 17599 10571 17625 10597
rect 17651 10571 17677 10597
rect 17703 10571 17729 10597
rect 9143 10487 9169 10513
rect 9311 10487 9337 10513
rect 10767 10487 10793 10513
rect 967 10431 993 10457
rect 8023 10431 8049 10457
rect 9031 10431 9057 10457
rect 9759 10431 9785 10457
rect 12951 10431 12977 10457
rect 2143 10375 2169 10401
rect 8135 10375 8161 10401
rect 9479 10375 9505 10401
rect 10095 10375 10121 10401
rect 10991 10375 11017 10401
rect 11775 10375 11801 10401
rect 7799 10319 7825 10345
rect 10823 10319 10849 10345
rect 11327 10319 11353 10345
rect 10263 10263 10289 10289
rect 10767 10263 10793 10289
rect 11159 10263 11185 10289
rect 11383 10263 11409 10289
rect 11495 10263 11521 10289
rect 9919 10179 9945 10205
rect 9971 10179 9997 10205
rect 10023 10179 10049 10205
rect 8751 10095 8777 10121
rect 9087 10095 9113 10121
rect 7351 10039 7377 10065
rect 7519 10039 7545 10065
rect 7799 10039 7825 10065
rect 7911 10039 7937 10065
rect 8359 10039 8385 10065
rect 8863 10039 8889 10065
rect 11719 10039 11745 10065
rect 13567 10039 13593 10065
rect 13791 10039 13817 10065
rect 13903 10039 13929 10065
rect 14015 10039 14041 10065
rect 6791 9983 6817 10009
rect 7239 9983 7265 10009
rect 7967 9983 7993 10009
rect 9031 9983 9057 10009
rect 9199 9983 9225 10009
rect 9703 9983 9729 10009
rect 13399 9983 13425 10009
rect 13679 9983 13705 10009
rect 5335 9927 5361 9953
rect 6399 9927 6425 9953
rect 7015 9927 7041 9953
rect 7183 9927 7209 9953
rect 9535 9927 9561 9953
rect 7631 9871 7657 9897
rect 7687 9871 7713 9897
rect 8415 9871 8441 9897
rect 8695 9871 8721 9897
rect 2239 9787 2265 9813
rect 2291 9787 2317 9813
rect 2343 9787 2369 9813
rect 17599 9787 17625 9813
rect 17651 9787 17677 9813
rect 17703 9787 17729 9813
rect 6175 9703 6201 9729
rect 6791 9703 6817 9729
rect 13735 9703 13761 9729
rect 6231 9647 6257 9673
rect 13119 9647 13145 9673
rect 13959 9647 13985 9673
rect 20007 9647 20033 9673
rect 7575 9591 7601 9617
rect 10039 9591 10065 9617
rect 11327 9591 11353 9617
rect 11607 9591 11633 9617
rect 12615 9591 12641 9617
rect 14127 9591 14153 9617
rect 18831 9591 18857 9617
rect 6847 9535 6873 9561
rect 8471 9535 8497 9561
rect 10823 9535 10849 9561
rect 11943 9535 11969 9561
rect 12783 9535 12809 9561
rect 13007 9535 13033 9561
rect 13903 9535 13929 9561
rect 14071 9535 14097 9561
rect 6791 9479 6817 9505
rect 7407 9479 7433 9505
rect 10655 9479 10681 9505
rect 11159 9479 11185 9505
rect 11495 9479 11521 9505
rect 11775 9479 11801 9505
rect 11887 9479 11913 9505
rect 13063 9479 13089 9505
rect 13623 9479 13649 9505
rect 13679 9479 13705 9505
rect 9919 9395 9945 9421
rect 9971 9395 9997 9421
rect 10023 9395 10049 9421
rect 7855 9311 7881 9337
rect 7967 9311 7993 9337
rect 8359 9311 8385 9337
rect 9199 9311 9225 9337
rect 9591 9311 9617 9337
rect 9983 9311 10009 9337
rect 8079 9255 8105 9281
rect 8303 9255 8329 9281
rect 9255 9255 9281 9281
rect 9759 9255 9785 9281
rect 9927 9255 9953 9281
rect 10263 9255 10289 9281
rect 10319 9255 10345 9281
rect 11999 9255 12025 9281
rect 13735 9255 13761 9281
rect 2143 9199 2169 9225
rect 6231 9199 6257 9225
rect 6623 9199 6649 9225
rect 6791 9199 6817 9225
rect 6847 9199 6873 9225
rect 6903 9199 6929 9225
rect 7071 9199 7097 9225
rect 7799 9199 7825 9225
rect 8639 9199 8665 9225
rect 8807 9199 8833 9225
rect 8975 9199 9001 9225
rect 10431 9199 10457 9225
rect 10655 9199 10681 9225
rect 10767 9199 10793 9225
rect 11215 9199 11241 9225
rect 11271 9199 11297 9225
rect 11495 9199 11521 9225
rect 11607 9199 11633 9225
rect 11775 9199 11801 9225
rect 12111 9199 12137 9225
rect 13343 9199 13369 9225
rect 15023 9199 15049 9225
rect 18831 9199 18857 9225
rect 5167 9143 5193 9169
rect 7295 9143 7321 9169
rect 8751 9143 8777 9169
rect 11103 9143 11129 9169
rect 11887 9143 11913 9169
rect 14799 9143 14825 9169
rect 967 9087 993 9113
rect 8359 9087 8385 9113
rect 9199 9087 9225 9113
rect 9983 9087 10009 9113
rect 10935 9087 10961 9113
rect 20007 9087 20033 9113
rect 2239 9003 2265 9029
rect 2291 9003 2317 9029
rect 2343 9003 2369 9029
rect 17599 9003 17625 9029
rect 17651 9003 17677 9029
rect 17703 9003 17729 9029
rect 6791 8919 6817 8945
rect 9143 8919 9169 8945
rect 13287 8919 13313 8945
rect 14071 8919 14097 8945
rect 9927 8863 9953 8889
rect 11943 8863 11969 8889
rect 13007 8863 13033 8889
rect 13175 8863 13201 8889
rect 20007 8863 20033 8889
rect 8583 8807 8609 8833
rect 9535 8807 9561 8833
rect 9983 8807 10009 8833
rect 11607 8807 11633 8833
rect 13791 8807 13817 8833
rect 14239 8807 14265 8833
rect 14575 8807 14601 8833
rect 14687 8807 14713 8833
rect 15135 8807 15161 8833
rect 18831 8807 18857 8833
rect 6791 8751 6817 8777
rect 6847 8751 6873 8777
rect 8303 8751 8329 8777
rect 9031 8751 9057 8777
rect 9367 8751 9393 8777
rect 9759 8751 9785 8777
rect 13679 8751 13705 8777
rect 14855 8751 14881 8777
rect 8247 8695 8273 8721
rect 8415 8695 8441 8721
rect 9087 8695 9113 8721
rect 9871 8695 9897 8721
rect 13455 8695 13481 8721
rect 15023 8695 15049 8721
rect 9919 8611 9945 8637
rect 9971 8611 9997 8637
rect 10023 8611 10049 8637
rect 7015 8527 7041 8553
rect 7351 8527 7377 8553
rect 7743 8527 7769 8553
rect 7855 8527 7881 8553
rect 9647 8527 9673 8553
rect 9759 8527 9785 8553
rect 11215 8527 11241 8553
rect 13119 8527 13145 8553
rect 7127 8471 7153 8497
rect 7463 8471 7489 8497
rect 8247 8471 8273 8497
rect 8303 8471 8329 8497
rect 14743 8471 14769 8497
rect 2143 8415 2169 8441
rect 6847 8415 6873 8441
rect 6903 8415 6929 8441
rect 6959 8415 6985 8441
rect 7295 8415 7321 8441
rect 7687 8415 7713 8441
rect 7967 8415 7993 8441
rect 8135 8415 8161 8441
rect 9983 8415 10009 8441
rect 11271 8415 11297 8441
rect 13511 8415 13537 8441
rect 15079 8415 15105 8441
rect 7799 8359 7825 8385
rect 9703 8359 9729 8385
rect 13679 8359 13705 8385
rect 967 8303 993 8329
rect 11215 8303 11241 8329
rect 2239 8219 2265 8245
rect 2291 8219 2317 8245
rect 2343 8219 2369 8245
rect 17599 8219 17625 8245
rect 17651 8219 17677 8245
rect 17703 8219 17729 8245
rect 11999 8135 12025 8161
rect 7127 8079 7153 8105
rect 8191 8079 8217 8105
rect 8415 8079 8441 8105
rect 10711 8079 10737 8105
rect 6791 8023 6817 8049
rect 10879 8023 10905 8049
rect 11047 8023 11073 8049
rect 11439 8023 11465 8049
rect 11551 8023 11577 8049
rect 11943 8023 11969 8049
rect 10655 7967 10681 7993
rect 10767 7939 10793 7965
rect 11495 7967 11521 7993
rect 11775 7911 11801 7937
rect 11999 7911 12025 7937
rect 9919 7827 9945 7853
rect 9971 7827 9997 7853
rect 10023 7827 10049 7853
rect 13511 7743 13537 7769
rect 13623 7743 13649 7769
rect 6567 7687 6593 7713
rect 9591 7687 9617 7713
rect 11663 7687 11689 7713
rect 6959 7631 6985 7657
rect 9199 7631 9225 7657
rect 11551 7631 11577 7657
rect 13399 7631 13425 7657
rect 18831 7631 18857 7657
rect 5503 7575 5529 7601
rect 7183 7575 7209 7601
rect 9031 7575 9057 7601
rect 10655 7575 10681 7601
rect 13455 7575 13481 7601
rect 20007 7575 20033 7601
rect 2239 7435 2265 7461
rect 2291 7435 2317 7461
rect 2343 7435 2369 7461
rect 17599 7435 17625 7461
rect 17651 7435 17677 7461
rect 17703 7435 17729 7461
rect 7967 7351 7993 7377
rect 8079 7351 8105 7377
rect 10879 7351 10905 7377
rect 13175 7351 13201 7377
rect 13343 7351 13369 7377
rect 8415 7295 8441 7321
rect 8527 7295 8553 7321
rect 8695 7295 8721 7321
rect 11719 7295 11745 7321
rect 12783 7295 12809 7321
rect 20007 7295 20033 7321
rect 8191 7239 8217 7265
rect 9367 7239 9393 7265
rect 10207 7239 10233 7265
rect 11047 7239 11073 7265
rect 11327 7239 11353 7265
rect 13343 7239 13369 7265
rect 13903 7239 13929 7265
rect 18831 7239 18857 7265
rect 7911 7183 7937 7209
rect 8751 7183 8777 7209
rect 8863 7183 8889 7209
rect 9423 7183 9449 7209
rect 9591 7183 9617 7209
rect 10375 7183 10401 7209
rect 10935 7183 10961 7209
rect 8415 7127 8441 7153
rect 9479 7127 9505 7153
rect 10319 7127 10345 7153
rect 13007 7127 13033 7153
rect 14015 7127 14041 7153
rect 9919 7043 9945 7069
rect 9971 7043 9997 7069
rect 10023 7043 10049 7069
rect 7351 6903 7377 6929
rect 10543 6903 10569 6929
rect 13175 6903 13201 6929
rect 7015 6847 7041 6873
rect 10207 6847 10233 6873
rect 11831 6847 11857 6873
rect 12783 6847 12809 6873
rect 14463 6847 14489 6873
rect 8415 6791 8441 6817
rect 8751 6791 8777 6817
rect 11607 6791 11633 6817
rect 14239 6791 14265 6817
rect 2239 6651 2265 6677
rect 2291 6651 2317 6677
rect 2343 6651 2369 6677
rect 17599 6651 17625 6677
rect 17651 6651 17677 6677
rect 17703 6651 17729 6677
rect 8639 6511 8665 6537
rect 9703 6511 9729 6537
rect 9927 6511 9953 6537
rect 8303 6455 8329 6481
rect 9919 6259 9945 6285
rect 9971 6259 9997 6285
rect 10023 6259 10049 6285
rect 2239 5867 2265 5893
rect 2291 5867 2317 5893
rect 2343 5867 2369 5893
rect 17599 5867 17625 5893
rect 17651 5867 17677 5893
rect 17703 5867 17729 5893
rect 9919 5475 9945 5501
rect 9971 5475 9997 5501
rect 10023 5475 10049 5501
rect 2239 5083 2265 5109
rect 2291 5083 2317 5109
rect 2343 5083 2369 5109
rect 17599 5083 17625 5109
rect 17651 5083 17677 5109
rect 17703 5083 17729 5109
rect 9919 4691 9945 4717
rect 9971 4691 9997 4717
rect 10023 4691 10049 4717
rect 2239 4299 2265 4325
rect 2291 4299 2317 4325
rect 2343 4299 2369 4325
rect 17599 4299 17625 4325
rect 17651 4299 17677 4325
rect 17703 4299 17729 4325
rect 9919 3907 9945 3933
rect 9971 3907 9997 3933
rect 10023 3907 10049 3933
rect 2239 3515 2265 3541
rect 2291 3515 2317 3541
rect 2343 3515 2369 3541
rect 17599 3515 17625 3541
rect 17651 3515 17677 3541
rect 17703 3515 17729 3541
rect 9919 3123 9945 3149
rect 9971 3123 9997 3149
rect 10023 3123 10049 3149
rect 2239 2731 2265 2757
rect 2291 2731 2317 2757
rect 2343 2731 2369 2757
rect 17599 2731 17625 2757
rect 17651 2731 17677 2757
rect 17703 2731 17729 2757
rect 8695 2591 8721 2617
rect 8191 2535 8217 2561
rect 9919 2339 9945 2365
rect 9971 2339 9997 2365
rect 10023 2339 10049 2365
rect 8695 2143 8721 2169
rect 10543 2143 10569 2169
rect 9199 2031 9225 2057
rect 11047 2031 11073 2057
rect 2239 1947 2265 1973
rect 2291 1947 2317 1973
rect 2343 1947 2369 1973
rect 17599 1947 17625 1973
rect 17651 1947 17677 1973
rect 17703 1947 17729 1973
rect 12783 1807 12809 1833
rect 8807 1751 8833 1777
rect 11943 1751 11969 1777
rect 12279 1751 12305 1777
rect 9703 1695 9729 1721
rect 11103 1695 11129 1721
rect 15247 1639 15273 1665
rect 9919 1555 9945 1581
rect 9971 1555 9997 1581
rect 10023 1555 10049 1581
<< metal2 >>
rect 8400 20600 8456 21000
rect 9072 20600 9128 21000
rect 10752 20600 10808 21000
rect 11088 20600 11144 21000
rect 12768 20600 12824 21000
rect 12950 20622 13146 20650
rect 2238 19222 2370 19227
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2238 19189 2370 19194
rect 8414 18746 8442 20600
rect 9086 19081 9114 20600
rect 9086 19055 9087 19081
rect 9113 19055 9114 19081
rect 9086 19049 9114 19055
rect 9870 19026 9898 19031
rect 9422 19025 9898 19026
rect 9422 18999 9871 19025
rect 9897 18999 9898 19025
rect 9422 18998 9898 18999
rect 8414 18713 8442 18718
rect 9198 18746 9226 18751
rect 9198 18699 9226 18718
rect 8806 18633 8834 18639
rect 8806 18607 8807 18633
rect 8833 18607 8834 18633
rect 2238 18438 2370 18443
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2238 18405 2370 18410
rect 2238 17654 2370 17659
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2238 17621 2370 17626
rect 2238 16870 2370 16875
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2238 16837 2370 16842
rect 2238 16086 2370 16091
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2238 16053 2370 16058
rect 2238 15302 2370 15307
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2238 15269 2370 15274
rect 2238 14518 2370 14523
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2238 14485 2370 14490
rect 2238 13734 2370 13739
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2238 13701 2370 13706
rect 8582 13594 8610 13599
rect 8806 13594 8834 18607
rect 8582 13593 8834 13594
rect 8582 13567 8583 13593
rect 8609 13567 8834 13593
rect 8582 13566 8834 13567
rect 8582 13561 8610 13566
rect 7182 13537 7210 13543
rect 7182 13511 7183 13537
rect 7209 13511 7210 13537
rect 2086 13482 2114 13487
rect 966 10457 994 10463
rect 966 10431 967 10457
rect 993 10431 994 10457
rect 966 10122 994 10431
rect 966 10089 994 10094
rect 2086 9954 2114 13454
rect 2238 12950 2370 12955
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2238 12917 2370 12922
rect 7182 12754 7210 13511
rect 7518 13481 7546 13487
rect 7518 13455 7519 13481
rect 7545 13455 7546 13481
rect 7518 13146 7546 13455
rect 8078 13482 8106 13487
rect 8078 13257 8106 13454
rect 8694 13482 8722 13487
rect 8694 13435 8722 13454
rect 8806 13481 8834 13566
rect 8806 13455 8807 13481
rect 8833 13455 8834 13481
rect 8806 13449 8834 13455
rect 8862 13481 8890 13487
rect 8862 13455 8863 13481
rect 8889 13455 8890 13481
rect 8078 13231 8079 13257
rect 8105 13231 8106 13257
rect 8078 13225 8106 13231
rect 8862 13258 8890 13455
rect 8862 13225 8890 13230
rect 9086 13481 9114 13487
rect 9086 13455 9087 13481
rect 9113 13455 9114 13481
rect 7518 13113 7546 13118
rect 8022 13145 8050 13151
rect 8022 13119 8023 13145
rect 8049 13119 8050 13145
rect 7182 12721 7210 12726
rect 7518 12754 7546 12759
rect 6006 12474 6034 12479
rect 6006 12473 6258 12474
rect 6006 12447 6007 12473
rect 6033 12447 6258 12473
rect 6006 12446 6258 12447
rect 6006 12441 6034 12446
rect 5894 12361 5922 12367
rect 5894 12335 5895 12361
rect 5921 12335 5922 12361
rect 2238 12166 2370 12171
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2238 12133 2370 12138
rect 5894 12082 5922 12335
rect 5894 12049 5922 12054
rect 6174 12361 6202 12367
rect 6174 12335 6175 12361
rect 6201 12335 6202 12361
rect 5894 11578 5922 11583
rect 6174 11578 6202 12335
rect 6230 11633 6258 12446
rect 6566 12362 6594 12367
rect 6566 12315 6594 12334
rect 6230 11607 6231 11633
rect 6257 11607 6258 11633
rect 6230 11601 6258 11607
rect 5894 11577 6202 11578
rect 5894 11551 5895 11577
rect 5921 11551 6202 11577
rect 5894 11550 6202 11551
rect 2238 11382 2370 11387
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2238 11349 2370 11354
rect 5894 10962 5922 11550
rect 7294 11521 7322 11527
rect 7294 11495 7295 11521
rect 7321 11495 7322 11521
rect 7294 11186 7322 11495
rect 7518 11521 7546 12726
rect 7798 12754 7826 12759
rect 7798 12707 7826 12726
rect 7966 12417 7994 12423
rect 7966 12391 7967 12417
rect 7993 12391 7994 12417
rect 7966 12362 7994 12391
rect 7910 12334 7966 12362
rect 7630 12306 7658 12311
rect 7630 12305 7770 12306
rect 7630 12279 7631 12305
rect 7657 12279 7770 12305
rect 7630 12278 7770 12279
rect 7630 12273 7658 12278
rect 7518 11495 7519 11521
rect 7545 11495 7546 11521
rect 7462 11186 7490 11191
rect 7294 11158 7462 11186
rect 7462 11139 7490 11158
rect 5838 10934 5922 10962
rect 7182 11130 7210 11135
rect 5838 10906 5866 10934
rect 5782 10794 5810 10799
rect 5838 10794 5866 10878
rect 5782 10793 5866 10794
rect 5782 10767 5783 10793
rect 5809 10767 5866 10793
rect 5782 10766 5866 10767
rect 5782 10761 5810 10766
rect 6118 10737 6146 10743
rect 6118 10711 6119 10737
rect 6145 10711 6146 10737
rect 2238 10598 2370 10603
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2238 10565 2370 10570
rect 2142 10402 2170 10407
rect 2142 10355 2170 10374
rect 5334 10402 5362 10407
rect 2086 9921 2114 9926
rect 5334 9953 5362 10374
rect 5334 9927 5335 9953
rect 5361 9927 5362 9953
rect 5334 9842 5362 9927
rect 2238 9814 2370 9819
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 5334 9809 5362 9814
rect 2238 9781 2370 9786
rect 6118 9786 6146 10711
rect 7182 10737 7210 11102
rect 7406 10906 7434 10911
rect 7518 10906 7546 11495
rect 7742 12025 7770 12278
rect 7742 11999 7743 12025
rect 7769 11999 7770 12025
rect 7742 11522 7770 11999
rect 7910 12025 7938 12334
rect 7966 12329 7994 12334
rect 8022 12305 8050 13119
rect 8190 13146 8218 13151
rect 8190 13099 8218 13118
rect 8414 12754 8442 12759
rect 8190 12697 8218 12703
rect 8190 12671 8191 12697
rect 8217 12671 8218 12697
rect 8190 12530 8218 12671
rect 8190 12497 8218 12502
rect 8414 12474 8442 12726
rect 8414 12427 8442 12446
rect 8750 12530 8778 12535
rect 8750 12473 8778 12502
rect 8750 12447 8751 12473
rect 8777 12447 8778 12473
rect 8750 12441 8778 12447
rect 9086 12474 9114 13455
rect 9422 13454 9450 18998
rect 9870 18993 9898 18998
rect 9918 18830 10050 18835
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 9918 18797 10050 18802
rect 10766 18746 10794 20600
rect 11102 19081 11130 20600
rect 12782 20538 12810 20600
rect 12950 20594 12978 20622
rect 12894 20566 12978 20594
rect 12894 20538 12922 20566
rect 12782 20510 12922 20538
rect 13118 19137 13146 20622
rect 17598 19222 17730 19227
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17598 19189 17730 19194
rect 13118 19111 13119 19137
rect 13145 19111 13146 19137
rect 13118 19105 13146 19111
rect 11102 19055 11103 19081
rect 11129 19055 11130 19081
rect 11102 19049 11130 19055
rect 11774 19025 11802 19031
rect 11774 18999 11775 19025
rect 11801 18999 11802 19025
rect 10766 18713 10794 18718
rect 11382 18746 11410 18751
rect 11382 18699 11410 18718
rect 10934 18633 10962 18639
rect 10934 18607 10935 18633
rect 10961 18607 10962 18633
rect 9918 18046 10050 18051
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 9918 18013 10050 18018
rect 9918 17262 10050 17267
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 9918 17229 10050 17234
rect 9918 16478 10050 16483
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 9918 16445 10050 16450
rect 9918 15694 10050 15699
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 9918 15661 10050 15666
rect 9918 14910 10050 14915
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 9918 14877 10050 14882
rect 9918 14126 10050 14131
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 9918 14093 10050 14098
rect 10654 13538 10682 13543
rect 10654 13537 10850 13538
rect 10654 13511 10655 13537
rect 10681 13511 10850 13537
rect 10654 13510 10850 13511
rect 10654 13505 10682 13510
rect 9254 13426 9450 13454
rect 9254 12810 9282 13426
rect 10710 13425 10738 13431
rect 10710 13399 10711 13425
rect 10737 13399 10738 13425
rect 9918 13342 10050 13347
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 9918 13309 10050 13314
rect 9310 13258 9338 13263
rect 9310 13211 9338 13230
rect 10206 13202 10234 13207
rect 10710 13202 10738 13399
rect 10206 13201 10738 13202
rect 10206 13175 10207 13201
rect 10233 13175 10738 13201
rect 10206 13174 10738 13175
rect 10766 13425 10794 13431
rect 10766 13399 10767 13425
rect 10793 13399 10794 13425
rect 10206 13169 10234 13174
rect 9478 13146 9506 13151
rect 9870 13146 9898 13151
rect 9478 13145 9562 13146
rect 9478 13119 9479 13145
rect 9505 13119 9562 13145
rect 9478 13118 9562 13119
rect 9478 13113 9506 13118
rect 9254 12809 9506 12810
rect 9254 12783 9255 12809
rect 9281 12783 9506 12809
rect 9254 12782 9506 12783
rect 9254 12777 9282 12782
rect 9478 12697 9506 12782
rect 9534 12754 9562 13118
rect 9870 13099 9898 13118
rect 9534 12707 9562 12726
rect 10262 12754 10290 12759
rect 9478 12671 9479 12697
rect 9505 12671 9506 12697
rect 9478 12665 9506 12671
rect 10262 12697 10290 12726
rect 10430 12754 10458 12759
rect 10598 12754 10626 12759
rect 10430 12753 10626 12754
rect 10430 12727 10431 12753
rect 10457 12727 10599 12753
rect 10625 12727 10626 12753
rect 10430 12726 10626 12727
rect 10430 12721 10458 12726
rect 10598 12721 10626 12726
rect 10262 12671 10263 12697
rect 10289 12671 10290 12697
rect 9366 12642 9394 12647
rect 9086 12441 9114 12446
rect 9198 12641 9394 12642
rect 9198 12615 9367 12641
rect 9393 12615 9394 12641
rect 9198 12614 9394 12615
rect 9198 12417 9226 12614
rect 9366 12609 9394 12614
rect 9758 12641 9786 12647
rect 9758 12615 9759 12641
rect 9785 12615 9786 12641
rect 9422 12474 9450 12479
rect 9422 12427 9450 12446
rect 9646 12474 9674 12479
rect 9758 12474 9786 12615
rect 10094 12642 10122 12647
rect 9918 12558 10050 12563
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 9918 12525 10050 12530
rect 10094 12474 10122 12614
rect 9674 12446 9786 12474
rect 9982 12446 10122 12474
rect 9198 12391 9199 12417
rect 9225 12391 9226 12417
rect 9198 12385 9226 12391
rect 8022 12279 8023 12305
rect 8049 12279 8050 12305
rect 8022 12273 8050 12279
rect 8078 12361 8106 12367
rect 8078 12335 8079 12361
rect 8105 12335 8106 12361
rect 8078 12250 8106 12335
rect 8078 12217 8106 12222
rect 8246 12361 8274 12367
rect 8246 12335 8247 12361
rect 8273 12335 8274 12361
rect 7910 11999 7911 12025
rect 7937 11999 7938 12025
rect 7910 11993 7938 11999
rect 7966 11746 7994 11751
rect 7742 11489 7770 11494
rect 7910 11577 7938 11583
rect 7910 11551 7911 11577
rect 7937 11551 7938 11577
rect 7434 10878 7546 10906
rect 7742 11185 7770 11191
rect 7742 11159 7743 11185
rect 7769 11159 7770 11185
rect 7406 10859 7434 10878
rect 7182 10711 7183 10737
rect 7209 10711 7210 10737
rect 7182 10705 7210 10711
rect 7350 10850 7378 10855
rect 7350 10065 7378 10822
rect 7462 10094 7490 10878
rect 7742 10850 7770 11159
rect 7854 11186 7882 11191
rect 7910 11186 7938 11551
rect 7882 11158 7938 11186
rect 7854 11139 7882 11158
rect 7966 10906 7994 11718
rect 8246 11746 8274 12335
rect 9142 12362 9170 12367
rect 8806 12306 8834 12311
rect 8806 12259 8834 12278
rect 8918 12250 8946 12255
rect 8246 11713 8274 11718
rect 8694 11746 8722 11751
rect 8078 11634 8106 11639
rect 8078 11587 8106 11606
rect 8246 11633 8274 11639
rect 8246 11607 8247 11633
rect 8273 11607 8274 11633
rect 8078 11522 8106 11527
rect 8022 11242 8050 11247
rect 8022 11073 8050 11214
rect 8078 11186 8106 11494
rect 8078 11139 8106 11158
rect 8134 11185 8162 11191
rect 8134 11159 8135 11185
rect 8161 11159 8162 11185
rect 8134 11130 8162 11159
rect 8134 11097 8162 11102
rect 8022 11047 8023 11073
rect 8049 11047 8050 11073
rect 8022 11041 8050 11047
rect 8246 10962 8274 11607
rect 8694 11633 8722 11718
rect 8694 11607 8695 11633
rect 8721 11607 8722 11633
rect 8694 11601 8722 11607
rect 8750 11634 8778 11639
rect 8358 11577 8386 11583
rect 8358 11551 8359 11577
rect 8385 11551 8386 11577
rect 8358 11130 8386 11551
rect 8414 11186 8442 11191
rect 8414 11139 8442 11158
rect 8750 11186 8778 11606
rect 8750 11139 8778 11158
rect 8806 11577 8834 11583
rect 8806 11551 8807 11577
rect 8833 11551 8834 11577
rect 8358 11097 8386 11102
rect 8078 10906 8106 10911
rect 7966 10905 8106 10906
rect 7966 10879 8079 10905
rect 8105 10879 8106 10905
rect 7966 10878 8106 10879
rect 7742 10817 7770 10822
rect 8022 10793 8050 10799
rect 8022 10767 8023 10793
rect 8049 10767 8050 10793
rect 8022 10458 8050 10767
rect 8022 10411 8050 10430
rect 7798 10345 7826 10351
rect 7798 10319 7799 10345
rect 7825 10319 7826 10345
rect 7798 10178 7826 10319
rect 7798 10150 7994 10178
rect 7350 10039 7351 10065
rect 7377 10039 7378 10065
rect 7350 10033 7378 10039
rect 7406 10066 7490 10094
rect 7518 10066 7546 10071
rect 7798 10066 7826 10071
rect 6790 10009 6818 10015
rect 6790 9983 6791 10009
rect 6817 9983 6818 10009
rect 6398 9954 6426 9959
rect 6118 9753 6146 9758
rect 6174 9953 6426 9954
rect 6174 9927 6399 9953
rect 6425 9927 6426 9953
rect 6174 9926 6426 9927
rect 6790 9954 6818 9983
rect 7014 10010 7042 10015
rect 7014 9954 7042 9982
rect 7238 10009 7266 10015
rect 7238 9983 7239 10009
rect 7265 9983 7266 10009
rect 6790 9953 7042 9954
rect 6790 9927 7015 9953
rect 7041 9927 7042 9953
rect 6790 9926 7042 9927
rect 6174 9729 6202 9926
rect 6398 9921 6426 9926
rect 6734 9786 6762 9791
rect 6762 9758 6818 9786
rect 6734 9753 6762 9758
rect 6174 9703 6175 9729
rect 6201 9703 6202 9729
rect 6174 9697 6202 9703
rect 6790 9729 6818 9758
rect 6790 9703 6791 9729
rect 6817 9703 6818 9729
rect 6790 9697 6818 9703
rect 6230 9674 6258 9679
rect 6230 9627 6258 9646
rect 6846 9562 6874 9567
rect 6846 9561 6930 9562
rect 6846 9535 6847 9561
rect 6873 9535 6930 9561
rect 6846 9534 6930 9535
rect 6846 9529 6874 9534
rect 6790 9506 6818 9511
rect 6734 9505 6818 9506
rect 6734 9479 6791 9505
rect 6817 9479 6818 9505
rect 6734 9478 6818 9479
rect 2142 9226 2170 9231
rect 2142 9179 2170 9198
rect 6230 9226 6258 9231
rect 6230 9179 6258 9198
rect 6622 9225 6650 9231
rect 6622 9199 6623 9225
rect 6649 9199 6650 9225
rect 5166 9170 5194 9175
rect 966 9114 994 9119
rect 966 9067 994 9086
rect 2238 9030 2370 9035
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2238 8997 2370 9002
rect 5166 8778 5194 9142
rect 6622 9170 6650 9199
rect 6622 9137 6650 9142
rect 5166 8745 5194 8750
rect 6734 8554 6762 9478
rect 6790 9473 6818 9478
rect 6902 9282 6930 9534
rect 6790 9225 6818 9231
rect 6790 9199 6791 9225
rect 6817 9199 6818 9225
rect 6790 8945 6818 9199
rect 6846 9226 6874 9231
rect 6846 9179 6874 9198
rect 6902 9225 6930 9254
rect 6902 9199 6903 9225
rect 6929 9199 6930 9225
rect 6902 9193 6930 9199
rect 6958 9394 6986 9399
rect 6790 8919 6791 8945
rect 6817 8919 6818 8945
rect 6790 8913 6818 8919
rect 6790 8778 6818 8783
rect 6790 8731 6818 8750
rect 6846 8778 6874 8783
rect 6958 8778 6986 9366
rect 7014 9170 7042 9926
rect 7182 9953 7210 9959
rect 7182 9927 7183 9953
rect 7209 9927 7210 9953
rect 7182 9674 7210 9927
rect 7182 9641 7210 9646
rect 7182 9394 7210 9399
rect 7238 9394 7266 9983
rect 7406 10010 7434 10066
rect 7518 10065 7826 10066
rect 7518 10039 7519 10065
rect 7545 10039 7799 10065
rect 7825 10039 7826 10065
rect 7518 10038 7826 10039
rect 7518 10033 7546 10038
rect 7798 10033 7826 10038
rect 7910 10066 7938 10071
rect 7406 9977 7434 9982
rect 7630 9897 7658 9903
rect 7630 9871 7631 9897
rect 7657 9871 7658 9897
rect 7630 9674 7658 9871
rect 7686 9898 7714 9903
rect 7686 9851 7714 9870
rect 7630 9641 7658 9646
rect 7574 9618 7602 9623
rect 7574 9571 7602 9590
rect 7210 9366 7266 9394
rect 7406 9505 7434 9511
rect 7406 9479 7407 9505
rect 7433 9479 7434 9505
rect 7182 9361 7210 9366
rect 7406 9282 7434 9479
rect 7854 9338 7882 9343
rect 7910 9338 7938 10038
rect 7966 10009 7994 10150
rect 7966 9983 7967 10009
rect 7993 9983 7994 10009
rect 7966 9618 7994 9983
rect 7966 9585 7994 9590
rect 7854 9337 7938 9338
rect 7854 9311 7855 9337
rect 7881 9311 7938 9337
rect 7854 9310 7938 9311
rect 7966 9506 7994 9511
rect 7966 9337 7994 9478
rect 7966 9311 7967 9337
rect 7993 9311 7994 9337
rect 7854 9305 7882 9310
rect 7966 9305 7994 9311
rect 7182 9254 7434 9282
rect 8078 9282 8106 10878
rect 8246 10794 8274 10934
rect 8134 10793 8274 10794
rect 8134 10767 8247 10793
rect 8273 10767 8274 10793
rect 8134 10766 8274 10767
rect 8134 10401 8162 10766
rect 8246 10761 8274 10766
rect 8526 11073 8554 11079
rect 8526 11047 8527 11073
rect 8553 11047 8554 11073
rect 8526 10794 8554 11047
rect 8526 10761 8554 10766
rect 8694 10850 8722 10855
rect 8806 10850 8834 11551
rect 8918 11578 8946 12222
rect 9142 11970 9170 12334
rect 9646 12361 9674 12446
rect 9982 12417 10010 12446
rect 9982 12391 9983 12417
rect 10009 12391 10010 12417
rect 9982 12385 10010 12391
rect 9646 12335 9647 12361
rect 9673 12335 9674 12361
rect 9646 12329 9674 12335
rect 9142 11942 9282 11970
rect 9086 11690 9114 11695
rect 9086 11643 9114 11662
rect 8974 11578 9002 11583
rect 8918 11577 9002 11578
rect 8918 11551 8975 11577
rect 9001 11551 9002 11577
rect 8918 11550 9002 11551
rect 8862 11074 8890 11079
rect 8918 11074 8946 11550
rect 8974 11545 9002 11550
rect 8974 11465 9002 11471
rect 8974 11439 8975 11465
rect 9001 11439 9002 11465
rect 8974 11298 9002 11439
rect 8974 11265 9002 11270
rect 8862 11073 8946 11074
rect 8862 11047 8863 11073
rect 8889 11047 8946 11073
rect 8862 11046 8946 11047
rect 9086 11186 9114 11191
rect 8862 10906 8890 11046
rect 8862 10873 8890 10878
rect 8694 10849 8834 10850
rect 8694 10823 8695 10849
rect 8721 10823 8834 10849
rect 8694 10822 8834 10823
rect 8134 10375 8135 10401
rect 8161 10375 8162 10401
rect 8134 10369 8162 10375
rect 8694 10122 8722 10822
rect 8862 10794 8890 10799
rect 8358 10066 8386 10071
rect 8358 10019 8386 10038
rect 8694 10010 8722 10094
rect 8750 10766 8862 10794
rect 8890 10766 9058 10794
rect 8750 10121 8778 10766
rect 8862 10747 8890 10766
rect 9030 10458 9058 10766
rect 9086 10514 9114 11158
rect 9198 11186 9226 11191
rect 9198 11139 9226 11158
rect 9142 11130 9170 11135
rect 9142 11083 9170 11102
rect 9254 10793 9282 11942
rect 10150 11802 10178 11807
rect 9918 11774 10050 11779
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 9918 11741 10050 11746
rect 10094 11634 10122 11639
rect 10150 11634 10178 11774
rect 10094 11633 10178 11634
rect 10094 11607 10095 11633
rect 10121 11607 10178 11633
rect 10094 11606 10178 11607
rect 10094 11601 10122 11606
rect 9422 11186 9450 11191
rect 10094 11186 10122 11191
rect 9422 11185 9506 11186
rect 9422 11159 9423 11185
rect 9449 11159 9506 11185
rect 9422 11158 9506 11159
rect 9422 11153 9450 11158
rect 9478 10962 9506 11158
rect 9310 10850 9338 10855
rect 9338 10822 9394 10850
rect 9310 10803 9338 10822
rect 9254 10767 9255 10793
rect 9281 10767 9282 10793
rect 9254 10761 9282 10767
rect 9142 10514 9170 10519
rect 9086 10513 9170 10514
rect 9086 10487 9143 10513
rect 9169 10487 9170 10513
rect 9086 10486 9170 10487
rect 9030 10457 9114 10458
rect 9030 10431 9031 10457
rect 9057 10431 9114 10457
rect 9030 10430 9114 10431
rect 9030 10425 9058 10430
rect 8750 10095 8751 10121
rect 8777 10095 8778 10121
rect 8750 10089 8778 10095
rect 8918 10122 8946 10127
rect 8862 10066 8890 10071
rect 8862 10019 8890 10038
rect 8694 9982 8834 10010
rect 8414 9898 8442 9903
rect 8414 9897 8666 9898
rect 8414 9871 8415 9897
rect 8441 9871 8666 9897
rect 8414 9870 8666 9871
rect 8414 9865 8442 9870
rect 8470 9561 8498 9567
rect 8470 9535 8471 9561
rect 8497 9535 8498 9561
rect 8358 9338 8386 9343
rect 8358 9291 8386 9310
rect 8302 9282 8330 9287
rect 8078 9281 8330 9282
rect 8078 9255 8079 9281
rect 8105 9255 8303 9281
rect 8329 9255 8330 9281
rect 8078 9254 8330 9255
rect 7014 9137 7042 9142
rect 7070 9226 7098 9231
rect 7182 9226 7210 9254
rect 8078 9249 8106 9254
rect 8302 9249 8330 9254
rect 7070 9225 7210 9226
rect 7070 9199 7071 9225
rect 7097 9199 7210 9225
rect 7070 9198 7210 9199
rect 7798 9226 7826 9231
rect 6846 8777 6986 8778
rect 6846 8751 6847 8777
rect 6873 8751 6986 8777
rect 6846 8750 6986 8751
rect 6734 8521 6762 8526
rect 6566 8498 6594 8503
rect 2142 8442 2170 8447
rect 2142 8395 2170 8414
rect 5502 8442 5530 8447
rect 966 8329 994 8335
rect 966 8303 967 8329
rect 993 8303 994 8329
rect 966 8106 994 8303
rect 2238 8246 2370 8251
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2238 8213 2370 8218
rect 966 8073 994 8078
rect 5502 7601 5530 8414
rect 6566 7713 6594 8470
rect 6846 8441 6874 8750
rect 7014 8554 7042 8559
rect 7070 8554 7098 9198
rect 7798 9179 7826 9198
rect 7238 9170 7266 9175
rect 7294 9170 7322 9175
rect 7266 9169 7322 9170
rect 7266 9143 7295 9169
rect 7321 9143 7322 9169
rect 7266 9142 7322 9143
rect 7126 8554 7154 8559
rect 7070 8526 7126 8554
rect 7014 8507 7042 8526
rect 7126 8497 7154 8526
rect 7126 8471 7127 8497
rect 7153 8471 7154 8497
rect 7126 8465 7154 8471
rect 6846 8415 6847 8441
rect 6873 8415 6874 8441
rect 6846 8218 6874 8415
rect 6902 8441 6930 8447
rect 6902 8415 6903 8441
rect 6929 8415 6930 8441
rect 6902 8386 6930 8415
rect 6958 8442 6986 8447
rect 6958 8395 6986 8414
rect 6902 8353 6930 8358
rect 6846 8185 6874 8190
rect 7126 8106 7154 8111
rect 7126 8059 7154 8078
rect 6566 7687 6567 7713
rect 6593 7687 6594 7713
rect 6566 7681 6594 7687
rect 6790 8049 6818 8055
rect 6790 8023 6791 8049
rect 6817 8023 6818 8049
rect 6790 7658 6818 8023
rect 6958 7658 6986 7663
rect 6790 7657 7042 7658
rect 6790 7631 6959 7657
rect 6985 7631 7042 7657
rect 6790 7630 7042 7631
rect 6958 7625 6986 7630
rect 5502 7575 5503 7601
rect 5529 7575 5530 7601
rect 5502 7569 5530 7575
rect 7014 7546 7042 7630
rect 7182 7601 7210 7607
rect 7182 7575 7183 7601
rect 7209 7575 7210 7601
rect 7182 7546 7210 7575
rect 7238 7546 7266 9142
rect 7294 9137 7322 9142
rect 8414 9170 8442 9175
rect 8358 9113 8386 9119
rect 8358 9087 8359 9113
rect 8385 9087 8386 9113
rect 8358 9002 8386 9087
rect 8358 8969 8386 8974
rect 8414 8834 8442 9142
rect 8358 8806 8442 8834
rect 8302 8778 8330 8783
rect 8302 8731 8330 8750
rect 7350 8722 7378 8727
rect 7350 8553 7378 8694
rect 8246 8722 8274 8727
rect 8246 8675 8274 8694
rect 7854 8666 7882 8671
rect 7350 8527 7351 8553
rect 7377 8527 7378 8553
rect 7350 8521 7378 8527
rect 7686 8610 7714 8615
rect 7462 8498 7490 8503
rect 7462 8451 7490 8470
rect 7294 8442 7322 8447
rect 7294 8395 7322 8414
rect 7686 8441 7714 8582
rect 7686 8415 7687 8441
rect 7713 8415 7714 8441
rect 7686 8409 7714 8415
rect 7742 8554 7770 8559
rect 7294 7546 7322 7551
rect 7014 7518 7294 7546
rect 2238 7462 2370 7467
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2238 7429 2370 7434
rect 7014 6873 7042 7518
rect 7294 7513 7322 7518
rect 7742 7378 7770 8526
rect 7854 8553 7882 8638
rect 7854 8527 7855 8553
rect 7881 8527 7882 8553
rect 7854 8521 7882 8527
rect 8246 8497 8274 8503
rect 8246 8471 8247 8497
rect 8273 8471 8274 8497
rect 7966 8442 7994 8447
rect 8134 8442 8162 8447
rect 7966 8441 8162 8442
rect 7966 8415 7967 8441
rect 7993 8415 8135 8441
rect 8161 8415 8162 8441
rect 7966 8414 8162 8415
rect 7966 8409 7994 8414
rect 8134 8409 8162 8414
rect 7798 8385 7826 8391
rect 7798 8359 7799 8385
rect 7825 8359 7826 8385
rect 7798 8106 7826 8359
rect 7798 8073 7826 8078
rect 8190 8106 8218 8111
rect 8246 8106 8274 8471
rect 8302 8498 8330 8503
rect 8358 8498 8386 8806
rect 8414 8722 8442 8727
rect 8414 8675 8442 8694
rect 8302 8497 8386 8498
rect 8302 8471 8303 8497
rect 8329 8471 8386 8497
rect 8302 8470 8386 8471
rect 8302 8465 8330 8470
rect 8190 8105 8274 8106
rect 8190 8079 8191 8105
rect 8217 8079 8274 8105
rect 8190 8078 8274 8079
rect 8190 8073 8218 8078
rect 7966 7378 7994 7383
rect 7742 7377 7994 7378
rect 7742 7351 7967 7377
rect 7993 7351 7994 7377
rect 7742 7350 7994 7351
rect 7966 7345 7994 7350
rect 8078 7378 8106 7383
rect 8078 7331 8106 7350
rect 8190 7266 8218 7271
rect 8190 7219 8218 7238
rect 7350 7210 7378 7215
rect 7350 6929 7378 7182
rect 7910 7210 7938 7215
rect 7910 7163 7938 7182
rect 7350 6903 7351 6929
rect 7377 6903 7378 6929
rect 7350 6897 7378 6903
rect 7014 6847 7015 6873
rect 7041 6847 7042 6873
rect 7014 6841 7042 6847
rect 2238 6678 2370 6683
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2238 6645 2370 6650
rect 2238 5894 2370 5899
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2238 5861 2370 5866
rect 2238 5110 2370 5115
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2238 5077 2370 5082
rect 2238 4326 2370 4331
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2238 4293 2370 4298
rect 8246 4214 8274 8078
rect 8414 8106 8442 8111
rect 8470 8106 8498 9535
rect 8638 9282 8666 9870
rect 8694 9897 8722 9903
rect 8694 9871 8695 9897
rect 8721 9871 8722 9897
rect 8694 9338 8722 9871
rect 8694 9305 8722 9310
rect 8638 9225 8666 9254
rect 8638 9199 8639 9225
rect 8665 9199 8666 9225
rect 8638 9193 8666 9199
rect 8806 9225 8834 9982
rect 8806 9199 8807 9225
rect 8833 9199 8834 9225
rect 8806 9193 8834 9199
rect 8750 9169 8778 9175
rect 8750 9143 8751 9169
rect 8777 9143 8778 9169
rect 8582 9002 8610 9007
rect 8582 8833 8610 8974
rect 8582 8807 8583 8833
rect 8609 8807 8610 8833
rect 8582 8801 8610 8807
rect 8414 8105 8498 8106
rect 8414 8079 8415 8105
rect 8441 8079 8498 8105
rect 8414 8078 8498 8079
rect 8358 7546 8386 7551
rect 8414 7546 8442 8078
rect 8386 7518 8442 7546
rect 8302 6818 8330 6823
rect 8358 6818 8386 7518
rect 8750 7378 8778 9143
rect 8918 8722 8946 10094
rect 9086 10121 9114 10430
rect 9086 10095 9087 10121
rect 9113 10095 9114 10121
rect 9086 10089 9114 10095
rect 9142 10066 9170 10486
rect 9310 10514 9338 10519
rect 9310 10467 9338 10486
rect 9142 10033 9170 10038
rect 9030 10010 9058 10015
rect 9030 9506 9058 9982
rect 9198 10010 9226 10015
rect 9366 10010 9394 10822
rect 9478 10401 9506 10934
rect 9478 10375 9479 10401
rect 9505 10375 9506 10401
rect 9478 10369 9506 10375
rect 9534 11073 9562 11079
rect 9534 11047 9535 11073
rect 9561 11047 9562 11073
rect 9534 10962 9562 11047
rect 9918 10990 10050 10995
rect 9590 10962 9618 10967
rect 9534 10934 9590 10962
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 9918 10957 10050 10962
rect 9534 10290 9562 10934
rect 9590 10929 9618 10934
rect 9814 10849 9842 10855
rect 9814 10823 9815 10849
rect 9841 10823 9842 10849
rect 9758 10458 9786 10463
rect 9814 10458 9842 10823
rect 9758 10457 9842 10458
rect 9758 10431 9759 10457
rect 9785 10431 9842 10457
rect 9758 10430 9842 10431
rect 9758 10425 9786 10430
rect 9198 10009 9282 10010
rect 9198 9983 9199 10009
rect 9225 9983 9282 10009
rect 9198 9982 9282 9983
rect 9198 9977 9226 9982
rect 9030 9473 9058 9478
rect 9254 9506 9282 9982
rect 9366 9977 9394 9982
rect 9478 10262 9562 10290
rect 8974 9338 9002 9343
rect 9198 9338 9226 9343
rect 9002 9310 9058 9338
rect 8974 9305 9002 9310
rect 8974 9225 9002 9231
rect 8974 9199 8975 9225
rect 9001 9199 9002 9225
rect 8974 9170 9002 9199
rect 8974 9137 9002 9142
rect 9030 8777 9058 9310
rect 9198 9291 9226 9310
rect 9254 9281 9282 9478
rect 9254 9255 9255 9281
rect 9281 9255 9282 9281
rect 9254 9249 9282 9255
rect 9198 9113 9226 9119
rect 9198 9087 9199 9113
rect 9225 9087 9226 9113
rect 9030 8751 9031 8777
rect 9057 8751 9058 8777
rect 9030 8745 9058 8751
rect 9142 8946 9170 8951
rect 9198 8946 9226 9087
rect 9142 8945 9226 8946
rect 9142 8919 9143 8945
rect 9169 8919 9226 8945
rect 9142 8918 9226 8919
rect 8918 8689 8946 8694
rect 9086 8721 9114 8727
rect 9086 8695 9087 8721
rect 9113 8695 9114 8721
rect 9086 8554 9114 8695
rect 9142 8610 9170 8918
rect 9142 8577 9170 8582
rect 9366 8778 9394 8783
rect 9086 8521 9114 8526
rect 9198 7658 9226 7663
rect 8414 7321 8442 7327
rect 8414 7295 8415 7321
rect 8441 7295 8442 7321
rect 8414 7266 8442 7295
rect 8526 7322 8554 7327
rect 8526 7275 8554 7294
rect 8694 7321 8722 7327
rect 8694 7295 8695 7321
rect 8721 7295 8722 7321
rect 8414 7233 8442 7238
rect 8330 6790 8386 6818
rect 8414 7153 8442 7159
rect 8414 7127 8415 7153
rect 8441 7127 8442 7153
rect 8414 6817 8442 7127
rect 8414 6791 8415 6817
rect 8441 6791 8442 6817
rect 8302 6481 8330 6790
rect 8302 6455 8303 6481
rect 8329 6455 8330 6481
rect 8302 6449 8330 6455
rect 8190 4186 8274 4214
rect 8414 4214 8442 6791
rect 8638 6538 8666 6543
rect 8694 6538 8722 7295
rect 8750 7209 8778 7350
rect 9030 7657 9226 7658
rect 9030 7631 9199 7657
rect 9225 7631 9226 7657
rect 9030 7630 9226 7631
rect 9030 7601 9058 7630
rect 9198 7625 9226 7630
rect 9030 7575 9031 7601
rect 9057 7575 9058 7601
rect 8750 7183 8751 7209
rect 8777 7183 8778 7209
rect 8750 7177 8778 7183
rect 8862 7210 8890 7215
rect 8862 7163 8890 7182
rect 8750 6818 8778 6823
rect 8750 6771 8778 6790
rect 9030 6818 9058 7575
rect 9366 7322 9394 8750
rect 9478 8274 9506 10262
rect 9702 10009 9730 10015
rect 9702 9983 9703 10009
rect 9729 9983 9730 10009
rect 9534 9954 9562 9959
rect 9702 9954 9730 9983
rect 9562 9926 9730 9954
rect 9534 9907 9562 9926
rect 9590 9338 9618 9343
rect 9590 9291 9618 9310
rect 9814 9338 9842 10430
rect 10094 10401 10122 11158
rect 10094 10375 10095 10401
rect 10121 10375 10122 10401
rect 10094 10369 10122 10375
rect 9918 10206 10050 10211
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 9918 10173 10050 10178
rect 10038 10066 10066 10071
rect 10038 9617 10066 10038
rect 10038 9591 10039 9617
rect 10065 9591 10066 9617
rect 10038 9585 10066 9591
rect 9918 9422 10050 9427
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 9918 9389 10050 9394
rect 9814 9305 9842 9310
rect 9982 9338 10010 9343
rect 10150 9338 10178 11606
rect 10206 11577 10234 11583
rect 10206 11551 10207 11577
rect 10233 11551 10234 11577
rect 10206 10514 10234 11551
rect 10262 11298 10290 12671
rect 10318 12698 10346 12703
rect 10318 12651 10346 12670
rect 10766 12306 10794 13399
rect 10654 12082 10682 12087
rect 10654 12035 10682 12054
rect 10654 11577 10682 11583
rect 10654 11551 10655 11577
rect 10681 11551 10682 11577
rect 10486 11522 10514 11527
rect 10486 11521 10570 11522
rect 10486 11495 10487 11521
rect 10513 11495 10570 11521
rect 10486 11494 10570 11495
rect 10486 11489 10514 11494
rect 10318 11298 10346 11317
rect 10262 11270 10318 11298
rect 10318 11265 10346 11270
rect 10318 11186 10346 11191
rect 10318 11139 10346 11158
rect 10206 10481 10234 10486
rect 10542 11130 10570 11494
rect 10654 11186 10682 11551
rect 10766 11354 10794 12278
rect 10822 12641 10850 13510
rect 10934 13454 10962 18607
rect 10990 13538 11018 13543
rect 10990 13537 11410 13538
rect 10990 13511 10991 13537
rect 11017 13511 11410 13537
rect 10990 13510 11410 13511
rect 10990 13505 11018 13510
rect 10934 13426 11074 13454
rect 11046 12698 11074 13426
rect 11382 13257 11410 13510
rect 11774 13454 11802 18999
rect 12838 19025 12866 19031
rect 12838 18999 12839 19025
rect 12865 18999 12866 19025
rect 12838 15974 12866 18999
rect 17598 18438 17730 18443
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17598 18405 17730 18410
rect 17598 17654 17730 17659
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17598 17621 17730 17626
rect 17598 16870 17730 16875
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17598 16837 17730 16842
rect 17598 16086 17730 16091
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17598 16053 17730 16058
rect 12838 15946 12978 15974
rect 12558 13481 12586 13487
rect 12558 13455 12559 13481
rect 12585 13455 12586 13481
rect 12558 13454 12586 13455
rect 11494 13426 11802 13454
rect 12334 13426 12586 13454
rect 12614 13482 12642 13487
rect 12614 13435 12642 13454
rect 11494 13258 11522 13426
rect 11382 13231 11383 13257
rect 11409 13231 11410 13257
rect 11382 13225 11410 13231
rect 11438 13257 11522 13258
rect 11438 13231 11495 13257
rect 11521 13231 11522 13257
rect 11438 13230 11522 13231
rect 11270 13090 11298 13095
rect 11438 13090 11466 13230
rect 11494 13225 11522 13230
rect 11550 13258 11578 13263
rect 11550 13201 11578 13230
rect 12334 13258 12362 13426
rect 11550 13175 11551 13201
rect 11577 13175 11578 13201
rect 11550 13169 11578 13175
rect 12278 13202 12306 13207
rect 12278 13155 12306 13174
rect 12334 13201 12362 13230
rect 12334 13175 12335 13201
rect 12361 13175 12362 13201
rect 12334 13169 12362 13175
rect 12726 13425 12754 13431
rect 12726 13399 12727 13425
rect 12753 13399 12754 13425
rect 11270 13089 11466 13090
rect 11270 13063 11271 13089
rect 11297 13063 11466 13089
rect 11270 13062 11466 13063
rect 11606 13146 11634 13151
rect 11270 13057 11298 13062
rect 11550 12754 11578 12759
rect 11606 12754 11634 13118
rect 11830 13146 11858 13151
rect 12166 13146 12194 13151
rect 11830 13099 11858 13118
rect 11942 13145 12194 13146
rect 11942 13119 12167 13145
rect 12193 13119 12194 13145
rect 11942 13118 12194 13119
rect 11550 12753 11634 12754
rect 11550 12727 11551 12753
rect 11577 12727 11634 12753
rect 11550 12726 11634 12727
rect 11550 12721 11578 12726
rect 11886 12698 11914 12703
rect 10822 12615 10823 12641
rect 10849 12615 10850 12641
rect 10822 12082 10850 12615
rect 10878 12642 10906 12647
rect 10878 12595 10906 12614
rect 10934 12641 10962 12647
rect 10934 12615 10935 12641
rect 10961 12615 10962 12641
rect 10934 12586 10962 12615
rect 10934 12553 10962 12558
rect 11046 12305 11074 12670
rect 11662 12697 11914 12698
rect 11662 12671 11887 12697
rect 11913 12671 11914 12697
rect 11662 12670 11914 12671
rect 11550 12586 11578 12591
rect 11578 12558 11634 12586
rect 11550 12553 11578 12558
rect 11046 12279 11047 12305
rect 11073 12279 11074 12305
rect 11046 12273 11074 12279
rect 11606 12473 11634 12558
rect 11606 12447 11607 12473
rect 11633 12447 11634 12473
rect 10822 12054 10906 12082
rect 10822 11970 10850 11975
rect 10878 11970 10906 12054
rect 10934 11970 10962 11975
rect 10878 11969 10962 11970
rect 10878 11943 10935 11969
rect 10961 11943 10962 11969
rect 10878 11942 10962 11943
rect 10822 11923 10850 11942
rect 10934 11802 10962 11942
rect 10934 11769 10962 11774
rect 11494 11970 11522 11975
rect 10654 11139 10682 11158
rect 10710 11326 10794 11354
rect 10878 11521 10906 11527
rect 10878 11495 10879 11521
rect 10905 11495 10906 11521
rect 10542 10794 10570 11102
rect 10598 10794 10626 10799
rect 10542 10793 10626 10794
rect 10542 10767 10599 10793
rect 10625 10767 10626 10793
rect 10542 10766 10626 10767
rect 10262 10290 10290 10295
rect 10262 10289 10346 10290
rect 10262 10263 10263 10289
rect 10289 10263 10346 10289
rect 10262 10262 10346 10263
rect 10262 10257 10290 10262
rect 10318 10234 10346 10262
rect 10262 10010 10290 10015
rect 9982 9291 10010 9310
rect 10038 9310 10178 9338
rect 10206 9674 10234 9679
rect 9758 9281 9786 9287
rect 9758 9255 9759 9281
rect 9785 9255 9786 9281
rect 9758 9058 9786 9255
rect 9926 9282 9954 9287
rect 9926 9235 9954 9254
rect 9982 9114 10010 9119
rect 9982 9067 10010 9086
rect 9590 9030 9758 9058
rect 9534 8834 9562 8839
rect 9534 8787 9562 8806
rect 9590 8666 9618 9030
rect 9758 9025 9786 9030
rect 9926 8890 9954 8895
rect 9478 8241 9506 8246
rect 9534 8638 9618 8666
rect 9646 8889 9954 8890
rect 9646 8863 9927 8889
rect 9953 8863 9954 8889
rect 9646 8862 9954 8863
rect 9366 7265 9394 7294
rect 9366 7239 9367 7265
rect 9393 7239 9394 7265
rect 9366 7233 9394 7239
rect 9422 7210 9450 7215
rect 9534 7210 9562 8638
rect 9646 8553 9674 8862
rect 9926 8857 9954 8862
rect 9982 8834 10010 8839
rect 10038 8834 10066 9310
rect 9982 8833 10066 8834
rect 9982 8807 9983 8833
rect 10009 8807 10066 8833
rect 9982 8806 10066 8807
rect 9982 8801 10010 8806
rect 9758 8777 9786 8783
rect 9758 8751 9759 8777
rect 9785 8751 9786 8777
rect 9702 8722 9730 8727
rect 9758 8722 9786 8751
rect 9870 8722 9898 8727
rect 9730 8694 9786 8722
rect 9814 8721 9898 8722
rect 9814 8695 9871 8721
rect 9897 8695 9898 8721
rect 9814 8694 9898 8695
rect 9702 8689 9730 8694
rect 9646 8527 9647 8553
rect 9673 8527 9674 8553
rect 9646 8521 9674 8527
rect 9758 8554 9786 8559
rect 9758 8507 9786 8526
rect 9702 8385 9730 8391
rect 9702 8359 9703 8385
rect 9729 8359 9730 8385
rect 9590 7714 9618 7719
rect 9702 7714 9730 8359
rect 9814 8274 9842 8694
rect 9870 8689 9898 8694
rect 9918 8638 10050 8643
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 9918 8605 10050 8610
rect 9982 8441 10010 8447
rect 9982 8415 9983 8441
rect 10009 8415 10010 8441
rect 9870 8274 9898 8279
rect 9814 8246 9870 8274
rect 9870 8241 9898 8246
rect 9982 8106 10010 8415
rect 9982 8073 10010 8078
rect 9918 7854 10050 7859
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 9918 7821 10050 7826
rect 9590 7713 9730 7714
rect 9590 7687 9591 7713
rect 9617 7687 9730 7713
rect 9590 7686 9730 7687
rect 9590 7681 9618 7686
rect 10206 7265 10234 9646
rect 10262 9281 10290 9982
rect 10262 9255 10263 9281
rect 10289 9255 10290 9281
rect 10262 9249 10290 9255
rect 10318 9281 10346 10206
rect 10318 9255 10319 9281
rect 10345 9255 10346 9281
rect 10318 7994 10346 9255
rect 10430 9226 10458 9231
rect 10430 9179 10458 9198
rect 10542 8834 10570 10766
rect 10598 10761 10626 10766
rect 10654 10738 10682 10743
rect 10654 10691 10682 10710
rect 10710 10514 10738 11326
rect 10878 11298 10906 11495
rect 10878 11270 11186 11298
rect 10766 11242 10794 11247
rect 10766 11195 10794 11214
rect 11102 11186 11130 11191
rect 11102 11139 11130 11158
rect 11158 11129 11186 11270
rect 11158 11103 11159 11129
rect 11185 11103 11186 11129
rect 10934 11074 10962 11079
rect 10934 11073 11074 11074
rect 10934 11047 10935 11073
rect 10961 11047 11074 11073
rect 10934 11046 11074 11047
rect 10934 11041 10962 11046
rect 10990 10962 11018 10967
rect 10934 10906 10962 10911
rect 10934 10859 10962 10878
rect 10822 10793 10850 10799
rect 10822 10767 10823 10793
rect 10849 10767 10850 10793
rect 10766 10514 10794 10519
rect 10710 10513 10794 10514
rect 10710 10487 10767 10513
rect 10793 10487 10794 10513
rect 10710 10486 10794 10487
rect 10654 9506 10682 9511
rect 10654 9459 10682 9478
rect 10654 9226 10682 9231
rect 10710 9226 10738 10486
rect 10766 10481 10794 10486
rect 10822 10514 10850 10767
rect 10878 10737 10906 10743
rect 10878 10711 10879 10737
rect 10905 10711 10906 10737
rect 10878 10682 10906 10711
rect 10878 10649 10906 10654
rect 10822 10481 10850 10486
rect 10990 10458 11018 10934
rect 10990 10401 11018 10430
rect 10990 10375 10991 10401
rect 11017 10375 11018 10401
rect 10990 10369 11018 10375
rect 10822 10345 10850 10351
rect 10822 10319 10823 10345
rect 10849 10319 10850 10345
rect 10766 10289 10794 10295
rect 10766 10263 10767 10289
rect 10793 10263 10794 10289
rect 10766 10234 10794 10263
rect 10822 10290 10850 10319
rect 10822 10257 10850 10262
rect 10766 10201 10794 10206
rect 10822 10178 10850 10183
rect 10822 9561 10850 10150
rect 10822 9535 10823 9561
rect 10849 9535 10850 9561
rect 10822 9529 10850 9535
rect 10990 9898 11018 9903
rect 10990 9506 11018 9870
rect 11046 9618 11074 11046
rect 11158 10962 11186 11103
rect 11158 10929 11186 10934
rect 11382 11073 11410 11079
rect 11382 11047 11383 11073
rect 11409 11047 11410 11073
rect 11382 10906 11410 11047
rect 11494 11074 11522 11942
rect 11550 11522 11578 11527
rect 11550 11241 11578 11494
rect 11550 11215 11551 11241
rect 11577 11215 11578 11241
rect 11550 11209 11578 11215
rect 11606 11298 11634 12447
rect 11662 12473 11690 12670
rect 11886 12665 11914 12670
rect 11662 12447 11663 12473
rect 11689 12447 11690 12473
rect 11662 12441 11690 12447
rect 11718 12361 11746 12367
rect 11718 12335 11719 12361
rect 11745 12335 11746 12361
rect 11718 11970 11746 12335
rect 11942 12361 11970 13118
rect 12166 13113 12194 13118
rect 12614 13146 12642 13151
rect 12614 13099 12642 13118
rect 12726 12922 12754 13399
rect 12614 12894 12754 12922
rect 12950 13202 12978 15946
rect 17598 15302 17730 15307
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17598 15269 17730 15274
rect 17598 14518 17730 14523
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17598 14485 17730 14490
rect 18830 13929 18858 13935
rect 18830 13903 18831 13929
rect 18857 13903 18858 13929
rect 17598 13734 17730 13739
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17598 13701 17730 13706
rect 13566 13650 13594 13655
rect 12614 12417 12642 12894
rect 12950 12809 12978 13174
rect 13454 13537 13482 13543
rect 13454 13511 13455 13537
rect 13481 13511 13482 13537
rect 13454 13482 13482 13511
rect 13174 13146 13202 13151
rect 12950 12783 12951 12809
rect 12977 12783 12978 12809
rect 12950 12777 12978 12783
rect 13006 13089 13034 13095
rect 13006 13063 13007 13089
rect 13033 13063 13034 13089
rect 13006 12642 13034 13063
rect 13174 12866 13202 13118
rect 13174 12809 13202 12838
rect 13174 12783 13175 12809
rect 13201 12783 13202 12809
rect 13174 12777 13202 12783
rect 13454 13090 13482 13454
rect 13566 13481 13594 13622
rect 18830 13650 18858 13903
rect 18830 13617 18858 13622
rect 19950 13873 19978 13879
rect 19950 13847 19951 13873
rect 19977 13847 19978 13873
rect 13566 13455 13567 13481
rect 13593 13455 13594 13481
rect 13566 13449 13594 13455
rect 18942 13537 18970 13543
rect 18942 13511 18943 13537
rect 18969 13511 18970 13537
rect 18830 13146 18858 13151
rect 18830 13099 18858 13118
rect 13454 12753 13482 13062
rect 14126 13090 14154 13095
rect 14126 13043 14154 13062
rect 14462 13089 14490 13095
rect 14462 13063 14463 13089
rect 14489 13063 14490 13089
rect 14462 12866 14490 13063
rect 17598 12950 17730 12955
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17598 12917 17730 12922
rect 14490 12838 14658 12866
rect 14462 12833 14490 12838
rect 13454 12727 13455 12753
rect 13481 12727 13482 12753
rect 13454 12721 13482 12727
rect 13566 12698 13594 12703
rect 13566 12651 13594 12670
rect 12782 12614 13034 12642
rect 12782 12473 12810 12614
rect 12782 12447 12783 12473
rect 12809 12447 12810 12473
rect 12782 12441 12810 12447
rect 12614 12391 12615 12417
rect 12641 12391 12642 12417
rect 12614 12385 12642 12391
rect 12670 12417 12698 12423
rect 12670 12391 12671 12417
rect 12697 12391 12698 12417
rect 11942 12335 11943 12361
rect 11969 12335 11970 12361
rect 11942 12329 11970 12335
rect 11718 11937 11746 11942
rect 12670 11690 12698 12391
rect 12614 11662 12698 11690
rect 12894 11690 12922 11695
rect 12334 11578 12362 11583
rect 12334 11531 12362 11550
rect 11942 11522 11970 11527
rect 11942 11475 11970 11494
rect 11606 11185 11634 11270
rect 11606 11159 11607 11185
rect 11633 11159 11634 11185
rect 11606 11153 11634 11159
rect 11718 11354 11746 11359
rect 11494 11073 11634 11074
rect 11494 11047 11495 11073
rect 11521 11047 11634 11073
rect 11494 11046 11634 11047
rect 11494 11041 11522 11046
rect 11382 10878 11578 10906
rect 11158 10793 11186 10799
rect 11326 10794 11354 10799
rect 11158 10767 11159 10793
rect 11185 10767 11186 10793
rect 11102 10738 11130 10743
rect 11102 10122 11130 10710
rect 11102 9618 11130 10094
rect 11158 10290 11186 10767
rect 11158 10010 11186 10262
rect 11158 9977 11186 9982
rect 11214 10766 11326 10794
rect 11214 9786 11242 10766
rect 11326 10761 11354 10766
rect 11382 10793 11410 10799
rect 11382 10767 11383 10793
rect 11409 10767 11410 10793
rect 11382 10738 11410 10767
rect 11438 10794 11466 10813
rect 11438 10761 11466 10766
rect 11494 10793 11522 10799
rect 11494 10767 11495 10793
rect 11521 10767 11522 10793
rect 11382 10705 11410 10710
rect 11494 10682 11522 10767
rect 11494 10649 11522 10654
rect 11326 10345 11354 10351
rect 11326 10319 11327 10345
rect 11353 10319 11354 10345
rect 11326 10178 11354 10319
rect 11326 10145 11354 10150
rect 11382 10289 11410 10295
rect 11382 10263 11383 10289
rect 11409 10263 11410 10289
rect 11158 9758 11242 9786
rect 11326 10010 11354 10015
rect 11158 9674 11186 9758
rect 11158 9646 11298 9674
rect 11102 9590 11242 9618
rect 11046 9585 11074 9590
rect 10934 9478 11074 9506
rect 10654 9225 10738 9226
rect 10654 9199 10655 9225
rect 10681 9199 10738 9225
rect 10654 9198 10738 9199
rect 10766 9450 10794 9455
rect 10766 9225 10794 9422
rect 10934 9226 10962 9478
rect 11046 9450 11074 9478
rect 11158 9505 11186 9511
rect 11158 9479 11159 9505
rect 11185 9479 11186 9505
rect 11158 9450 11186 9479
rect 11046 9422 11186 9450
rect 10766 9199 10767 9225
rect 10793 9199 10794 9225
rect 10654 9193 10682 9198
rect 10766 9193 10794 9199
rect 10878 9198 10962 9226
rect 11158 9226 11186 9231
rect 10542 8801 10570 8806
rect 10878 9170 10906 9198
rect 10710 8106 10738 8111
rect 10710 8059 10738 8078
rect 10878 8049 10906 9142
rect 10990 9170 11018 9175
rect 10934 9113 10962 9119
rect 10934 9087 10935 9113
rect 10961 9087 10962 9113
rect 10934 8330 10962 9087
rect 10990 9058 11018 9142
rect 10990 9025 11018 9030
rect 11102 9169 11130 9175
rect 11102 9143 11103 9169
rect 11129 9143 11130 9169
rect 11102 8834 11130 9143
rect 11102 8801 11130 8806
rect 11158 8554 11186 9198
rect 11214 9225 11242 9590
rect 11214 9199 11215 9225
rect 11241 9199 11242 9225
rect 11214 9193 11242 9199
rect 11270 9225 11298 9646
rect 11326 9618 11354 9982
rect 11382 9898 11410 10263
rect 11494 10290 11522 10295
rect 11550 10290 11578 10878
rect 11494 10289 11578 10290
rect 11494 10263 11495 10289
rect 11521 10263 11578 10289
rect 11494 10262 11578 10263
rect 11494 10094 11522 10262
rect 11550 10178 11578 10183
rect 11606 10178 11634 11046
rect 11718 10905 11746 11326
rect 11830 11298 11858 11303
rect 11830 11251 11858 11270
rect 11774 11130 11802 11135
rect 11774 11083 11802 11102
rect 11830 11073 11858 11079
rect 11830 11047 11831 11073
rect 11857 11047 11858 11073
rect 11830 11018 11858 11047
rect 11830 10985 11858 10990
rect 12614 10962 12642 11662
rect 12894 11633 12922 11662
rect 12894 11607 12895 11633
rect 12921 11607 12922 11633
rect 12894 11601 12922 11607
rect 12670 11578 12698 11583
rect 13062 11578 13090 11597
rect 12698 11550 12866 11578
rect 12670 11531 12698 11550
rect 12838 11186 12866 11550
rect 13062 11545 13090 11550
rect 13230 11577 13258 11583
rect 13230 11551 13231 11577
rect 13257 11551 13258 11577
rect 13062 11466 13090 11471
rect 13062 11465 13202 11466
rect 13062 11439 13063 11465
rect 13089 11439 13202 11465
rect 13062 11438 13202 11439
rect 13062 11433 13090 11438
rect 13174 11242 13202 11438
rect 13230 11354 13258 11551
rect 13734 11577 13762 11583
rect 13734 11551 13735 11577
rect 13761 11551 13762 11577
rect 13230 11321 13258 11326
rect 13342 11521 13370 11527
rect 13342 11495 13343 11521
rect 13369 11495 13370 11521
rect 13230 11242 13258 11247
rect 13174 11241 13258 11242
rect 13174 11215 13231 11241
rect 13257 11215 13258 11241
rect 13174 11214 13258 11215
rect 13230 11209 13258 11214
rect 12838 11185 12978 11186
rect 12838 11159 12839 11185
rect 12865 11159 12978 11185
rect 12838 11158 12978 11159
rect 12838 11153 12866 11158
rect 12614 10929 12642 10934
rect 11718 10879 11719 10905
rect 11745 10879 11746 10905
rect 11718 10873 11746 10879
rect 12950 10793 12978 11158
rect 13342 10849 13370 11495
rect 13342 10823 13343 10849
rect 13369 10823 13370 10849
rect 13342 10817 13370 10823
rect 13398 11465 13426 11471
rect 13398 11439 13399 11465
rect 13425 11439 13426 11465
rect 12950 10767 12951 10793
rect 12977 10767 12978 10793
rect 12950 10457 12978 10767
rect 13398 10794 13426 11439
rect 13398 10761 13426 10766
rect 12950 10431 12951 10457
rect 12977 10431 12978 10457
rect 11578 10150 11634 10178
rect 11774 10401 11802 10407
rect 11774 10375 11775 10401
rect 11801 10375 11802 10401
rect 11550 10145 11578 10150
rect 11494 10066 11690 10094
rect 11382 9865 11410 9870
rect 11606 9618 11634 9623
rect 11326 9617 11634 9618
rect 11326 9591 11327 9617
rect 11353 9591 11607 9617
rect 11633 9591 11634 9617
rect 11326 9590 11634 9591
rect 11326 9585 11354 9590
rect 11606 9585 11634 9590
rect 11494 9506 11522 9511
rect 11270 9199 11271 9225
rect 11297 9199 11298 9225
rect 11270 9002 11298 9199
rect 11270 8969 11298 8974
rect 11438 9505 11522 9506
rect 11438 9479 11495 9505
rect 11521 9479 11522 9505
rect 11438 9478 11522 9479
rect 11214 8554 11242 8559
rect 10934 8297 10962 8302
rect 11046 8553 11242 8554
rect 11046 8527 11215 8553
rect 11241 8527 11242 8553
rect 11046 8526 11242 8527
rect 10878 8023 10879 8049
rect 10905 8023 10906 8049
rect 10878 8017 10906 8023
rect 11046 8049 11074 8526
rect 11214 8521 11242 8526
rect 11270 8442 11298 8447
rect 11270 8395 11298 8414
rect 11214 8330 11242 8335
rect 11214 8329 11410 8330
rect 11214 8303 11215 8329
rect 11241 8303 11410 8329
rect 11214 8302 11410 8303
rect 11214 8297 11242 8302
rect 11046 8023 11047 8049
rect 11073 8023 11074 8049
rect 11046 8017 11074 8023
rect 10318 7961 10346 7966
rect 10654 7994 10682 7999
rect 10654 7947 10682 7966
rect 10766 7965 10794 7971
rect 10766 7939 10767 7965
rect 10793 7939 10794 7965
rect 10206 7239 10207 7265
rect 10233 7239 10234 7265
rect 10206 7233 10234 7239
rect 10654 7602 10682 7607
rect 10766 7602 10794 7939
rect 10654 7601 10794 7602
rect 10654 7575 10655 7601
rect 10681 7575 10794 7601
rect 10654 7574 10794 7575
rect 10878 7938 10906 7943
rect 11382 7938 11410 8302
rect 11438 8218 11466 9478
rect 11494 9473 11522 9478
rect 11606 9338 11634 9343
rect 11494 9226 11522 9231
rect 11494 9179 11522 9198
rect 11606 9225 11634 9310
rect 11662 9282 11690 10066
rect 11718 10066 11746 10071
rect 11774 10066 11802 10375
rect 11746 10038 11802 10066
rect 11718 10019 11746 10038
rect 12782 9674 12810 9679
rect 12614 9618 12642 9623
rect 12614 9571 12642 9590
rect 11942 9561 11970 9567
rect 11942 9535 11943 9561
rect 11969 9535 11970 9561
rect 11662 9249 11690 9254
rect 11774 9505 11802 9511
rect 11886 9506 11914 9511
rect 11774 9479 11775 9505
rect 11801 9479 11802 9505
rect 11606 9199 11607 9225
rect 11633 9199 11634 9225
rect 11606 9193 11634 9199
rect 11774 9225 11802 9479
rect 11774 9199 11775 9225
rect 11801 9199 11802 9225
rect 11774 9193 11802 9199
rect 11830 9505 11914 9506
rect 11830 9479 11887 9505
rect 11913 9479 11914 9505
rect 11830 9478 11914 9479
rect 11830 9226 11858 9478
rect 11886 9473 11914 9478
rect 11942 9394 11970 9535
rect 12782 9561 12810 9646
rect 12782 9535 12783 9561
rect 12809 9535 12810 9561
rect 12782 9529 12810 9535
rect 12110 9506 12138 9511
rect 11942 9366 12082 9394
rect 11998 9282 12026 9287
rect 11998 9235 12026 9254
rect 11830 9193 11858 9198
rect 11886 9170 11914 9175
rect 11886 9169 11970 9170
rect 11886 9143 11887 9169
rect 11913 9143 11970 9169
rect 11886 9142 11970 9143
rect 11886 9137 11914 9142
rect 11942 8889 11970 9142
rect 11998 9114 12026 9119
rect 12054 9114 12082 9366
rect 12110 9225 12138 9478
rect 12110 9199 12111 9225
rect 12137 9199 12138 9225
rect 12110 9193 12138 9199
rect 12950 9226 12978 10431
rect 13734 10094 13762 11551
rect 13846 11578 13874 11583
rect 13846 11531 13874 11550
rect 13958 11577 13986 11583
rect 13958 11551 13959 11577
rect 13985 11551 13986 11577
rect 13958 11186 13986 11551
rect 13958 11153 13986 11158
rect 14014 11577 14042 11583
rect 14014 11551 14015 11577
rect 14041 11551 14042 11577
rect 13174 10066 13202 10071
rect 13118 9674 13146 9679
rect 13118 9627 13146 9646
rect 12950 9193 12978 9198
rect 13006 9562 13034 9567
rect 12026 9086 12082 9114
rect 11998 9081 12026 9086
rect 11942 8863 11943 8889
rect 11969 8863 11970 8889
rect 11942 8857 11970 8863
rect 13006 8889 13034 9534
rect 13062 9506 13090 9511
rect 13062 9459 13090 9478
rect 13006 8863 13007 8889
rect 13033 8863 13034 8889
rect 13006 8857 13034 8863
rect 13118 9226 13146 9231
rect 11606 8834 11634 8839
rect 11606 8787 11634 8806
rect 13118 8834 13146 9198
rect 13174 8889 13202 10038
rect 13566 10066 13594 10071
rect 13566 10019 13594 10038
rect 13678 10066 13762 10094
rect 13790 10794 13818 10799
rect 13398 10009 13426 10015
rect 13398 9983 13399 10009
rect 13425 9983 13426 10009
rect 13174 8863 13175 8889
rect 13201 8863 13202 8889
rect 13174 8857 13202 8863
rect 13230 9674 13258 9679
rect 13118 8553 13146 8806
rect 13230 8778 13258 9646
rect 13398 9618 13426 9983
rect 13678 10009 13706 10066
rect 13790 10065 13818 10766
rect 13790 10039 13791 10065
rect 13817 10039 13818 10065
rect 13790 10033 13818 10039
rect 13902 10738 13930 10743
rect 13902 10065 13930 10710
rect 13902 10039 13903 10065
rect 13929 10039 13930 10065
rect 13902 10033 13930 10039
rect 13958 10066 13986 10071
rect 14014 10066 14042 11551
rect 14294 11241 14322 11247
rect 14294 11215 14295 11241
rect 14321 11215 14322 11241
rect 14294 11186 14322 11215
rect 14294 11153 14322 11158
rect 14630 11241 14658 12838
rect 18942 12698 18970 13511
rect 19950 13482 19978 13847
rect 19950 13449 19978 13454
rect 20006 13593 20034 13599
rect 20006 13567 20007 13593
rect 20033 13567 20034 13593
rect 20006 13146 20034 13567
rect 20006 13113 20034 13118
rect 20006 13033 20034 13039
rect 20006 13007 20007 13033
rect 20033 13007 20034 13033
rect 20006 12810 20034 13007
rect 20006 12777 20034 12782
rect 18942 12665 18970 12670
rect 20118 12417 20146 12423
rect 20118 12391 20119 12417
rect 20145 12391 20146 12417
rect 17598 12166 17730 12171
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17598 12133 17730 12138
rect 20118 12138 20146 12391
rect 20118 12105 20146 12110
rect 17598 11382 17730 11387
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17598 11349 17730 11354
rect 14630 11215 14631 11241
rect 14657 11215 14658 11241
rect 14630 10905 14658 11215
rect 20006 11241 20034 11247
rect 20006 11215 20007 11241
rect 20033 11215 20034 11241
rect 18830 11186 18858 11191
rect 18830 11139 18858 11158
rect 20006 11130 20034 11215
rect 20006 11097 20034 11102
rect 14630 10879 14631 10905
rect 14657 10879 14658 10905
rect 14406 10738 14434 10743
rect 14406 10691 14434 10710
rect 13986 10065 14154 10066
rect 13986 10039 14015 10065
rect 14041 10039 14154 10065
rect 13986 10038 14154 10039
rect 13958 10033 13986 10038
rect 14014 10019 14042 10038
rect 13678 9983 13679 10009
rect 13705 9983 13706 10009
rect 13678 9618 13706 9983
rect 13734 9730 13762 9735
rect 13734 9729 13986 9730
rect 13734 9703 13735 9729
rect 13761 9703 13986 9729
rect 13734 9702 13986 9703
rect 13734 9697 13762 9702
rect 13958 9673 13986 9702
rect 13958 9647 13959 9673
rect 13985 9647 13986 9673
rect 13958 9641 13986 9647
rect 13678 9590 13762 9618
rect 13398 9394 13426 9590
rect 13734 9562 13762 9590
rect 14126 9617 14154 10038
rect 14126 9591 14127 9617
rect 14153 9591 14154 9617
rect 14126 9585 14154 9591
rect 13902 9562 13930 9567
rect 13734 9561 13930 9562
rect 13734 9535 13903 9561
rect 13929 9535 13930 9561
rect 13734 9534 13930 9535
rect 13398 9361 13426 9366
rect 13622 9505 13650 9511
rect 13622 9479 13623 9505
rect 13649 9479 13650 9505
rect 13622 9338 13650 9479
rect 13622 9305 13650 9310
rect 13678 9505 13706 9511
rect 13678 9479 13679 9505
rect 13705 9479 13706 9505
rect 13678 9282 13706 9479
rect 13734 9394 13762 9399
rect 13762 9366 13818 9394
rect 13734 9361 13762 9366
rect 13734 9282 13762 9287
rect 13678 9281 13762 9282
rect 13678 9255 13735 9281
rect 13761 9255 13762 9281
rect 13678 9254 13762 9255
rect 13734 9249 13762 9254
rect 13342 9226 13370 9231
rect 13342 9179 13370 9198
rect 13286 9114 13314 9119
rect 13286 8945 13314 9086
rect 13286 8919 13287 8945
rect 13313 8919 13314 8945
rect 13286 8913 13314 8919
rect 13790 8833 13818 9366
rect 13846 9170 13874 9175
rect 13902 9170 13930 9534
rect 13874 9142 13930 9170
rect 14070 9561 14098 9567
rect 14070 9535 14071 9561
rect 14097 9535 14098 9561
rect 14070 9170 14098 9535
rect 14630 9226 14658 10879
rect 18830 10794 18858 10799
rect 18830 10747 18858 10766
rect 20006 10794 20034 10799
rect 20006 10737 20034 10766
rect 20006 10711 20007 10737
rect 20033 10711 20034 10737
rect 20006 10705 20034 10711
rect 17598 10598 17730 10603
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17598 10565 17730 10570
rect 17598 9814 17730 9819
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17598 9781 17730 9786
rect 20006 9673 20034 9679
rect 20006 9647 20007 9673
rect 20033 9647 20034 9673
rect 18830 9618 18858 9623
rect 18830 9571 18858 9590
rect 20006 9450 20034 9647
rect 20006 9417 20034 9422
rect 14630 9193 14658 9198
rect 15022 9226 15050 9231
rect 18830 9226 18858 9231
rect 15050 9198 15106 9226
rect 15022 9179 15050 9198
rect 13846 9137 13874 9142
rect 14070 9137 14098 9142
rect 14798 9170 14826 9175
rect 14798 9123 14826 9142
rect 14070 9002 14098 9007
rect 14070 8945 14098 8974
rect 14070 8919 14071 8945
rect 14097 8919 14098 8945
rect 14070 8913 14098 8919
rect 13790 8807 13791 8833
rect 13817 8807 13818 8833
rect 13790 8801 13818 8807
rect 14238 8834 14266 8839
rect 14238 8787 14266 8806
rect 14574 8833 14602 8839
rect 14574 8807 14575 8833
rect 14601 8807 14602 8833
rect 13118 8527 13119 8553
rect 13145 8527 13146 8553
rect 13118 8442 13146 8527
rect 11998 8386 12026 8391
rect 11438 8049 11466 8190
rect 11438 8023 11439 8049
rect 11465 8023 11466 8049
rect 11438 8017 11466 8023
rect 11550 8330 11578 8335
rect 11550 8050 11578 8302
rect 11550 8003 11578 8022
rect 11942 8274 11970 8279
rect 11942 8049 11970 8246
rect 11998 8161 12026 8358
rect 11998 8135 11999 8161
rect 12025 8135 12026 8161
rect 11998 8129 12026 8135
rect 11942 8023 11943 8049
rect 11969 8023 11970 8049
rect 11942 8017 11970 8023
rect 11494 7993 11522 7999
rect 11494 7967 11495 7993
rect 11521 7967 11522 7993
rect 11494 7938 11522 7967
rect 11774 7938 11802 7943
rect 11382 7910 11522 7938
rect 11606 7937 11802 7938
rect 11606 7911 11775 7937
rect 11801 7911 11802 7937
rect 11606 7910 11802 7911
rect 9590 7210 9618 7215
rect 9534 7209 9618 7210
rect 9534 7183 9591 7209
rect 9617 7183 9618 7209
rect 9534 7182 9618 7183
rect 9422 7163 9450 7182
rect 9590 7177 9618 7182
rect 10374 7210 10402 7215
rect 10374 7163 10402 7182
rect 9030 6785 9058 6790
rect 9478 7153 9506 7159
rect 9478 7127 9479 7153
rect 9505 7127 9506 7153
rect 8638 6537 8722 6538
rect 8638 6511 8639 6537
rect 8665 6511 8722 6537
rect 8638 6510 8722 6511
rect 8806 6538 8834 6543
rect 8638 6505 8666 6510
rect 8414 4186 8498 4214
rect 2238 3542 2370 3547
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2238 3509 2370 3514
rect 2238 2758 2370 2763
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2238 2725 2370 2730
rect 8078 2618 8106 2623
rect 2238 1974 2370 1979
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2238 1941 2370 1946
rect 8078 400 8106 2590
rect 8190 2561 8218 4186
rect 8190 2535 8191 2561
rect 8217 2535 8218 2561
rect 8190 2529 8218 2535
rect 8470 2170 8498 4186
rect 8694 2618 8722 2623
rect 8694 2571 8722 2590
rect 8694 2170 8722 2175
rect 8470 2169 8722 2170
rect 8470 2143 8695 2169
rect 8721 2143 8722 2169
rect 8470 2142 8722 2143
rect 8694 2137 8722 2142
rect 8414 2058 8442 2063
rect 8414 400 8442 2030
rect 8806 1777 8834 6510
rect 9478 6538 9506 7127
rect 10318 7153 10346 7159
rect 10318 7127 10319 7153
rect 10345 7127 10346 7153
rect 9918 7070 10050 7075
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 9918 7037 10050 7042
rect 10318 6986 10346 7127
rect 10318 6958 10570 6986
rect 10542 6929 10570 6958
rect 10542 6903 10543 6929
rect 10569 6903 10570 6929
rect 10542 6897 10570 6903
rect 10206 6874 10234 6879
rect 10206 6827 10234 6846
rect 9926 6818 9954 6823
rect 9478 6505 9506 6510
rect 9702 6538 9730 6543
rect 9702 6491 9730 6510
rect 9926 6537 9954 6790
rect 9926 6511 9927 6537
rect 9953 6511 9954 6537
rect 9926 6505 9954 6511
rect 9918 6286 10050 6291
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 9918 6253 10050 6258
rect 9918 5502 10050 5507
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 9918 5469 10050 5474
rect 9918 4718 10050 4723
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 9918 4685 10050 4690
rect 10654 4214 10682 7574
rect 10878 7377 10906 7910
rect 11550 7658 11578 7663
rect 11606 7658 11634 7910
rect 11774 7905 11802 7910
rect 11998 7937 12026 7943
rect 11998 7911 11999 7937
rect 12025 7911 12026 7937
rect 11550 7657 11634 7658
rect 11550 7631 11551 7657
rect 11577 7631 11634 7657
rect 11550 7630 11634 7631
rect 11662 7713 11690 7719
rect 11662 7687 11663 7713
rect 11689 7687 11690 7713
rect 11550 7625 11578 7630
rect 11662 7574 11690 7687
rect 11662 7546 11746 7574
rect 10878 7351 10879 7377
rect 10905 7351 10906 7377
rect 10878 7345 10906 7351
rect 11718 7321 11746 7546
rect 11718 7295 11719 7321
rect 11745 7295 11746 7321
rect 11718 7289 11746 7295
rect 11998 7322 12026 7911
rect 11998 7289 12026 7294
rect 12278 7322 12306 7327
rect 11046 7265 11074 7271
rect 11046 7239 11047 7265
rect 11073 7239 11074 7265
rect 10934 7210 10962 7215
rect 10934 7163 10962 7182
rect 11046 6762 11074 7239
rect 11326 7265 11354 7271
rect 11326 7239 11327 7265
rect 11353 7239 11354 7265
rect 11326 6874 11354 7239
rect 11326 6841 11354 6846
rect 11830 6874 11858 6879
rect 11830 6827 11858 6846
rect 11046 6729 11074 6734
rect 11606 6817 11634 6823
rect 11606 6791 11607 6817
rect 11633 6791 11634 6817
rect 11606 6762 11634 6791
rect 11606 6729 11634 6734
rect 11942 6762 11970 6767
rect 10542 4186 10682 4214
rect 9918 3934 10050 3939
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 9918 3901 10050 3906
rect 9918 3150 10050 3155
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 9918 3117 10050 3122
rect 9918 2366 10050 2371
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 9918 2333 10050 2338
rect 10542 2169 10570 4186
rect 10542 2143 10543 2169
rect 10569 2143 10570 2169
rect 10542 2137 10570 2143
rect 9198 2058 9226 2063
rect 9198 2011 9226 2030
rect 10430 2058 10458 2063
rect 8806 1751 8807 1777
rect 8833 1751 8834 1777
rect 8806 1745 8834 1751
rect 9702 1722 9730 1727
rect 9702 1721 9786 1722
rect 9702 1695 9703 1721
rect 9729 1695 9786 1721
rect 9702 1694 9786 1695
rect 9702 1689 9730 1694
rect 9758 400 9786 1694
rect 9918 1582 10050 1587
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 9918 1549 10050 1554
rect 10430 400 10458 2030
rect 11046 2058 11074 2063
rect 11046 2011 11074 2030
rect 11774 1834 11802 1839
rect 11102 1721 11130 1727
rect 11102 1695 11103 1721
rect 11129 1695 11130 1721
rect 11102 400 11130 1695
rect 11774 400 11802 1806
rect 11942 1777 11970 6734
rect 11942 1751 11943 1777
rect 11969 1751 11970 1777
rect 11942 1745 11970 1751
rect 12278 1777 12306 7294
rect 12782 7322 12810 7327
rect 12782 7275 12810 7294
rect 13006 7154 13034 7159
rect 13118 7154 13146 8414
rect 13174 8750 13258 8778
rect 13678 8777 13706 8783
rect 13678 8751 13679 8777
rect 13705 8751 13706 8777
rect 13174 7377 13202 8750
rect 13454 8721 13482 8727
rect 13454 8695 13455 8721
rect 13481 8695 13482 8721
rect 13454 7770 13482 8695
rect 13678 8498 13706 8751
rect 13510 8442 13538 8447
rect 13510 8395 13538 8414
rect 13678 8385 13706 8470
rect 13678 8359 13679 8385
rect 13705 8359 13706 8385
rect 13678 8353 13706 8359
rect 13622 8050 13650 8055
rect 13510 7770 13538 7775
rect 13454 7769 13538 7770
rect 13454 7743 13511 7769
rect 13537 7743 13538 7769
rect 13454 7742 13538 7743
rect 13510 7737 13538 7742
rect 13622 7769 13650 8022
rect 14574 8050 14602 8807
rect 14686 8834 14714 8839
rect 14686 8787 14714 8806
rect 14854 8778 14882 8783
rect 14854 8731 14882 8750
rect 15022 8722 15050 8727
rect 14910 8721 15050 8722
rect 14910 8695 15023 8721
rect 15049 8695 15050 8721
rect 14910 8694 15050 8695
rect 14742 8498 14770 8503
rect 14910 8498 14938 8694
rect 15022 8689 15050 8694
rect 14742 8497 14938 8498
rect 14742 8471 14743 8497
rect 14769 8471 14938 8497
rect 14742 8470 14938 8471
rect 14742 8465 14770 8470
rect 15078 8441 15106 9198
rect 18830 9179 18858 9198
rect 20006 9114 20034 9119
rect 20006 9067 20034 9086
rect 17598 9030 17730 9035
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17598 8997 17730 9002
rect 20006 8889 20034 8895
rect 20006 8863 20007 8889
rect 20033 8863 20034 8889
rect 15134 8833 15162 8839
rect 15134 8807 15135 8833
rect 15161 8807 15162 8833
rect 15134 8778 15162 8807
rect 15134 8745 15162 8750
rect 18830 8833 18858 8839
rect 18830 8807 18831 8833
rect 18857 8807 18858 8833
rect 18830 8498 18858 8807
rect 20006 8778 20034 8863
rect 20006 8745 20034 8750
rect 18830 8465 18858 8470
rect 15078 8415 15079 8441
rect 15105 8415 15106 8441
rect 15078 8409 15106 8415
rect 17598 8246 17730 8251
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17598 8213 17730 8218
rect 14574 8017 14602 8022
rect 13622 7743 13623 7769
rect 13649 7743 13650 7769
rect 13622 7737 13650 7743
rect 13398 7657 13426 7663
rect 18830 7658 18858 7663
rect 13398 7631 13399 7657
rect 13425 7631 13426 7657
rect 13174 7351 13175 7377
rect 13201 7351 13202 7377
rect 13174 7345 13202 7351
rect 13230 7602 13258 7607
rect 13006 7153 13146 7154
rect 13006 7127 13007 7153
rect 13033 7127 13146 7153
rect 13006 7126 13146 7127
rect 12782 6874 12810 6879
rect 13006 6874 13034 7126
rect 13174 6930 13202 6935
rect 13230 6930 13258 7574
rect 13342 7378 13370 7383
rect 13398 7378 13426 7631
rect 18718 7657 18858 7658
rect 18718 7631 18831 7657
rect 18857 7631 18858 7657
rect 18718 7630 18858 7631
rect 13454 7602 13482 7607
rect 13454 7555 13482 7574
rect 17598 7462 17730 7467
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17598 7429 17730 7434
rect 13342 7377 13426 7378
rect 13342 7351 13343 7377
rect 13369 7351 13426 7377
rect 13342 7350 13426 7351
rect 13342 7345 13370 7350
rect 13342 7265 13370 7271
rect 13342 7239 13343 7265
rect 13369 7239 13370 7265
rect 13342 7210 13370 7239
rect 13342 7177 13370 7182
rect 13902 7265 13930 7271
rect 13902 7239 13903 7265
rect 13929 7239 13930 7265
rect 13902 7210 13930 7239
rect 13902 7177 13930 7182
rect 14238 7210 14266 7215
rect 14014 7154 14042 7159
rect 14014 7107 14042 7126
rect 13174 6929 13258 6930
rect 13174 6903 13175 6929
rect 13201 6903 13258 6929
rect 13174 6902 13258 6903
rect 13174 6897 13202 6902
rect 12810 6846 13034 6874
rect 12782 6827 12810 6846
rect 14238 6817 14266 7182
rect 18718 7210 18746 7630
rect 18830 7625 18858 7630
rect 20006 7601 20034 7607
rect 20006 7575 20007 7601
rect 20033 7575 20034 7601
rect 20006 7434 20034 7575
rect 20006 7401 20034 7406
rect 20006 7321 20034 7327
rect 20006 7295 20007 7321
rect 20033 7295 20034 7321
rect 18830 7266 18858 7271
rect 18830 7219 18858 7238
rect 18718 7177 18746 7182
rect 20006 7098 20034 7295
rect 20006 7065 20034 7070
rect 14462 6874 14490 6879
rect 14462 6827 14490 6846
rect 14238 6791 14239 6817
rect 14265 6791 14266 6817
rect 14238 6785 14266 6791
rect 17598 6678 17730 6683
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17598 6645 17730 6650
rect 17598 5894 17730 5899
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17598 5861 17730 5866
rect 17598 5110 17730 5115
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17598 5077 17730 5082
rect 17598 4326 17730 4331
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17598 4293 17730 4298
rect 17598 3542 17730 3547
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17598 3509 17730 3514
rect 17598 2758 17730 2763
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17598 2725 17730 2730
rect 17598 1974 17730 1979
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17598 1941 17730 1946
rect 12782 1834 12810 1839
rect 12782 1787 12810 1806
rect 12278 1751 12279 1777
rect 12305 1751 12306 1777
rect 12278 1745 12306 1751
rect 15246 1666 15274 1671
rect 15134 1665 15274 1666
rect 15134 1639 15247 1665
rect 15273 1639 15274 1665
rect 15134 1638 15274 1639
rect 15134 400 15162 1638
rect 15246 1633 15274 1638
rect 8064 0 8120 400
rect 8400 0 8456 400
rect 9744 0 9800 400
rect 10416 0 10472 400
rect 11088 0 11144 400
rect 11760 0 11816 400
rect 15120 0 15176 400
<< via2 >>
rect 2238 19221 2266 19222
rect 2238 19195 2239 19221
rect 2239 19195 2265 19221
rect 2265 19195 2266 19221
rect 2238 19194 2266 19195
rect 2290 19221 2318 19222
rect 2290 19195 2291 19221
rect 2291 19195 2317 19221
rect 2317 19195 2318 19221
rect 2290 19194 2318 19195
rect 2342 19221 2370 19222
rect 2342 19195 2343 19221
rect 2343 19195 2369 19221
rect 2369 19195 2370 19221
rect 2342 19194 2370 19195
rect 8414 18718 8442 18746
rect 9198 18745 9226 18746
rect 9198 18719 9199 18745
rect 9199 18719 9225 18745
rect 9225 18719 9226 18745
rect 9198 18718 9226 18719
rect 2238 18437 2266 18438
rect 2238 18411 2239 18437
rect 2239 18411 2265 18437
rect 2265 18411 2266 18437
rect 2238 18410 2266 18411
rect 2290 18437 2318 18438
rect 2290 18411 2291 18437
rect 2291 18411 2317 18437
rect 2317 18411 2318 18437
rect 2290 18410 2318 18411
rect 2342 18437 2370 18438
rect 2342 18411 2343 18437
rect 2343 18411 2369 18437
rect 2369 18411 2370 18437
rect 2342 18410 2370 18411
rect 2238 17653 2266 17654
rect 2238 17627 2239 17653
rect 2239 17627 2265 17653
rect 2265 17627 2266 17653
rect 2238 17626 2266 17627
rect 2290 17653 2318 17654
rect 2290 17627 2291 17653
rect 2291 17627 2317 17653
rect 2317 17627 2318 17653
rect 2290 17626 2318 17627
rect 2342 17653 2370 17654
rect 2342 17627 2343 17653
rect 2343 17627 2369 17653
rect 2369 17627 2370 17653
rect 2342 17626 2370 17627
rect 2238 16869 2266 16870
rect 2238 16843 2239 16869
rect 2239 16843 2265 16869
rect 2265 16843 2266 16869
rect 2238 16842 2266 16843
rect 2290 16869 2318 16870
rect 2290 16843 2291 16869
rect 2291 16843 2317 16869
rect 2317 16843 2318 16869
rect 2290 16842 2318 16843
rect 2342 16869 2370 16870
rect 2342 16843 2343 16869
rect 2343 16843 2369 16869
rect 2369 16843 2370 16869
rect 2342 16842 2370 16843
rect 2238 16085 2266 16086
rect 2238 16059 2239 16085
rect 2239 16059 2265 16085
rect 2265 16059 2266 16085
rect 2238 16058 2266 16059
rect 2290 16085 2318 16086
rect 2290 16059 2291 16085
rect 2291 16059 2317 16085
rect 2317 16059 2318 16085
rect 2290 16058 2318 16059
rect 2342 16085 2370 16086
rect 2342 16059 2343 16085
rect 2343 16059 2369 16085
rect 2369 16059 2370 16085
rect 2342 16058 2370 16059
rect 2238 15301 2266 15302
rect 2238 15275 2239 15301
rect 2239 15275 2265 15301
rect 2265 15275 2266 15301
rect 2238 15274 2266 15275
rect 2290 15301 2318 15302
rect 2290 15275 2291 15301
rect 2291 15275 2317 15301
rect 2317 15275 2318 15301
rect 2290 15274 2318 15275
rect 2342 15301 2370 15302
rect 2342 15275 2343 15301
rect 2343 15275 2369 15301
rect 2369 15275 2370 15301
rect 2342 15274 2370 15275
rect 2238 14517 2266 14518
rect 2238 14491 2239 14517
rect 2239 14491 2265 14517
rect 2265 14491 2266 14517
rect 2238 14490 2266 14491
rect 2290 14517 2318 14518
rect 2290 14491 2291 14517
rect 2291 14491 2317 14517
rect 2317 14491 2318 14517
rect 2290 14490 2318 14491
rect 2342 14517 2370 14518
rect 2342 14491 2343 14517
rect 2343 14491 2369 14517
rect 2369 14491 2370 14517
rect 2342 14490 2370 14491
rect 2238 13733 2266 13734
rect 2238 13707 2239 13733
rect 2239 13707 2265 13733
rect 2265 13707 2266 13733
rect 2238 13706 2266 13707
rect 2290 13733 2318 13734
rect 2290 13707 2291 13733
rect 2291 13707 2317 13733
rect 2317 13707 2318 13733
rect 2290 13706 2318 13707
rect 2342 13733 2370 13734
rect 2342 13707 2343 13733
rect 2343 13707 2369 13733
rect 2369 13707 2370 13733
rect 2342 13706 2370 13707
rect 2086 13454 2114 13482
rect 966 10094 994 10122
rect 2238 12949 2266 12950
rect 2238 12923 2239 12949
rect 2239 12923 2265 12949
rect 2265 12923 2266 12949
rect 2238 12922 2266 12923
rect 2290 12949 2318 12950
rect 2290 12923 2291 12949
rect 2291 12923 2317 12949
rect 2317 12923 2318 12949
rect 2290 12922 2318 12923
rect 2342 12949 2370 12950
rect 2342 12923 2343 12949
rect 2343 12923 2369 12949
rect 2369 12923 2370 12949
rect 2342 12922 2370 12923
rect 8078 13454 8106 13482
rect 8694 13481 8722 13482
rect 8694 13455 8695 13481
rect 8695 13455 8721 13481
rect 8721 13455 8722 13481
rect 8694 13454 8722 13455
rect 8862 13230 8890 13258
rect 7518 13118 7546 13146
rect 7182 12726 7210 12754
rect 7518 12726 7546 12754
rect 2238 12165 2266 12166
rect 2238 12139 2239 12165
rect 2239 12139 2265 12165
rect 2265 12139 2266 12165
rect 2238 12138 2266 12139
rect 2290 12165 2318 12166
rect 2290 12139 2291 12165
rect 2291 12139 2317 12165
rect 2317 12139 2318 12165
rect 2290 12138 2318 12139
rect 2342 12165 2370 12166
rect 2342 12139 2343 12165
rect 2343 12139 2369 12165
rect 2369 12139 2370 12165
rect 2342 12138 2370 12139
rect 5894 12054 5922 12082
rect 6566 12361 6594 12362
rect 6566 12335 6567 12361
rect 6567 12335 6593 12361
rect 6593 12335 6594 12361
rect 6566 12334 6594 12335
rect 2238 11381 2266 11382
rect 2238 11355 2239 11381
rect 2239 11355 2265 11381
rect 2265 11355 2266 11381
rect 2238 11354 2266 11355
rect 2290 11381 2318 11382
rect 2290 11355 2291 11381
rect 2291 11355 2317 11381
rect 2317 11355 2318 11381
rect 2290 11354 2318 11355
rect 2342 11381 2370 11382
rect 2342 11355 2343 11381
rect 2343 11355 2369 11381
rect 2369 11355 2370 11381
rect 2342 11354 2370 11355
rect 7798 12753 7826 12754
rect 7798 12727 7799 12753
rect 7799 12727 7825 12753
rect 7825 12727 7826 12753
rect 7798 12726 7826 12727
rect 7966 12334 7994 12362
rect 7462 11185 7490 11186
rect 7462 11159 7463 11185
rect 7463 11159 7489 11185
rect 7489 11159 7490 11185
rect 7462 11158 7490 11159
rect 7182 11102 7210 11130
rect 5838 10878 5866 10906
rect 2238 10597 2266 10598
rect 2238 10571 2239 10597
rect 2239 10571 2265 10597
rect 2265 10571 2266 10597
rect 2238 10570 2266 10571
rect 2290 10597 2318 10598
rect 2290 10571 2291 10597
rect 2291 10571 2317 10597
rect 2317 10571 2318 10597
rect 2290 10570 2318 10571
rect 2342 10597 2370 10598
rect 2342 10571 2343 10597
rect 2343 10571 2369 10597
rect 2369 10571 2370 10597
rect 2342 10570 2370 10571
rect 2142 10401 2170 10402
rect 2142 10375 2143 10401
rect 2143 10375 2169 10401
rect 2169 10375 2170 10401
rect 2142 10374 2170 10375
rect 5334 10374 5362 10402
rect 2086 9926 2114 9954
rect 2238 9813 2266 9814
rect 2238 9787 2239 9813
rect 2239 9787 2265 9813
rect 2265 9787 2266 9813
rect 2238 9786 2266 9787
rect 2290 9813 2318 9814
rect 2290 9787 2291 9813
rect 2291 9787 2317 9813
rect 2317 9787 2318 9813
rect 2290 9786 2318 9787
rect 2342 9813 2370 9814
rect 2342 9787 2343 9813
rect 2343 9787 2369 9813
rect 2369 9787 2370 9813
rect 5334 9814 5362 9842
rect 2342 9786 2370 9787
rect 8190 13145 8218 13146
rect 8190 13119 8191 13145
rect 8191 13119 8217 13145
rect 8217 13119 8218 13145
rect 8190 13118 8218 13119
rect 8414 12726 8442 12754
rect 8190 12502 8218 12530
rect 8414 12473 8442 12474
rect 8414 12447 8415 12473
rect 8415 12447 8441 12473
rect 8441 12447 8442 12473
rect 8414 12446 8442 12447
rect 8750 12502 8778 12530
rect 9918 18829 9946 18830
rect 9918 18803 9919 18829
rect 9919 18803 9945 18829
rect 9945 18803 9946 18829
rect 9918 18802 9946 18803
rect 9970 18829 9998 18830
rect 9970 18803 9971 18829
rect 9971 18803 9997 18829
rect 9997 18803 9998 18829
rect 9970 18802 9998 18803
rect 10022 18829 10050 18830
rect 10022 18803 10023 18829
rect 10023 18803 10049 18829
rect 10049 18803 10050 18829
rect 10022 18802 10050 18803
rect 17598 19221 17626 19222
rect 17598 19195 17599 19221
rect 17599 19195 17625 19221
rect 17625 19195 17626 19221
rect 17598 19194 17626 19195
rect 17650 19221 17678 19222
rect 17650 19195 17651 19221
rect 17651 19195 17677 19221
rect 17677 19195 17678 19221
rect 17650 19194 17678 19195
rect 17702 19221 17730 19222
rect 17702 19195 17703 19221
rect 17703 19195 17729 19221
rect 17729 19195 17730 19221
rect 17702 19194 17730 19195
rect 10766 18718 10794 18746
rect 11382 18745 11410 18746
rect 11382 18719 11383 18745
rect 11383 18719 11409 18745
rect 11409 18719 11410 18745
rect 11382 18718 11410 18719
rect 9918 18045 9946 18046
rect 9918 18019 9919 18045
rect 9919 18019 9945 18045
rect 9945 18019 9946 18045
rect 9918 18018 9946 18019
rect 9970 18045 9998 18046
rect 9970 18019 9971 18045
rect 9971 18019 9997 18045
rect 9997 18019 9998 18045
rect 9970 18018 9998 18019
rect 10022 18045 10050 18046
rect 10022 18019 10023 18045
rect 10023 18019 10049 18045
rect 10049 18019 10050 18045
rect 10022 18018 10050 18019
rect 9918 17261 9946 17262
rect 9918 17235 9919 17261
rect 9919 17235 9945 17261
rect 9945 17235 9946 17261
rect 9918 17234 9946 17235
rect 9970 17261 9998 17262
rect 9970 17235 9971 17261
rect 9971 17235 9997 17261
rect 9997 17235 9998 17261
rect 9970 17234 9998 17235
rect 10022 17261 10050 17262
rect 10022 17235 10023 17261
rect 10023 17235 10049 17261
rect 10049 17235 10050 17261
rect 10022 17234 10050 17235
rect 9918 16477 9946 16478
rect 9918 16451 9919 16477
rect 9919 16451 9945 16477
rect 9945 16451 9946 16477
rect 9918 16450 9946 16451
rect 9970 16477 9998 16478
rect 9970 16451 9971 16477
rect 9971 16451 9997 16477
rect 9997 16451 9998 16477
rect 9970 16450 9998 16451
rect 10022 16477 10050 16478
rect 10022 16451 10023 16477
rect 10023 16451 10049 16477
rect 10049 16451 10050 16477
rect 10022 16450 10050 16451
rect 9918 15693 9946 15694
rect 9918 15667 9919 15693
rect 9919 15667 9945 15693
rect 9945 15667 9946 15693
rect 9918 15666 9946 15667
rect 9970 15693 9998 15694
rect 9970 15667 9971 15693
rect 9971 15667 9997 15693
rect 9997 15667 9998 15693
rect 9970 15666 9998 15667
rect 10022 15693 10050 15694
rect 10022 15667 10023 15693
rect 10023 15667 10049 15693
rect 10049 15667 10050 15693
rect 10022 15666 10050 15667
rect 9918 14909 9946 14910
rect 9918 14883 9919 14909
rect 9919 14883 9945 14909
rect 9945 14883 9946 14909
rect 9918 14882 9946 14883
rect 9970 14909 9998 14910
rect 9970 14883 9971 14909
rect 9971 14883 9997 14909
rect 9997 14883 9998 14909
rect 9970 14882 9998 14883
rect 10022 14909 10050 14910
rect 10022 14883 10023 14909
rect 10023 14883 10049 14909
rect 10049 14883 10050 14909
rect 10022 14882 10050 14883
rect 9918 14125 9946 14126
rect 9918 14099 9919 14125
rect 9919 14099 9945 14125
rect 9945 14099 9946 14125
rect 9918 14098 9946 14099
rect 9970 14125 9998 14126
rect 9970 14099 9971 14125
rect 9971 14099 9997 14125
rect 9997 14099 9998 14125
rect 9970 14098 9998 14099
rect 10022 14125 10050 14126
rect 10022 14099 10023 14125
rect 10023 14099 10049 14125
rect 10049 14099 10050 14125
rect 10022 14098 10050 14099
rect 9918 13341 9946 13342
rect 9918 13315 9919 13341
rect 9919 13315 9945 13341
rect 9945 13315 9946 13341
rect 9918 13314 9946 13315
rect 9970 13341 9998 13342
rect 9970 13315 9971 13341
rect 9971 13315 9997 13341
rect 9997 13315 9998 13341
rect 9970 13314 9998 13315
rect 10022 13341 10050 13342
rect 10022 13315 10023 13341
rect 10023 13315 10049 13341
rect 10049 13315 10050 13341
rect 10022 13314 10050 13315
rect 9310 13257 9338 13258
rect 9310 13231 9311 13257
rect 9311 13231 9337 13257
rect 9337 13231 9338 13257
rect 9310 13230 9338 13231
rect 9870 13145 9898 13146
rect 9870 13119 9871 13145
rect 9871 13119 9897 13145
rect 9897 13119 9898 13145
rect 9870 13118 9898 13119
rect 9534 12753 9562 12754
rect 9534 12727 9535 12753
rect 9535 12727 9561 12753
rect 9561 12727 9562 12753
rect 9534 12726 9562 12727
rect 10262 12726 10290 12754
rect 9086 12446 9114 12474
rect 9422 12473 9450 12474
rect 9422 12447 9423 12473
rect 9423 12447 9449 12473
rect 9449 12447 9450 12473
rect 9422 12446 9450 12447
rect 10094 12614 10122 12642
rect 9918 12557 9946 12558
rect 9918 12531 9919 12557
rect 9919 12531 9945 12557
rect 9945 12531 9946 12557
rect 9918 12530 9946 12531
rect 9970 12557 9998 12558
rect 9970 12531 9971 12557
rect 9971 12531 9997 12557
rect 9997 12531 9998 12557
rect 9970 12530 9998 12531
rect 10022 12557 10050 12558
rect 10022 12531 10023 12557
rect 10023 12531 10049 12557
rect 10049 12531 10050 12557
rect 10022 12530 10050 12531
rect 9646 12446 9674 12474
rect 8078 12222 8106 12250
rect 7966 11718 7994 11746
rect 7742 11494 7770 11522
rect 7406 10905 7434 10906
rect 7406 10879 7407 10905
rect 7407 10879 7433 10905
rect 7433 10879 7434 10905
rect 7406 10878 7434 10879
rect 7350 10822 7378 10850
rect 7854 11185 7882 11186
rect 7854 11159 7855 11185
rect 7855 11159 7881 11185
rect 7881 11159 7882 11185
rect 7854 11158 7882 11159
rect 9142 12361 9170 12362
rect 9142 12335 9143 12361
rect 9143 12335 9169 12361
rect 9169 12335 9170 12361
rect 9142 12334 9170 12335
rect 8806 12305 8834 12306
rect 8806 12279 8807 12305
rect 8807 12279 8833 12305
rect 8833 12279 8834 12305
rect 8806 12278 8834 12279
rect 8918 12249 8946 12250
rect 8918 12223 8919 12249
rect 8919 12223 8945 12249
rect 8945 12223 8946 12249
rect 8918 12222 8946 12223
rect 8246 11718 8274 11746
rect 8694 11718 8722 11746
rect 8078 11633 8106 11634
rect 8078 11607 8079 11633
rect 8079 11607 8105 11633
rect 8105 11607 8106 11633
rect 8078 11606 8106 11607
rect 8078 11494 8106 11522
rect 8022 11214 8050 11242
rect 8078 11185 8106 11186
rect 8078 11159 8079 11185
rect 8079 11159 8105 11185
rect 8105 11159 8106 11185
rect 8078 11158 8106 11159
rect 8134 11102 8162 11130
rect 8750 11606 8778 11634
rect 8414 11185 8442 11186
rect 8414 11159 8415 11185
rect 8415 11159 8441 11185
rect 8441 11159 8442 11185
rect 8414 11158 8442 11159
rect 8750 11185 8778 11186
rect 8750 11159 8751 11185
rect 8751 11159 8777 11185
rect 8777 11159 8778 11185
rect 8750 11158 8778 11159
rect 8358 11102 8386 11130
rect 8246 10934 8274 10962
rect 7742 10822 7770 10850
rect 8022 10457 8050 10458
rect 8022 10431 8023 10457
rect 8023 10431 8049 10457
rect 8049 10431 8050 10457
rect 8022 10430 8050 10431
rect 6118 9758 6146 9786
rect 7014 9982 7042 10010
rect 6734 9758 6762 9786
rect 6230 9673 6258 9674
rect 6230 9647 6231 9673
rect 6231 9647 6257 9673
rect 6257 9647 6258 9673
rect 6230 9646 6258 9647
rect 2142 9225 2170 9226
rect 2142 9199 2143 9225
rect 2143 9199 2169 9225
rect 2169 9199 2170 9225
rect 2142 9198 2170 9199
rect 6230 9225 6258 9226
rect 6230 9199 6231 9225
rect 6231 9199 6257 9225
rect 6257 9199 6258 9225
rect 6230 9198 6258 9199
rect 5166 9169 5194 9170
rect 5166 9143 5167 9169
rect 5167 9143 5193 9169
rect 5193 9143 5194 9169
rect 5166 9142 5194 9143
rect 966 9113 994 9114
rect 966 9087 967 9113
rect 967 9087 993 9113
rect 993 9087 994 9113
rect 966 9086 994 9087
rect 2238 9029 2266 9030
rect 2238 9003 2239 9029
rect 2239 9003 2265 9029
rect 2265 9003 2266 9029
rect 2238 9002 2266 9003
rect 2290 9029 2318 9030
rect 2290 9003 2291 9029
rect 2291 9003 2317 9029
rect 2317 9003 2318 9029
rect 2290 9002 2318 9003
rect 2342 9029 2370 9030
rect 2342 9003 2343 9029
rect 2343 9003 2369 9029
rect 2369 9003 2370 9029
rect 2342 9002 2370 9003
rect 6622 9142 6650 9170
rect 5166 8750 5194 8778
rect 6902 9254 6930 9282
rect 6846 9225 6874 9226
rect 6846 9199 6847 9225
rect 6847 9199 6873 9225
rect 6873 9199 6874 9225
rect 6846 9198 6874 9199
rect 6958 9366 6986 9394
rect 6790 8777 6818 8778
rect 6790 8751 6791 8777
rect 6791 8751 6817 8777
rect 6817 8751 6818 8777
rect 6790 8750 6818 8751
rect 7182 9646 7210 9674
rect 7910 10065 7938 10066
rect 7910 10039 7911 10065
rect 7911 10039 7937 10065
rect 7937 10039 7938 10065
rect 7910 10038 7938 10039
rect 7406 9982 7434 10010
rect 7686 9897 7714 9898
rect 7686 9871 7687 9897
rect 7687 9871 7713 9897
rect 7713 9871 7714 9897
rect 7686 9870 7714 9871
rect 7630 9646 7658 9674
rect 7574 9617 7602 9618
rect 7574 9591 7575 9617
rect 7575 9591 7601 9617
rect 7601 9591 7602 9617
rect 7574 9590 7602 9591
rect 7182 9366 7210 9394
rect 7966 9590 7994 9618
rect 7966 9478 7994 9506
rect 8526 10766 8554 10794
rect 9086 11689 9114 11690
rect 9086 11663 9087 11689
rect 9087 11663 9113 11689
rect 9113 11663 9114 11689
rect 9086 11662 9114 11663
rect 8974 11270 9002 11298
rect 9086 11158 9114 11186
rect 8862 10878 8890 10906
rect 8694 10094 8722 10122
rect 8358 10065 8386 10066
rect 8358 10039 8359 10065
rect 8359 10039 8385 10065
rect 8385 10039 8386 10065
rect 8358 10038 8386 10039
rect 8862 10793 8890 10794
rect 8862 10767 8863 10793
rect 8863 10767 8889 10793
rect 8889 10767 8890 10793
rect 8862 10766 8890 10767
rect 9198 11185 9226 11186
rect 9198 11159 9199 11185
rect 9199 11159 9225 11185
rect 9225 11159 9226 11185
rect 9198 11158 9226 11159
rect 9142 11129 9170 11130
rect 9142 11103 9143 11129
rect 9143 11103 9169 11129
rect 9169 11103 9170 11129
rect 9142 11102 9170 11103
rect 9918 11773 9946 11774
rect 9918 11747 9919 11773
rect 9919 11747 9945 11773
rect 9945 11747 9946 11773
rect 9918 11746 9946 11747
rect 9970 11773 9998 11774
rect 9970 11747 9971 11773
rect 9971 11747 9997 11773
rect 9997 11747 9998 11773
rect 9970 11746 9998 11747
rect 10022 11773 10050 11774
rect 10022 11747 10023 11773
rect 10023 11747 10049 11773
rect 10049 11747 10050 11773
rect 10022 11746 10050 11747
rect 10150 11774 10178 11802
rect 10094 11185 10122 11186
rect 10094 11159 10095 11185
rect 10095 11159 10121 11185
rect 10121 11159 10122 11185
rect 10094 11158 10122 11159
rect 9478 10934 9506 10962
rect 9310 10849 9338 10850
rect 9310 10823 9311 10849
rect 9311 10823 9337 10849
rect 9337 10823 9338 10849
rect 9310 10822 9338 10823
rect 8918 10094 8946 10122
rect 8862 10065 8890 10066
rect 8862 10039 8863 10065
rect 8863 10039 8889 10065
rect 8889 10039 8890 10065
rect 8862 10038 8890 10039
rect 8358 9337 8386 9338
rect 8358 9311 8359 9337
rect 8359 9311 8385 9337
rect 8385 9311 8386 9337
rect 8358 9310 8386 9311
rect 7014 9142 7042 9170
rect 7798 9225 7826 9226
rect 7798 9199 7799 9225
rect 7799 9199 7825 9225
rect 7825 9199 7826 9225
rect 7798 9198 7826 9199
rect 6734 8526 6762 8554
rect 6566 8470 6594 8498
rect 2142 8441 2170 8442
rect 2142 8415 2143 8441
rect 2143 8415 2169 8441
rect 2169 8415 2170 8441
rect 2142 8414 2170 8415
rect 5502 8414 5530 8442
rect 2238 8245 2266 8246
rect 2238 8219 2239 8245
rect 2239 8219 2265 8245
rect 2265 8219 2266 8245
rect 2238 8218 2266 8219
rect 2290 8245 2318 8246
rect 2290 8219 2291 8245
rect 2291 8219 2317 8245
rect 2317 8219 2318 8245
rect 2290 8218 2318 8219
rect 2342 8245 2370 8246
rect 2342 8219 2343 8245
rect 2343 8219 2369 8245
rect 2369 8219 2370 8245
rect 2342 8218 2370 8219
rect 966 8078 994 8106
rect 7014 8553 7042 8554
rect 7014 8527 7015 8553
rect 7015 8527 7041 8553
rect 7041 8527 7042 8553
rect 7014 8526 7042 8527
rect 7238 9142 7266 9170
rect 7126 8526 7154 8554
rect 6958 8441 6986 8442
rect 6958 8415 6959 8441
rect 6959 8415 6985 8441
rect 6985 8415 6986 8441
rect 6958 8414 6986 8415
rect 6902 8358 6930 8386
rect 6846 8190 6874 8218
rect 7126 8105 7154 8106
rect 7126 8079 7127 8105
rect 7127 8079 7153 8105
rect 7153 8079 7154 8105
rect 7126 8078 7154 8079
rect 8414 9142 8442 9170
rect 8358 8974 8386 9002
rect 8302 8777 8330 8778
rect 8302 8751 8303 8777
rect 8303 8751 8329 8777
rect 8329 8751 8330 8777
rect 8302 8750 8330 8751
rect 7350 8694 7378 8722
rect 8246 8721 8274 8722
rect 8246 8695 8247 8721
rect 8247 8695 8273 8721
rect 8273 8695 8274 8721
rect 8246 8694 8274 8695
rect 7854 8638 7882 8666
rect 7686 8582 7714 8610
rect 7462 8497 7490 8498
rect 7462 8471 7463 8497
rect 7463 8471 7489 8497
rect 7489 8471 7490 8497
rect 7462 8470 7490 8471
rect 7294 8441 7322 8442
rect 7294 8415 7295 8441
rect 7295 8415 7321 8441
rect 7321 8415 7322 8441
rect 7294 8414 7322 8415
rect 7742 8553 7770 8554
rect 7742 8527 7743 8553
rect 7743 8527 7769 8553
rect 7769 8527 7770 8553
rect 7742 8526 7770 8527
rect 7294 7518 7322 7546
rect 2238 7461 2266 7462
rect 2238 7435 2239 7461
rect 2239 7435 2265 7461
rect 2265 7435 2266 7461
rect 2238 7434 2266 7435
rect 2290 7461 2318 7462
rect 2290 7435 2291 7461
rect 2291 7435 2317 7461
rect 2317 7435 2318 7461
rect 2290 7434 2318 7435
rect 2342 7461 2370 7462
rect 2342 7435 2343 7461
rect 2343 7435 2369 7461
rect 2369 7435 2370 7461
rect 2342 7434 2370 7435
rect 7798 8078 7826 8106
rect 8414 8721 8442 8722
rect 8414 8695 8415 8721
rect 8415 8695 8441 8721
rect 8441 8695 8442 8721
rect 8414 8694 8442 8695
rect 8078 7377 8106 7378
rect 8078 7351 8079 7377
rect 8079 7351 8105 7377
rect 8105 7351 8106 7377
rect 8078 7350 8106 7351
rect 8190 7265 8218 7266
rect 8190 7239 8191 7265
rect 8191 7239 8217 7265
rect 8217 7239 8218 7265
rect 8190 7238 8218 7239
rect 7350 7182 7378 7210
rect 7910 7209 7938 7210
rect 7910 7183 7911 7209
rect 7911 7183 7937 7209
rect 7937 7183 7938 7209
rect 7910 7182 7938 7183
rect 2238 6677 2266 6678
rect 2238 6651 2239 6677
rect 2239 6651 2265 6677
rect 2265 6651 2266 6677
rect 2238 6650 2266 6651
rect 2290 6677 2318 6678
rect 2290 6651 2291 6677
rect 2291 6651 2317 6677
rect 2317 6651 2318 6677
rect 2290 6650 2318 6651
rect 2342 6677 2370 6678
rect 2342 6651 2343 6677
rect 2343 6651 2369 6677
rect 2369 6651 2370 6677
rect 2342 6650 2370 6651
rect 2238 5893 2266 5894
rect 2238 5867 2239 5893
rect 2239 5867 2265 5893
rect 2265 5867 2266 5893
rect 2238 5866 2266 5867
rect 2290 5893 2318 5894
rect 2290 5867 2291 5893
rect 2291 5867 2317 5893
rect 2317 5867 2318 5893
rect 2290 5866 2318 5867
rect 2342 5893 2370 5894
rect 2342 5867 2343 5893
rect 2343 5867 2369 5893
rect 2369 5867 2370 5893
rect 2342 5866 2370 5867
rect 2238 5109 2266 5110
rect 2238 5083 2239 5109
rect 2239 5083 2265 5109
rect 2265 5083 2266 5109
rect 2238 5082 2266 5083
rect 2290 5109 2318 5110
rect 2290 5083 2291 5109
rect 2291 5083 2317 5109
rect 2317 5083 2318 5109
rect 2290 5082 2318 5083
rect 2342 5109 2370 5110
rect 2342 5083 2343 5109
rect 2343 5083 2369 5109
rect 2369 5083 2370 5109
rect 2342 5082 2370 5083
rect 2238 4325 2266 4326
rect 2238 4299 2239 4325
rect 2239 4299 2265 4325
rect 2265 4299 2266 4325
rect 2238 4298 2266 4299
rect 2290 4325 2318 4326
rect 2290 4299 2291 4325
rect 2291 4299 2317 4325
rect 2317 4299 2318 4325
rect 2290 4298 2318 4299
rect 2342 4325 2370 4326
rect 2342 4299 2343 4325
rect 2343 4299 2369 4325
rect 2369 4299 2370 4325
rect 2342 4298 2370 4299
rect 8694 9310 8722 9338
rect 8638 9254 8666 9282
rect 8582 8974 8610 9002
rect 8358 7518 8386 7546
rect 9310 10513 9338 10514
rect 9310 10487 9311 10513
rect 9311 10487 9337 10513
rect 9337 10487 9338 10513
rect 9310 10486 9338 10487
rect 9142 10038 9170 10066
rect 9030 10009 9058 10010
rect 9030 9983 9031 10009
rect 9031 9983 9057 10009
rect 9057 9983 9058 10009
rect 9030 9982 9058 9983
rect 9918 10989 9946 10990
rect 9590 10934 9618 10962
rect 9918 10963 9919 10989
rect 9919 10963 9945 10989
rect 9945 10963 9946 10989
rect 9918 10962 9946 10963
rect 9970 10989 9998 10990
rect 9970 10963 9971 10989
rect 9971 10963 9997 10989
rect 9997 10963 9998 10989
rect 9970 10962 9998 10963
rect 10022 10989 10050 10990
rect 10022 10963 10023 10989
rect 10023 10963 10049 10989
rect 10049 10963 10050 10989
rect 10022 10962 10050 10963
rect 9030 9478 9058 9506
rect 9366 9982 9394 10010
rect 9254 9478 9282 9506
rect 8974 9310 9002 9338
rect 8974 9142 9002 9170
rect 9198 9337 9226 9338
rect 9198 9311 9199 9337
rect 9199 9311 9225 9337
rect 9225 9311 9226 9337
rect 9198 9310 9226 9311
rect 8918 8694 8946 8722
rect 9142 8582 9170 8610
rect 9366 8777 9394 8778
rect 9366 8751 9367 8777
rect 9367 8751 9393 8777
rect 9393 8751 9394 8777
rect 9366 8750 9394 8751
rect 9086 8526 9114 8554
rect 8750 7350 8778 7378
rect 8526 7321 8554 7322
rect 8526 7295 8527 7321
rect 8527 7295 8553 7321
rect 8553 7295 8554 7321
rect 8526 7294 8554 7295
rect 8414 7238 8442 7266
rect 8302 6790 8330 6818
rect 8862 7209 8890 7210
rect 8862 7183 8863 7209
rect 8863 7183 8889 7209
rect 8889 7183 8890 7209
rect 8862 7182 8890 7183
rect 8750 6817 8778 6818
rect 8750 6791 8751 6817
rect 8751 6791 8777 6817
rect 8777 6791 8778 6817
rect 8750 6790 8778 6791
rect 9534 9953 9562 9954
rect 9534 9927 9535 9953
rect 9535 9927 9561 9953
rect 9561 9927 9562 9953
rect 9534 9926 9562 9927
rect 9590 9337 9618 9338
rect 9590 9311 9591 9337
rect 9591 9311 9617 9337
rect 9617 9311 9618 9337
rect 9590 9310 9618 9311
rect 9918 10205 9946 10206
rect 9918 10179 9919 10205
rect 9919 10179 9945 10205
rect 9945 10179 9946 10205
rect 9918 10178 9946 10179
rect 9970 10205 9998 10206
rect 9970 10179 9971 10205
rect 9971 10179 9997 10205
rect 9997 10179 9998 10205
rect 9970 10178 9998 10179
rect 10022 10205 10050 10206
rect 10022 10179 10023 10205
rect 10023 10179 10049 10205
rect 10049 10179 10050 10205
rect 10022 10178 10050 10179
rect 10038 10038 10066 10066
rect 9918 9421 9946 9422
rect 9918 9395 9919 9421
rect 9919 9395 9945 9421
rect 9945 9395 9946 9421
rect 9918 9394 9946 9395
rect 9970 9421 9998 9422
rect 9970 9395 9971 9421
rect 9971 9395 9997 9421
rect 9997 9395 9998 9421
rect 9970 9394 9998 9395
rect 10022 9421 10050 9422
rect 10022 9395 10023 9421
rect 10023 9395 10049 9421
rect 10049 9395 10050 9421
rect 10022 9394 10050 9395
rect 9814 9310 9842 9338
rect 10318 12697 10346 12698
rect 10318 12671 10319 12697
rect 10319 12671 10345 12697
rect 10345 12671 10346 12697
rect 10318 12670 10346 12671
rect 10766 12278 10794 12306
rect 10654 12081 10682 12082
rect 10654 12055 10655 12081
rect 10655 12055 10681 12081
rect 10681 12055 10682 12081
rect 10654 12054 10682 12055
rect 10318 11297 10346 11298
rect 10318 11271 10319 11297
rect 10319 11271 10345 11297
rect 10345 11271 10346 11297
rect 10318 11270 10346 11271
rect 10318 11185 10346 11186
rect 10318 11159 10319 11185
rect 10319 11159 10345 11185
rect 10345 11159 10346 11185
rect 10318 11158 10346 11159
rect 10206 10486 10234 10514
rect 17598 18437 17626 18438
rect 17598 18411 17599 18437
rect 17599 18411 17625 18437
rect 17625 18411 17626 18437
rect 17598 18410 17626 18411
rect 17650 18437 17678 18438
rect 17650 18411 17651 18437
rect 17651 18411 17677 18437
rect 17677 18411 17678 18437
rect 17650 18410 17678 18411
rect 17702 18437 17730 18438
rect 17702 18411 17703 18437
rect 17703 18411 17729 18437
rect 17729 18411 17730 18437
rect 17702 18410 17730 18411
rect 17598 17653 17626 17654
rect 17598 17627 17599 17653
rect 17599 17627 17625 17653
rect 17625 17627 17626 17653
rect 17598 17626 17626 17627
rect 17650 17653 17678 17654
rect 17650 17627 17651 17653
rect 17651 17627 17677 17653
rect 17677 17627 17678 17653
rect 17650 17626 17678 17627
rect 17702 17653 17730 17654
rect 17702 17627 17703 17653
rect 17703 17627 17729 17653
rect 17729 17627 17730 17653
rect 17702 17626 17730 17627
rect 17598 16869 17626 16870
rect 17598 16843 17599 16869
rect 17599 16843 17625 16869
rect 17625 16843 17626 16869
rect 17598 16842 17626 16843
rect 17650 16869 17678 16870
rect 17650 16843 17651 16869
rect 17651 16843 17677 16869
rect 17677 16843 17678 16869
rect 17650 16842 17678 16843
rect 17702 16869 17730 16870
rect 17702 16843 17703 16869
rect 17703 16843 17729 16869
rect 17729 16843 17730 16869
rect 17702 16842 17730 16843
rect 17598 16085 17626 16086
rect 17598 16059 17599 16085
rect 17599 16059 17625 16085
rect 17625 16059 17626 16085
rect 17598 16058 17626 16059
rect 17650 16085 17678 16086
rect 17650 16059 17651 16085
rect 17651 16059 17677 16085
rect 17677 16059 17678 16085
rect 17650 16058 17678 16059
rect 17702 16085 17730 16086
rect 17702 16059 17703 16085
rect 17703 16059 17729 16085
rect 17729 16059 17730 16085
rect 17702 16058 17730 16059
rect 12614 13481 12642 13482
rect 12614 13455 12615 13481
rect 12615 13455 12641 13481
rect 12641 13455 12642 13481
rect 12614 13454 12642 13455
rect 11550 13230 11578 13258
rect 12334 13230 12362 13258
rect 12278 13201 12306 13202
rect 12278 13175 12279 13201
rect 12279 13175 12305 13201
rect 12305 13175 12306 13201
rect 12278 13174 12306 13175
rect 11606 13118 11634 13146
rect 11830 13145 11858 13146
rect 11830 13119 11831 13145
rect 11831 13119 11857 13145
rect 11857 13119 11858 13145
rect 11830 13118 11858 13119
rect 11046 12670 11074 12698
rect 10878 12641 10906 12642
rect 10878 12615 10879 12641
rect 10879 12615 10905 12641
rect 10905 12615 10906 12641
rect 10878 12614 10906 12615
rect 10934 12558 10962 12586
rect 11550 12558 11578 12586
rect 10822 11969 10850 11970
rect 10822 11943 10823 11969
rect 10823 11943 10849 11969
rect 10849 11943 10850 11969
rect 10822 11942 10850 11943
rect 10934 11774 10962 11802
rect 11494 11942 11522 11970
rect 10654 11185 10682 11186
rect 10654 11159 10655 11185
rect 10655 11159 10681 11185
rect 10681 11159 10682 11185
rect 10654 11158 10682 11159
rect 10542 11102 10570 11130
rect 10318 10206 10346 10234
rect 10262 9982 10290 10010
rect 9982 9337 10010 9338
rect 9982 9311 9983 9337
rect 9983 9311 10009 9337
rect 10009 9311 10010 9337
rect 9982 9310 10010 9311
rect 10206 9646 10234 9674
rect 9926 9281 9954 9282
rect 9926 9255 9927 9281
rect 9927 9255 9953 9281
rect 9953 9255 9954 9281
rect 9926 9254 9954 9255
rect 9982 9113 10010 9114
rect 9982 9087 9983 9113
rect 9983 9087 10009 9113
rect 10009 9087 10010 9113
rect 9982 9086 10010 9087
rect 9758 9030 9786 9058
rect 9534 8833 9562 8834
rect 9534 8807 9535 8833
rect 9535 8807 9561 8833
rect 9561 8807 9562 8833
rect 9534 8806 9562 8807
rect 9478 8246 9506 8274
rect 9366 7294 9394 7322
rect 9422 7209 9450 7210
rect 9422 7183 9423 7209
rect 9423 7183 9449 7209
rect 9449 7183 9450 7209
rect 9422 7182 9450 7183
rect 9702 8694 9730 8722
rect 9758 8553 9786 8554
rect 9758 8527 9759 8553
rect 9759 8527 9785 8553
rect 9785 8527 9786 8553
rect 9758 8526 9786 8527
rect 9918 8637 9946 8638
rect 9918 8611 9919 8637
rect 9919 8611 9945 8637
rect 9945 8611 9946 8637
rect 9918 8610 9946 8611
rect 9970 8637 9998 8638
rect 9970 8611 9971 8637
rect 9971 8611 9997 8637
rect 9997 8611 9998 8637
rect 9970 8610 9998 8611
rect 10022 8637 10050 8638
rect 10022 8611 10023 8637
rect 10023 8611 10049 8637
rect 10049 8611 10050 8637
rect 10022 8610 10050 8611
rect 9870 8246 9898 8274
rect 9982 8078 10010 8106
rect 9918 7853 9946 7854
rect 9918 7827 9919 7853
rect 9919 7827 9945 7853
rect 9945 7827 9946 7853
rect 9918 7826 9946 7827
rect 9970 7853 9998 7854
rect 9970 7827 9971 7853
rect 9971 7827 9997 7853
rect 9997 7827 9998 7853
rect 9970 7826 9998 7827
rect 10022 7853 10050 7854
rect 10022 7827 10023 7853
rect 10023 7827 10049 7853
rect 10049 7827 10050 7853
rect 10022 7826 10050 7827
rect 10430 9225 10458 9226
rect 10430 9199 10431 9225
rect 10431 9199 10457 9225
rect 10457 9199 10458 9225
rect 10430 9198 10458 9199
rect 10654 10737 10682 10738
rect 10654 10711 10655 10737
rect 10655 10711 10681 10737
rect 10681 10711 10682 10737
rect 10654 10710 10682 10711
rect 10766 11241 10794 11242
rect 10766 11215 10767 11241
rect 10767 11215 10793 11241
rect 10793 11215 10794 11241
rect 10766 11214 10794 11215
rect 11102 11185 11130 11186
rect 11102 11159 11103 11185
rect 11103 11159 11129 11185
rect 11129 11159 11130 11185
rect 11102 11158 11130 11159
rect 10990 10934 11018 10962
rect 10934 10905 10962 10906
rect 10934 10879 10935 10905
rect 10935 10879 10961 10905
rect 10961 10879 10962 10905
rect 10934 10878 10962 10879
rect 10654 9505 10682 9506
rect 10654 9479 10655 9505
rect 10655 9479 10681 9505
rect 10681 9479 10682 9505
rect 10654 9478 10682 9479
rect 10878 10654 10906 10682
rect 10822 10486 10850 10514
rect 10990 10430 11018 10458
rect 10822 10262 10850 10290
rect 10766 10206 10794 10234
rect 10822 10150 10850 10178
rect 10990 9870 11018 9898
rect 11158 10934 11186 10962
rect 11550 11494 11578 11522
rect 12614 13145 12642 13146
rect 12614 13119 12615 13145
rect 12615 13119 12641 13145
rect 12641 13119 12642 13145
rect 12614 13118 12642 13119
rect 17598 15301 17626 15302
rect 17598 15275 17599 15301
rect 17599 15275 17625 15301
rect 17625 15275 17626 15301
rect 17598 15274 17626 15275
rect 17650 15301 17678 15302
rect 17650 15275 17651 15301
rect 17651 15275 17677 15301
rect 17677 15275 17678 15301
rect 17650 15274 17678 15275
rect 17702 15301 17730 15302
rect 17702 15275 17703 15301
rect 17703 15275 17729 15301
rect 17729 15275 17730 15301
rect 17702 15274 17730 15275
rect 17598 14517 17626 14518
rect 17598 14491 17599 14517
rect 17599 14491 17625 14517
rect 17625 14491 17626 14517
rect 17598 14490 17626 14491
rect 17650 14517 17678 14518
rect 17650 14491 17651 14517
rect 17651 14491 17677 14517
rect 17677 14491 17678 14517
rect 17650 14490 17678 14491
rect 17702 14517 17730 14518
rect 17702 14491 17703 14517
rect 17703 14491 17729 14517
rect 17729 14491 17730 14517
rect 17702 14490 17730 14491
rect 17598 13733 17626 13734
rect 17598 13707 17599 13733
rect 17599 13707 17625 13733
rect 17625 13707 17626 13733
rect 17598 13706 17626 13707
rect 17650 13733 17678 13734
rect 17650 13707 17651 13733
rect 17651 13707 17677 13733
rect 17677 13707 17678 13733
rect 17650 13706 17678 13707
rect 17702 13733 17730 13734
rect 17702 13707 17703 13733
rect 17703 13707 17729 13733
rect 17729 13707 17730 13733
rect 17702 13706 17730 13707
rect 13566 13622 13594 13650
rect 12950 13174 12978 13202
rect 13454 13454 13482 13482
rect 13174 13118 13202 13146
rect 13174 12838 13202 12866
rect 18830 13622 18858 13650
rect 18830 13145 18858 13146
rect 18830 13119 18831 13145
rect 18831 13119 18857 13145
rect 18857 13119 18858 13145
rect 18830 13118 18858 13119
rect 13454 13062 13482 13090
rect 14126 13089 14154 13090
rect 14126 13063 14127 13089
rect 14127 13063 14153 13089
rect 14153 13063 14154 13089
rect 14126 13062 14154 13063
rect 17598 12949 17626 12950
rect 17598 12923 17599 12949
rect 17599 12923 17625 12949
rect 17625 12923 17626 12949
rect 17598 12922 17626 12923
rect 17650 12949 17678 12950
rect 17650 12923 17651 12949
rect 17651 12923 17677 12949
rect 17677 12923 17678 12949
rect 17650 12922 17678 12923
rect 17702 12949 17730 12950
rect 17702 12923 17703 12949
rect 17703 12923 17729 12949
rect 17729 12923 17730 12949
rect 17702 12922 17730 12923
rect 14462 12838 14490 12866
rect 13566 12697 13594 12698
rect 13566 12671 13567 12697
rect 13567 12671 13593 12697
rect 13593 12671 13594 12697
rect 13566 12670 13594 12671
rect 11718 11942 11746 11970
rect 12894 11662 12922 11690
rect 12334 11577 12362 11578
rect 12334 11551 12335 11577
rect 12335 11551 12361 11577
rect 12361 11551 12362 11577
rect 12334 11550 12362 11551
rect 11942 11521 11970 11522
rect 11942 11495 11943 11521
rect 11943 11495 11969 11521
rect 11969 11495 11970 11521
rect 11942 11494 11970 11495
rect 11606 11270 11634 11298
rect 11718 11326 11746 11354
rect 11046 9590 11074 9618
rect 11102 10710 11130 10738
rect 11102 10094 11130 10122
rect 11158 10289 11186 10290
rect 11158 10263 11159 10289
rect 11159 10263 11185 10289
rect 11185 10263 11186 10289
rect 11158 10262 11186 10263
rect 11158 9982 11186 10010
rect 11326 10766 11354 10794
rect 11438 10793 11466 10794
rect 11438 10767 11439 10793
rect 11439 10767 11465 10793
rect 11465 10767 11466 10793
rect 11438 10766 11466 10767
rect 11382 10710 11410 10738
rect 11494 10654 11522 10682
rect 11326 10150 11354 10178
rect 11326 9982 11354 10010
rect 10766 9422 10794 9450
rect 11158 9198 11186 9226
rect 10542 8806 10570 8834
rect 10878 9142 10906 9170
rect 10710 8105 10738 8106
rect 10710 8079 10711 8105
rect 10711 8079 10737 8105
rect 10737 8079 10738 8105
rect 10710 8078 10738 8079
rect 10990 9142 11018 9170
rect 10990 9030 11018 9058
rect 11102 8806 11130 8834
rect 11830 11297 11858 11298
rect 11830 11271 11831 11297
rect 11831 11271 11857 11297
rect 11857 11271 11858 11297
rect 11830 11270 11858 11271
rect 11774 11129 11802 11130
rect 11774 11103 11775 11129
rect 11775 11103 11801 11129
rect 11801 11103 11802 11129
rect 11774 11102 11802 11103
rect 11830 10990 11858 11018
rect 12670 11577 12698 11578
rect 12670 11551 12671 11577
rect 12671 11551 12697 11577
rect 12697 11551 12698 11577
rect 12670 11550 12698 11551
rect 13062 11577 13090 11578
rect 13062 11551 13063 11577
rect 13063 11551 13089 11577
rect 13089 11551 13090 11577
rect 13062 11550 13090 11551
rect 13230 11326 13258 11354
rect 12614 10934 12642 10962
rect 13398 10766 13426 10794
rect 11550 10150 11578 10178
rect 11382 9870 11410 9898
rect 11270 8974 11298 9002
rect 10934 8302 10962 8330
rect 11270 8441 11298 8442
rect 11270 8415 11271 8441
rect 11271 8415 11297 8441
rect 11297 8415 11298 8441
rect 11270 8414 11298 8415
rect 10318 7966 10346 7994
rect 10654 7993 10682 7994
rect 10654 7967 10655 7993
rect 10655 7967 10681 7993
rect 10681 7967 10682 7993
rect 10654 7966 10682 7967
rect 10878 7910 10906 7938
rect 11606 9310 11634 9338
rect 11494 9225 11522 9226
rect 11494 9199 11495 9225
rect 11495 9199 11521 9225
rect 11521 9199 11522 9225
rect 11494 9198 11522 9199
rect 11718 10065 11746 10066
rect 11718 10039 11719 10065
rect 11719 10039 11745 10065
rect 11745 10039 11746 10065
rect 11718 10038 11746 10039
rect 12782 9646 12810 9674
rect 12614 9617 12642 9618
rect 12614 9591 12615 9617
rect 12615 9591 12641 9617
rect 12641 9591 12642 9617
rect 12614 9590 12642 9591
rect 11662 9254 11690 9282
rect 12110 9478 12138 9506
rect 11998 9281 12026 9282
rect 11998 9255 11999 9281
rect 11999 9255 12025 9281
rect 12025 9255 12026 9281
rect 11998 9254 12026 9255
rect 11830 9198 11858 9226
rect 13846 11577 13874 11578
rect 13846 11551 13847 11577
rect 13847 11551 13873 11577
rect 13873 11551 13874 11577
rect 13846 11550 13874 11551
rect 13958 11158 13986 11186
rect 13174 10038 13202 10066
rect 13118 9673 13146 9674
rect 13118 9647 13119 9673
rect 13119 9647 13145 9673
rect 13145 9647 13146 9673
rect 13118 9646 13146 9647
rect 12950 9198 12978 9226
rect 13006 9561 13034 9562
rect 13006 9535 13007 9561
rect 13007 9535 13033 9561
rect 13033 9535 13034 9561
rect 13006 9534 13034 9535
rect 11998 9086 12026 9114
rect 13062 9505 13090 9506
rect 13062 9479 13063 9505
rect 13063 9479 13089 9505
rect 13089 9479 13090 9505
rect 13062 9478 13090 9479
rect 13118 9198 13146 9226
rect 11606 8833 11634 8834
rect 11606 8807 11607 8833
rect 11607 8807 11633 8833
rect 11633 8807 11634 8833
rect 11606 8806 11634 8807
rect 13566 10065 13594 10066
rect 13566 10039 13567 10065
rect 13567 10039 13593 10065
rect 13593 10039 13594 10065
rect 13566 10038 13594 10039
rect 13790 10766 13818 10794
rect 13230 9646 13258 9674
rect 13118 8806 13146 8834
rect 13398 9590 13426 9618
rect 13902 10710 13930 10738
rect 14294 11158 14322 11186
rect 19950 13454 19978 13482
rect 20006 13118 20034 13146
rect 20006 12782 20034 12810
rect 18942 12670 18970 12698
rect 17598 12165 17626 12166
rect 17598 12139 17599 12165
rect 17599 12139 17625 12165
rect 17625 12139 17626 12165
rect 17598 12138 17626 12139
rect 17650 12165 17678 12166
rect 17650 12139 17651 12165
rect 17651 12139 17677 12165
rect 17677 12139 17678 12165
rect 17650 12138 17678 12139
rect 17702 12165 17730 12166
rect 17702 12139 17703 12165
rect 17703 12139 17729 12165
rect 17729 12139 17730 12165
rect 17702 12138 17730 12139
rect 20118 12110 20146 12138
rect 17598 11381 17626 11382
rect 17598 11355 17599 11381
rect 17599 11355 17625 11381
rect 17625 11355 17626 11381
rect 17598 11354 17626 11355
rect 17650 11381 17678 11382
rect 17650 11355 17651 11381
rect 17651 11355 17677 11381
rect 17677 11355 17678 11381
rect 17650 11354 17678 11355
rect 17702 11381 17730 11382
rect 17702 11355 17703 11381
rect 17703 11355 17729 11381
rect 17729 11355 17730 11381
rect 17702 11354 17730 11355
rect 18830 11185 18858 11186
rect 18830 11159 18831 11185
rect 18831 11159 18857 11185
rect 18857 11159 18858 11185
rect 18830 11158 18858 11159
rect 20006 11102 20034 11130
rect 14406 10737 14434 10738
rect 14406 10711 14407 10737
rect 14407 10711 14433 10737
rect 14433 10711 14434 10737
rect 14406 10710 14434 10711
rect 13958 10038 13986 10066
rect 13398 9366 13426 9394
rect 13622 9310 13650 9338
rect 13734 9366 13762 9394
rect 13342 9225 13370 9226
rect 13342 9199 13343 9225
rect 13343 9199 13369 9225
rect 13369 9199 13370 9225
rect 13342 9198 13370 9199
rect 13286 9086 13314 9114
rect 13846 9142 13874 9170
rect 18830 10793 18858 10794
rect 18830 10767 18831 10793
rect 18831 10767 18857 10793
rect 18857 10767 18858 10793
rect 18830 10766 18858 10767
rect 20006 10766 20034 10794
rect 17598 10597 17626 10598
rect 17598 10571 17599 10597
rect 17599 10571 17625 10597
rect 17625 10571 17626 10597
rect 17598 10570 17626 10571
rect 17650 10597 17678 10598
rect 17650 10571 17651 10597
rect 17651 10571 17677 10597
rect 17677 10571 17678 10597
rect 17650 10570 17678 10571
rect 17702 10597 17730 10598
rect 17702 10571 17703 10597
rect 17703 10571 17729 10597
rect 17729 10571 17730 10597
rect 17702 10570 17730 10571
rect 17598 9813 17626 9814
rect 17598 9787 17599 9813
rect 17599 9787 17625 9813
rect 17625 9787 17626 9813
rect 17598 9786 17626 9787
rect 17650 9813 17678 9814
rect 17650 9787 17651 9813
rect 17651 9787 17677 9813
rect 17677 9787 17678 9813
rect 17650 9786 17678 9787
rect 17702 9813 17730 9814
rect 17702 9787 17703 9813
rect 17703 9787 17729 9813
rect 17729 9787 17730 9813
rect 17702 9786 17730 9787
rect 18830 9617 18858 9618
rect 18830 9591 18831 9617
rect 18831 9591 18857 9617
rect 18857 9591 18858 9617
rect 18830 9590 18858 9591
rect 20006 9422 20034 9450
rect 14630 9198 14658 9226
rect 15022 9225 15050 9226
rect 15022 9199 15023 9225
rect 15023 9199 15049 9225
rect 15049 9199 15050 9225
rect 15022 9198 15050 9199
rect 14070 9142 14098 9170
rect 14798 9169 14826 9170
rect 14798 9143 14799 9169
rect 14799 9143 14825 9169
rect 14825 9143 14826 9169
rect 14798 9142 14826 9143
rect 14070 8974 14098 9002
rect 14238 8833 14266 8834
rect 14238 8807 14239 8833
rect 14239 8807 14265 8833
rect 14265 8807 14266 8833
rect 14238 8806 14266 8807
rect 13118 8414 13146 8442
rect 11998 8358 12026 8386
rect 11438 8190 11466 8218
rect 11550 8302 11578 8330
rect 11550 8049 11578 8050
rect 11550 8023 11551 8049
rect 11551 8023 11577 8049
rect 11577 8023 11578 8049
rect 11550 8022 11578 8023
rect 11942 8246 11970 8274
rect 10374 7209 10402 7210
rect 10374 7183 10375 7209
rect 10375 7183 10401 7209
rect 10401 7183 10402 7209
rect 10374 7182 10402 7183
rect 9030 6790 9058 6818
rect 8806 6510 8834 6538
rect 2238 3541 2266 3542
rect 2238 3515 2239 3541
rect 2239 3515 2265 3541
rect 2265 3515 2266 3541
rect 2238 3514 2266 3515
rect 2290 3541 2318 3542
rect 2290 3515 2291 3541
rect 2291 3515 2317 3541
rect 2317 3515 2318 3541
rect 2290 3514 2318 3515
rect 2342 3541 2370 3542
rect 2342 3515 2343 3541
rect 2343 3515 2369 3541
rect 2369 3515 2370 3541
rect 2342 3514 2370 3515
rect 2238 2757 2266 2758
rect 2238 2731 2239 2757
rect 2239 2731 2265 2757
rect 2265 2731 2266 2757
rect 2238 2730 2266 2731
rect 2290 2757 2318 2758
rect 2290 2731 2291 2757
rect 2291 2731 2317 2757
rect 2317 2731 2318 2757
rect 2290 2730 2318 2731
rect 2342 2757 2370 2758
rect 2342 2731 2343 2757
rect 2343 2731 2369 2757
rect 2369 2731 2370 2757
rect 2342 2730 2370 2731
rect 8078 2590 8106 2618
rect 2238 1973 2266 1974
rect 2238 1947 2239 1973
rect 2239 1947 2265 1973
rect 2265 1947 2266 1973
rect 2238 1946 2266 1947
rect 2290 1973 2318 1974
rect 2290 1947 2291 1973
rect 2291 1947 2317 1973
rect 2317 1947 2318 1973
rect 2290 1946 2318 1947
rect 2342 1973 2370 1974
rect 2342 1947 2343 1973
rect 2343 1947 2369 1973
rect 2369 1947 2370 1973
rect 2342 1946 2370 1947
rect 8694 2617 8722 2618
rect 8694 2591 8695 2617
rect 8695 2591 8721 2617
rect 8721 2591 8722 2617
rect 8694 2590 8722 2591
rect 8414 2030 8442 2058
rect 9918 7069 9946 7070
rect 9918 7043 9919 7069
rect 9919 7043 9945 7069
rect 9945 7043 9946 7069
rect 9918 7042 9946 7043
rect 9970 7069 9998 7070
rect 9970 7043 9971 7069
rect 9971 7043 9997 7069
rect 9997 7043 9998 7069
rect 9970 7042 9998 7043
rect 10022 7069 10050 7070
rect 10022 7043 10023 7069
rect 10023 7043 10049 7069
rect 10049 7043 10050 7069
rect 10022 7042 10050 7043
rect 10206 6873 10234 6874
rect 10206 6847 10207 6873
rect 10207 6847 10233 6873
rect 10233 6847 10234 6873
rect 10206 6846 10234 6847
rect 9926 6790 9954 6818
rect 9478 6510 9506 6538
rect 9702 6537 9730 6538
rect 9702 6511 9703 6537
rect 9703 6511 9729 6537
rect 9729 6511 9730 6537
rect 9702 6510 9730 6511
rect 9918 6285 9946 6286
rect 9918 6259 9919 6285
rect 9919 6259 9945 6285
rect 9945 6259 9946 6285
rect 9918 6258 9946 6259
rect 9970 6285 9998 6286
rect 9970 6259 9971 6285
rect 9971 6259 9997 6285
rect 9997 6259 9998 6285
rect 9970 6258 9998 6259
rect 10022 6285 10050 6286
rect 10022 6259 10023 6285
rect 10023 6259 10049 6285
rect 10049 6259 10050 6285
rect 10022 6258 10050 6259
rect 9918 5501 9946 5502
rect 9918 5475 9919 5501
rect 9919 5475 9945 5501
rect 9945 5475 9946 5501
rect 9918 5474 9946 5475
rect 9970 5501 9998 5502
rect 9970 5475 9971 5501
rect 9971 5475 9997 5501
rect 9997 5475 9998 5501
rect 9970 5474 9998 5475
rect 10022 5501 10050 5502
rect 10022 5475 10023 5501
rect 10023 5475 10049 5501
rect 10049 5475 10050 5501
rect 10022 5474 10050 5475
rect 9918 4717 9946 4718
rect 9918 4691 9919 4717
rect 9919 4691 9945 4717
rect 9945 4691 9946 4717
rect 9918 4690 9946 4691
rect 9970 4717 9998 4718
rect 9970 4691 9971 4717
rect 9971 4691 9997 4717
rect 9997 4691 9998 4717
rect 9970 4690 9998 4691
rect 10022 4717 10050 4718
rect 10022 4691 10023 4717
rect 10023 4691 10049 4717
rect 10049 4691 10050 4717
rect 10022 4690 10050 4691
rect 11998 7294 12026 7322
rect 12278 7294 12306 7322
rect 10934 7209 10962 7210
rect 10934 7183 10935 7209
rect 10935 7183 10961 7209
rect 10961 7183 10962 7209
rect 10934 7182 10962 7183
rect 11326 6846 11354 6874
rect 11830 6873 11858 6874
rect 11830 6847 11831 6873
rect 11831 6847 11857 6873
rect 11857 6847 11858 6873
rect 11830 6846 11858 6847
rect 11046 6734 11074 6762
rect 11606 6734 11634 6762
rect 11942 6734 11970 6762
rect 9918 3933 9946 3934
rect 9918 3907 9919 3933
rect 9919 3907 9945 3933
rect 9945 3907 9946 3933
rect 9918 3906 9946 3907
rect 9970 3933 9998 3934
rect 9970 3907 9971 3933
rect 9971 3907 9997 3933
rect 9997 3907 9998 3933
rect 9970 3906 9998 3907
rect 10022 3933 10050 3934
rect 10022 3907 10023 3933
rect 10023 3907 10049 3933
rect 10049 3907 10050 3933
rect 10022 3906 10050 3907
rect 9918 3149 9946 3150
rect 9918 3123 9919 3149
rect 9919 3123 9945 3149
rect 9945 3123 9946 3149
rect 9918 3122 9946 3123
rect 9970 3149 9998 3150
rect 9970 3123 9971 3149
rect 9971 3123 9997 3149
rect 9997 3123 9998 3149
rect 9970 3122 9998 3123
rect 10022 3149 10050 3150
rect 10022 3123 10023 3149
rect 10023 3123 10049 3149
rect 10049 3123 10050 3149
rect 10022 3122 10050 3123
rect 9918 2365 9946 2366
rect 9918 2339 9919 2365
rect 9919 2339 9945 2365
rect 9945 2339 9946 2365
rect 9918 2338 9946 2339
rect 9970 2365 9998 2366
rect 9970 2339 9971 2365
rect 9971 2339 9997 2365
rect 9997 2339 9998 2365
rect 9970 2338 9998 2339
rect 10022 2365 10050 2366
rect 10022 2339 10023 2365
rect 10023 2339 10049 2365
rect 10049 2339 10050 2365
rect 10022 2338 10050 2339
rect 9198 2057 9226 2058
rect 9198 2031 9199 2057
rect 9199 2031 9225 2057
rect 9225 2031 9226 2057
rect 9198 2030 9226 2031
rect 10430 2030 10458 2058
rect 9918 1581 9946 1582
rect 9918 1555 9919 1581
rect 9919 1555 9945 1581
rect 9945 1555 9946 1581
rect 9918 1554 9946 1555
rect 9970 1581 9998 1582
rect 9970 1555 9971 1581
rect 9971 1555 9997 1581
rect 9997 1555 9998 1581
rect 9970 1554 9998 1555
rect 10022 1581 10050 1582
rect 10022 1555 10023 1581
rect 10023 1555 10049 1581
rect 10049 1555 10050 1581
rect 10022 1554 10050 1555
rect 11046 2057 11074 2058
rect 11046 2031 11047 2057
rect 11047 2031 11073 2057
rect 11073 2031 11074 2057
rect 11046 2030 11074 2031
rect 11774 1806 11802 1834
rect 12782 7321 12810 7322
rect 12782 7295 12783 7321
rect 12783 7295 12809 7321
rect 12809 7295 12810 7321
rect 12782 7294 12810 7295
rect 13678 8470 13706 8498
rect 13510 8441 13538 8442
rect 13510 8415 13511 8441
rect 13511 8415 13537 8441
rect 13537 8415 13538 8441
rect 13510 8414 13538 8415
rect 13622 8022 13650 8050
rect 14686 8833 14714 8834
rect 14686 8807 14687 8833
rect 14687 8807 14713 8833
rect 14713 8807 14714 8833
rect 14686 8806 14714 8807
rect 14854 8777 14882 8778
rect 14854 8751 14855 8777
rect 14855 8751 14881 8777
rect 14881 8751 14882 8777
rect 14854 8750 14882 8751
rect 18830 9225 18858 9226
rect 18830 9199 18831 9225
rect 18831 9199 18857 9225
rect 18857 9199 18858 9225
rect 18830 9198 18858 9199
rect 20006 9113 20034 9114
rect 20006 9087 20007 9113
rect 20007 9087 20033 9113
rect 20033 9087 20034 9113
rect 20006 9086 20034 9087
rect 17598 9029 17626 9030
rect 17598 9003 17599 9029
rect 17599 9003 17625 9029
rect 17625 9003 17626 9029
rect 17598 9002 17626 9003
rect 17650 9029 17678 9030
rect 17650 9003 17651 9029
rect 17651 9003 17677 9029
rect 17677 9003 17678 9029
rect 17650 9002 17678 9003
rect 17702 9029 17730 9030
rect 17702 9003 17703 9029
rect 17703 9003 17729 9029
rect 17729 9003 17730 9029
rect 17702 9002 17730 9003
rect 15134 8750 15162 8778
rect 20006 8750 20034 8778
rect 18830 8470 18858 8498
rect 17598 8245 17626 8246
rect 17598 8219 17599 8245
rect 17599 8219 17625 8245
rect 17625 8219 17626 8245
rect 17598 8218 17626 8219
rect 17650 8245 17678 8246
rect 17650 8219 17651 8245
rect 17651 8219 17677 8245
rect 17677 8219 17678 8245
rect 17650 8218 17678 8219
rect 17702 8245 17730 8246
rect 17702 8219 17703 8245
rect 17703 8219 17729 8245
rect 17729 8219 17730 8245
rect 17702 8218 17730 8219
rect 14574 8022 14602 8050
rect 13230 7574 13258 7602
rect 13454 7601 13482 7602
rect 13454 7575 13455 7601
rect 13455 7575 13481 7601
rect 13481 7575 13482 7601
rect 13454 7574 13482 7575
rect 17598 7461 17626 7462
rect 17598 7435 17599 7461
rect 17599 7435 17625 7461
rect 17625 7435 17626 7461
rect 17598 7434 17626 7435
rect 17650 7461 17678 7462
rect 17650 7435 17651 7461
rect 17651 7435 17677 7461
rect 17677 7435 17678 7461
rect 17650 7434 17678 7435
rect 17702 7461 17730 7462
rect 17702 7435 17703 7461
rect 17703 7435 17729 7461
rect 17729 7435 17730 7461
rect 17702 7434 17730 7435
rect 13342 7182 13370 7210
rect 13902 7182 13930 7210
rect 14238 7182 14266 7210
rect 14014 7153 14042 7154
rect 14014 7127 14015 7153
rect 14015 7127 14041 7153
rect 14041 7127 14042 7153
rect 14014 7126 14042 7127
rect 12782 6873 12810 6874
rect 12782 6847 12783 6873
rect 12783 6847 12809 6873
rect 12809 6847 12810 6873
rect 12782 6846 12810 6847
rect 20006 7406 20034 7434
rect 18830 7265 18858 7266
rect 18830 7239 18831 7265
rect 18831 7239 18857 7265
rect 18857 7239 18858 7265
rect 18830 7238 18858 7239
rect 18718 7182 18746 7210
rect 20006 7070 20034 7098
rect 14462 6873 14490 6874
rect 14462 6847 14463 6873
rect 14463 6847 14489 6873
rect 14489 6847 14490 6873
rect 14462 6846 14490 6847
rect 17598 6677 17626 6678
rect 17598 6651 17599 6677
rect 17599 6651 17625 6677
rect 17625 6651 17626 6677
rect 17598 6650 17626 6651
rect 17650 6677 17678 6678
rect 17650 6651 17651 6677
rect 17651 6651 17677 6677
rect 17677 6651 17678 6677
rect 17650 6650 17678 6651
rect 17702 6677 17730 6678
rect 17702 6651 17703 6677
rect 17703 6651 17729 6677
rect 17729 6651 17730 6677
rect 17702 6650 17730 6651
rect 17598 5893 17626 5894
rect 17598 5867 17599 5893
rect 17599 5867 17625 5893
rect 17625 5867 17626 5893
rect 17598 5866 17626 5867
rect 17650 5893 17678 5894
rect 17650 5867 17651 5893
rect 17651 5867 17677 5893
rect 17677 5867 17678 5893
rect 17650 5866 17678 5867
rect 17702 5893 17730 5894
rect 17702 5867 17703 5893
rect 17703 5867 17729 5893
rect 17729 5867 17730 5893
rect 17702 5866 17730 5867
rect 17598 5109 17626 5110
rect 17598 5083 17599 5109
rect 17599 5083 17625 5109
rect 17625 5083 17626 5109
rect 17598 5082 17626 5083
rect 17650 5109 17678 5110
rect 17650 5083 17651 5109
rect 17651 5083 17677 5109
rect 17677 5083 17678 5109
rect 17650 5082 17678 5083
rect 17702 5109 17730 5110
rect 17702 5083 17703 5109
rect 17703 5083 17729 5109
rect 17729 5083 17730 5109
rect 17702 5082 17730 5083
rect 17598 4325 17626 4326
rect 17598 4299 17599 4325
rect 17599 4299 17625 4325
rect 17625 4299 17626 4325
rect 17598 4298 17626 4299
rect 17650 4325 17678 4326
rect 17650 4299 17651 4325
rect 17651 4299 17677 4325
rect 17677 4299 17678 4325
rect 17650 4298 17678 4299
rect 17702 4325 17730 4326
rect 17702 4299 17703 4325
rect 17703 4299 17729 4325
rect 17729 4299 17730 4325
rect 17702 4298 17730 4299
rect 17598 3541 17626 3542
rect 17598 3515 17599 3541
rect 17599 3515 17625 3541
rect 17625 3515 17626 3541
rect 17598 3514 17626 3515
rect 17650 3541 17678 3542
rect 17650 3515 17651 3541
rect 17651 3515 17677 3541
rect 17677 3515 17678 3541
rect 17650 3514 17678 3515
rect 17702 3541 17730 3542
rect 17702 3515 17703 3541
rect 17703 3515 17729 3541
rect 17729 3515 17730 3541
rect 17702 3514 17730 3515
rect 17598 2757 17626 2758
rect 17598 2731 17599 2757
rect 17599 2731 17625 2757
rect 17625 2731 17626 2757
rect 17598 2730 17626 2731
rect 17650 2757 17678 2758
rect 17650 2731 17651 2757
rect 17651 2731 17677 2757
rect 17677 2731 17678 2757
rect 17650 2730 17678 2731
rect 17702 2757 17730 2758
rect 17702 2731 17703 2757
rect 17703 2731 17729 2757
rect 17729 2731 17730 2757
rect 17702 2730 17730 2731
rect 17598 1973 17626 1974
rect 17598 1947 17599 1973
rect 17599 1947 17625 1973
rect 17625 1947 17626 1973
rect 17598 1946 17626 1947
rect 17650 1973 17678 1974
rect 17650 1947 17651 1973
rect 17651 1947 17677 1973
rect 17677 1947 17678 1973
rect 17650 1946 17678 1947
rect 17702 1973 17730 1974
rect 17702 1947 17703 1973
rect 17703 1947 17729 1973
rect 17729 1947 17730 1973
rect 17702 1946 17730 1947
rect 12782 1833 12810 1834
rect 12782 1807 12783 1833
rect 12783 1807 12809 1833
rect 12809 1807 12810 1833
rect 12782 1806 12810 1807
<< metal3 >>
rect 2233 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2375 19222
rect 17593 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17735 19222
rect 9913 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10055 18830
rect 8409 18718 8414 18746
rect 8442 18718 9198 18746
rect 9226 18718 9231 18746
rect 10761 18718 10766 18746
rect 10794 18718 11382 18746
rect 11410 18718 11415 18746
rect 2233 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2375 18438
rect 17593 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17735 18438
rect 9913 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10055 18046
rect 2233 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2375 17654
rect 17593 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17735 17654
rect 9913 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10055 17262
rect 2233 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2375 16870
rect 17593 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17735 16870
rect 9913 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10055 16478
rect 2233 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2375 16086
rect 17593 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17735 16086
rect 9913 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10055 15694
rect 2233 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2375 15302
rect 17593 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17735 15302
rect 9913 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10055 14910
rect 2233 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2375 14518
rect 17593 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17735 14518
rect 9913 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10055 14126
rect 2233 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2375 13734
rect 17593 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17735 13734
rect 13561 13622 13566 13650
rect 13594 13622 18830 13650
rect 18858 13622 18863 13650
rect 0 13482 400 13496
rect 20600 13482 21000 13496
rect 0 13454 2086 13482
rect 2114 13454 2119 13482
rect 8073 13454 8078 13482
rect 8106 13454 8694 13482
rect 8722 13454 8727 13482
rect 12609 13454 12614 13482
rect 12642 13454 13454 13482
rect 13482 13454 13487 13482
rect 19945 13454 19950 13482
rect 19978 13454 21000 13482
rect 0 13440 400 13454
rect 20600 13440 21000 13454
rect 9913 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10055 13342
rect 8857 13230 8862 13258
rect 8890 13230 9310 13258
rect 9338 13230 11550 13258
rect 11578 13230 12334 13258
rect 12362 13230 12367 13258
rect 12273 13174 12278 13202
rect 12306 13174 12950 13202
rect 12978 13174 12983 13202
rect 20600 13146 21000 13160
rect 7513 13118 7518 13146
rect 7546 13118 8190 13146
rect 8218 13118 8223 13146
rect 9865 13118 9870 13146
rect 9898 13118 11606 13146
rect 11634 13118 11830 13146
rect 11858 13118 12614 13146
rect 12642 13118 13174 13146
rect 13202 13118 13207 13146
rect 15946 13118 18830 13146
rect 18858 13118 18863 13146
rect 20001 13118 20006 13146
rect 20034 13118 21000 13146
rect 15946 13090 15974 13118
rect 20600 13104 21000 13118
rect 13449 13062 13454 13090
rect 13482 13062 14126 13090
rect 14154 13062 15974 13090
rect 2233 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2375 12950
rect 17593 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17735 12950
rect 13169 12838 13174 12866
rect 13202 12838 14462 12866
rect 14490 12838 14495 12866
rect 20600 12810 21000 12824
rect 20001 12782 20006 12810
rect 20034 12782 21000 12810
rect 20600 12768 21000 12782
rect 7177 12726 7182 12754
rect 7210 12726 7518 12754
rect 7546 12726 7798 12754
rect 7826 12726 8414 12754
rect 8442 12726 8447 12754
rect 9529 12726 9534 12754
rect 9562 12726 10262 12754
rect 10290 12726 10295 12754
rect 10313 12670 10318 12698
rect 10346 12670 11046 12698
rect 11074 12670 11079 12698
rect 13561 12670 13566 12698
rect 13594 12670 18942 12698
rect 18970 12670 18975 12698
rect 10089 12614 10094 12642
rect 10122 12614 10878 12642
rect 10906 12614 10911 12642
rect 10929 12558 10934 12586
rect 10962 12558 11550 12586
rect 11578 12558 11583 12586
rect 9913 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10055 12558
rect 8185 12502 8190 12530
rect 8218 12502 8750 12530
rect 8778 12502 8783 12530
rect 8409 12446 8414 12474
rect 8442 12446 9086 12474
rect 9114 12446 9422 12474
rect 9450 12446 9646 12474
rect 9674 12446 9679 12474
rect 6561 12334 6566 12362
rect 6594 12334 7966 12362
rect 7994 12334 9142 12362
rect 9170 12334 9175 12362
rect 8801 12278 8806 12306
rect 8834 12278 10766 12306
rect 10794 12278 10799 12306
rect 8073 12222 8078 12250
rect 8106 12222 8918 12250
rect 8946 12222 8951 12250
rect 2233 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2375 12166
rect 17593 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17735 12166
rect 20600 12138 21000 12152
rect 20113 12110 20118 12138
rect 20146 12110 21000 12138
rect 20600 12096 21000 12110
rect 5889 12054 5894 12082
rect 5922 12054 10654 12082
rect 10682 12054 10687 12082
rect 10817 11942 10822 11970
rect 10850 11942 11494 11970
rect 11522 11942 11718 11970
rect 11746 11942 11751 11970
rect 10145 11774 10150 11802
rect 10178 11774 10934 11802
rect 10962 11774 10967 11802
rect 9913 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10055 11774
rect 7961 11718 7966 11746
rect 7994 11718 8246 11746
rect 8274 11718 8694 11746
rect 8722 11718 8727 11746
rect 9081 11662 9086 11690
rect 9114 11662 12894 11690
rect 12922 11662 12927 11690
rect 8073 11606 8078 11634
rect 8106 11606 8750 11634
rect 8778 11606 8783 11634
rect 12329 11550 12334 11578
rect 12362 11550 12670 11578
rect 12698 11550 12703 11578
rect 13057 11550 13062 11578
rect 13090 11550 13846 11578
rect 13874 11550 13879 11578
rect 7737 11494 7742 11522
rect 7770 11494 8078 11522
rect 8106 11494 8111 11522
rect 11545 11494 11550 11522
rect 11578 11494 11942 11522
rect 11970 11494 11975 11522
rect 2233 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2375 11382
rect 17593 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17735 11382
rect 11713 11326 11718 11354
rect 11746 11326 13230 11354
rect 13258 11326 13263 11354
rect 8969 11270 8974 11298
rect 9002 11270 10318 11298
rect 10346 11270 10351 11298
rect 11601 11270 11606 11298
rect 11634 11270 11830 11298
rect 11858 11270 11863 11298
rect 8017 11214 8022 11242
rect 8050 11214 10766 11242
rect 10794 11214 10799 11242
rect 7457 11158 7462 11186
rect 7490 11158 7854 11186
rect 7882 11158 7887 11186
rect 8073 11158 8078 11186
rect 8106 11158 8414 11186
rect 8442 11158 8447 11186
rect 8745 11158 8750 11186
rect 8778 11158 9086 11186
rect 9114 11158 9119 11186
rect 9193 11158 9198 11186
rect 9226 11158 10094 11186
rect 10122 11158 10127 11186
rect 10313 11158 10318 11186
rect 10346 11158 10654 11186
rect 10682 11158 11102 11186
rect 11130 11158 11135 11186
rect 13953 11158 13958 11186
rect 13986 11158 14294 11186
rect 14322 11158 18830 11186
rect 18858 11158 18863 11186
rect 20600 11130 21000 11144
rect 7177 11102 7182 11130
rect 7210 11102 8134 11130
rect 8162 11102 8358 11130
rect 8386 11102 9142 11130
rect 9170 11102 9175 11130
rect 10537 11102 10542 11130
rect 10570 11102 11774 11130
rect 11802 11102 11807 11130
rect 20001 11102 20006 11130
rect 20034 11102 21000 11130
rect 20600 11088 21000 11102
rect 10878 10990 11830 11018
rect 11858 10990 11863 11018
rect 9913 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10055 10990
rect 10878 10962 10906 10990
rect 8241 10934 8246 10962
rect 8274 10934 9478 10962
rect 9506 10934 9511 10962
rect 9585 10934 9590 10962
rect 9618 10934 9842 10962
rect 9814 10906 9842 10934
rect 10094 10934 10906 10962
rect 10985 10934 10990 10962
rect 11018 10934 11158 10962
rect 11186 10934 11191 10962
rect 11438 10934 12614 10962
rect 12642 10934 12647 10962
rect 10094 10906 10122 10934
rect 5833 10878 5838 10906
rect 5866 10878 7406 10906
rect 7434 10878 7439 10906
rect 7546 10878 8862 10906
rect 8890 10878 8895 10906
rect 9814 10878 10122 10906
rect 10878 10906 10906 10934
rect 10878 10878 10934 10906
rect 10962 10878 10967 10906
rect 7546 10850 7574 10878
rect 7345 10822 7350 10850
rect 7378 10822 7574 10850
rect 7737 10822 7742 10850
rect 7770 10822 9310 10850
rect 9338 10822 9343 10850
rect 11438 10794 11466 10934
rect 20600 10794 21000 10808
rect 8521 10766 8526 10794
rect 8554 10766 8862 10794
rect 8890 10766 8895 10794
rect 11321 10766 11326 10794
rect 11354 10766 11438 10794
rect 11466 10766 11471 10794
rect 13393 10766 13398 10794
rect 13426 10766 13790 10794
rect 13818 10766 13823 10794
rect 15946 10766 18830 10794
rect 18858 10766 18863 10794
rect 20001 10766 20006 10794
rect 20034 10766 21000 10794
rect 15946 10738 15974 10766
rect 20600 10752 21000 10766
rect 10649 10710 10654 10738
rect 10682 10710 11102 10738
rect 11130 10710 11382 10738
rect 11410 10710 11415 10738
rect 13897 10710 13902 10738
rect 13930 10710 14406 10738
rect 14434 10710 15974 10738
rect 10873 10654 10878 10682
rect 10906 10654 11494 10682
rect 11522 10654 11527 10682
rect 2233 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2375 10598
rect 17593 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17735 10598
rect 9305 10486 9310 10514
rect 9338 10486 10206 10514
rect 10234 10486 10822 10514
rect 10850 10486 10855 10514
rect 8017 10430 8022 10458
rect 8050 10430 10990 10458
rect 11018 10430 11023 10458
rect 2137 10374 2142 10402
rect 2170 10374 5334 10402
rect 5362 10374 5367 10402
rect 10817 10262 10822 10290
rect 10850 10262 11158 10290
rect 11186 10262 11191 10290
rect 10313 10206 10318 10234
rect 10346 10206 10766 10234
rect 10794 10206 10799 10234
rect 9913 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10055 10206
rect 10817 10150 10822 10178
rect 10850 10150 11326 10178
rect 11354 10150 11550 10178
rect 11578 10150 11583 10178
rect 0 10122 400 10136
rect 0 10094 966 10122
rect 994 10094 999 10122
rect 7910 10094 8694 10122
rect 8722 10094 8727 10122
rect 8913 10094 8918 10122
rect 8946 10094 11102 10122
rect 11130 10094 11135 10122
rect 0 10080 400 10094
rect 7910 10066 7938 10094
rect 7905 10038 7910 10066
rect 7938 10038 7943 10066
rect 8353 10038 8358 10066
rect 8386 10038 8862 10066
rect 8890 10038 9142 10066
rect 9170 10038 9175 10066
rect 10033 10038 10038 10066
rect 10066 10038 11718 10066
rect 11746 10038 11751 10066
rect 13169 10038 13174 10066
rect 13202 10038 13566 10066
rect 13594 10038 13958 10066
rect 13986 10038 13991 10066
rect 7009 9982 7014 10010
rect 7042 9982 7406 10010
rect 7434 9982 7439 10010
rect 9025 9982 9030 10010
rect 9058 9982 9366 10010
rect 9394 9982 10262 10010
rect 10290 9982 10295 10010
rect 11153 9982 11158 10010
rect 11186 9982 11326 10010
rect 11354 9982 11359 10010
rect 2081 9926 2086 9954
rect 2114 9926 9534 9954
rect 9562 9926 9567 9954
rect 7546 9870 7686 9898
rect 7714 9870 7719 9898
rect 10985 9870 10990 9898
rect 11018 9870 11382 9898
rect 11410 9870 11415 9898
rect 7546 9842 7574 9870
rect 5329 9814 5334 9842
rect 5362 9814 7574 9842
rect 2233 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2375 9814
rect 17593 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17735 9814
rect 6113 9758 6118 9786
rect 6146 9758 6734 9786
rect 6762 9758 6767 9786
rect 6225 9646 6230 9674
rect 6258 9646 7182 9674
rect 7210 9646 7215 9674
rect 7625 9646 7630 9674
rect 7658 9646 10206 9674
rect 10234 9646 12782 9674
rect 12810 9646 13118 9674
rect 13146 9646 13230 9674
rect 13258 9646 13263 9674
rect 7569 9590 7574 9618
rect 7602 9590 7966 9618
rect 7994 9590 7999 9618
rect 11041 9590 11046 9618
rect 11074 9590 12614 9618
rect 12642 9590 13398 9618
rect 13426 9590 13431 9618
rect 15946 9590 18830 9618
rect 18858 9590 18863 9618
rect 15946 9562 15974 9590
rect 13001 9534 13006 9562
rect 13034 9534 15974 9562
rect 7961 9478 7966 9506
rect 7994 9478 9030 9506
rect 9058 9478 9063 9506
rect 9249 9478 9254 9506
rect 9282 9478 10654 9506
rect 10682 9478 10687 9506
rect 12105 9478 12110 9506
rect 12138 9478 13062 9506
rect 13090 9478 13095 9506
rect 10654 9450 10682 9478
rect 20600 9450 21000 9464
rect 10654 9422 10766 9450
rect 10794 9422 10799 9450
rect 20001 9422 20006 9450
rect 20034 9422 21000 9450
rect 9913 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10055 9422
rect 20600 9408 21000 9422
rect 6953 9366 6958 9394
rect 6986 9366 7182 9394
rect 7210 9366 7215 9394
rect 13393 9366 13398 9394
rect 13426 9366 13734 9394
rect 13762 9366 13767 9394
rect 8353 9310 8358 9338
rect 8386 9310 8694 9338
rect 8722 9310 8974 9338
rect 9002 9310 9007 9338
rect 9193 9310 9198 9338
rect 9226 9310 9590 9338
rect 9618 9310 9814 9338
rect 9842 9310 9982 9338
rect 10010 9310 10015 9338
rect 11601 9310 11606 9338
rect 11634 9310 13622 9338
rect 13650 9310 13655 9338
rect 6897 9254 6902 9282
rect 6930 9254 6986 9282
rect 8633 9254 8638 9282
rect 8666 9254 9926 9282
rect 9954 9254 9959 9282
rect 11657 9254 11662 9282
rect 11690 9254 11998 9282
rect 12026 9254 12031 9282
rect 6958 9226 6986 9254
rect 2137 9198 2142 9226
rect 2170 9198 4214 9226
rect 6225 9198 6230 9226
rect 6258 9198 6846 9226
rect 6874 9198 6879 9226
rect 6958 9198 7798 9226
rect 7826 9198 7831 9226
rect 10425 9198 10430 9226
rect 10458 9198 11158 9226
rect 11186 9198 11494 9226
rect 11522 9198 11830 9226
rect 11858 9198 11863 9226
rect 12945 9198 12950 9226
rect 12978 9198 13118 9226
rect 13146 9198 13342 9226
rect 13370 9198 14630 9226
rect 14658 9198 15022 9226
rect 15050 9198 15055 9226
rect 15946 9198 18830 9226
rect 18858 9198 18863 9226
rect 4186 9170 4214 9198
rect 15946 9170 15974 9198
rect 4186 9142 5166 9170
rect 5194 9142 5199 9170
rect 6617 9142 6622 9170
rect 6650 9142 7014 9170
rect 7042 9142 7238 9170
rect 7266 9142 7271 9170
rect 8409 9142 8414 9170
rect 8442 9142 8974 9170
rect 9002 9142 10878 9170
rect 10906 9142 10911 9170
rect 10985 9142 10990 9170
rect 11018 9142 13846 9170
rect 13874 9142 13879 9170
rect 14065 9142 14070 9170
rect 14098 9142 14798 9170
rect 14826 9142 15974 9170
rect 0 9114 400 9128
rect 20600 9114 21000 9128
rect 0 9086 966 9114
rect 994 9086 999 9114
rect 9977 9086 9982 9114
rect 10010 9086 11998 9114
rect 12026 9086 13286 9114
rect 13314 9086 13454 9114
rect 20001 9086 20006 9114
rect 20034 9086 21000 9114
rect 0 9072 400 9086
rect 9753 9030 9758 9058
rect 9786 9030 10990 9058
rect 11018 9030 11023 9058
rect 2233 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2375 9030
rect 13426 9002 13454 9086
rect 20600 9072 21000 9086
rect 17593 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17735 9030
rect 8353 8974 8358 9002
rect 8386 8974 8582 9002
rect 8610 8974 11270 9002
rect 11298 8974 11303 9002
rect 13426 8974 14070 9002
rect 14098 8974 14103 9002
rect 9529 8806 9534 8834
rect 9562 8806 10542 8834
rect 10570 8806 11102 8834
rect 11130 8806 11135 8834
rect 11601 8806 11606 8834
rect 11634 8806 13118 8834
rect 13146 8806 13151 8834
rect 14233 8806 14238 8834
rect 14266 8806 14686 8834
rect 14714 8806 14719 8834
rect 20600 8778 21000 8792
rect 5161 8750 5166 8778
rect 5194 8750 6790 8778
rect 6818 8750 6823 8778
rect 8297 8750 8302 8778
rect 8330 8750 9366 8778
rect 9394 8750 9399 8778
rect 14849 8750 14854 8778
rect 14882 8750 15134 8778
rect 15162 8750 15167 8778
rect 20001 8750 20006 8778
rect 20034 8750 21000 8778
rect 9366 8722 9394 8750
rect 20600 8736 21000 8750
rect 7345 8694 7350 8722
rect 7378 8694 8246 8722
rect 8274 8694 8279 8722
rect 8409 8694 8414 8722
rect 8442 8694 8918 8722
rect 8946 8694 8951 8722
rect 9366 8694 9702 8722
rect 9730 8694 9735 8722
rect 8414 8666 8442 8694
rect 7849 8638 7854 8666
rect 7882 8638 8442 8666
rect 9913 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10055 8638
rect 7014 8582 7686 8610
rect 7714 8582 9142 8610
rect 9170 8582 9175 8610
rect 7014 8554 7042 8582
rect 6729 8526 6734 8554
rect 6762 8526 7014 8554
rect 7042 8526 7047 8554
rect 7121 8526 7126 8554
rect 7154 8526 7742 8554
rect 7770 8526 7775 8554
rect 9081 8526 9086 8554
rect 9114 8526 9758 8554
rect 9786 8526 9791 8554
rect 6561 8470 6566 8498
rect 6594 8470 7462 8498
rect 7490 8470 7495 8498
rect 13673 8470 13678 8498
rect 13706 8470 18830 8498
rect 18858 8470 18863 8498
rect 2137 8414 2142 8442
rect 2170 8414 5502 8442
rect 5530 8414 6874 8442
rect 6953 8414 6958 8442
rect 6986 8414 7294 8442
rect 7322 8414 7327 8442
rect 11265 8414 11270 8442
rect 11298 8414 11303 8442
rect 13113 8414 13118 8442
rect 13146 8414 13510 8442
rect 13538 8414 13543 8442
rect 6846 8386 6874 8414
rect 11270 8386 11298 8414
rect 6846 8358 6902 8386
rect 6930 8358 6935 8386
rect 11270 8358 11998 8386
rect 12026 8358 12031 8386
rect 10929 8302 10934 8330
rect 10962 8302 11550 8330
rect 11578 8302 11583 8330
rect 9473 8246 9478 8274
rect 9506 8246 9870 8274
rect 9898 8246 11942 8274
rect 11970 8246 11975 8274
rect 2233 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2375 8246
rect 17593 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17735 8246
rect 6841 8190 6846 8218
rect 6874 8190 11438 8218
rect 11466 8190 11471 8218
rect 0 8106 400 8120
rect 0 8078 966 8106
rect 994 8078 999 8106
rect 7121 8078 7126 8106
rect 7154 8078 7798 8106
rect 7826 8078 7831 8106
rect 9977 8078 9982 8106
rect 10010 8078 10710 8106
rect 10738 8078 10743 8106
rect 0 8064 400 8078
rect 11545 8022 11550 8050
rect 11578 8022 13622 8050
rect 13650 8022 14574 8050
rect 14602 8022 14607 8050
rect 10313 7966 10318 7994
rect 10346 7966 10654 7994
rect 10682 7966 10687 7994
rect 10654 7938 10682 7966
rect 10654 7910 10878 7938
rect 10906 7910 10911 7938
rect 9913 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10055 7854
rect 13225 7574 13230 7602
rect 13258 7574 13454 7602
rect 13482 7574 13487 7602
rect 7289 7518 7294 7546
rect 7322 7518 8358 7546
rect 8386 7518 8391 7546
rect 2233 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2375 7462
rect 17593 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17735 7462
rect 20600 7434 21000 7448
rect 20001 7406 20006 7434
rect 20034 7406 21000 7434
rect 20600 7392 21000 7406
rect 8073 7350 8078 7378
rect 8106 7350 8750 7378
rect 8778 7350 8783 7378
rect 8521 7294 8526 7322
rect 8554 7294 9366 7322
rect 9394 7294 9399 7322
rect 11993 7294 11998 7322
rect 12026 7294 12278 7322
rect 12306 7294 12782 7322
rect 12810 7294 12815 7322
rect 8185 7238 8190 7266
rect 8218 7238 8414 7266
rect 8442 7238 8447 7266
rect 18825 7238 18830 7266
rect 18858 7238 18863 7266
rect 7345 7182 7350 7210
rect 7378 7182 7910 7210
rect 7938 7182 7943 7210
rect 8857 7182 8862 7210
rect 8890 7182 9422 7210
rect 9450 7182 9455 7210
rect 10369 7182 10374 7210
rect 10402 7182 10934 7210
rect 10962 7182 10967 7210
rect 13337 7182 13342 7210
rect 13370 7182 13902 7210
rect 13930 7182 14238 7210
rect 14266 7182 18718 7210
rect 18746 7182 18751 7210
rect 18830 7154 18858 7238
rect 14009 7126 14014 7154
rect 14042 7126 18858 7154
rect 20600 7098 21000 7112
rect 20001 7070 20006 7098
rect 20034 7070 21000 7098
rect 9913 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10055 7070
rect 20600 7056 21000 7070
rect 10201 6846 10206 6874
rect 10234 6846 11326 6874
rect 11354 6846 11830 6874
rect 11858 6846 12782 6874
rect 12810 6846 14462 6874
rect 14490 6846 14495 6874
rect 8297 6790 8302 6818
rect 8330 6790 8750 6818
rect 8778 6790 9030 6818
rect 9058 6790 9926 6818
rect 9954 6790 9959 6818
rect 11041 6734 11046 6762
rect 11074 6734 11606 6762
rect 11634 6734 11942 6762
rect 11970 6734 11975 6762
rect 2233 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2375 6678
rect 17593 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17735 6678
rect 8801 6510 8806 6538
rect 8834 6510 9478 6538
rect 9506 6510 9702 6538
rect 9730 6510 9735 6538
rect 9913 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10055 6286
rect 2233 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2375 5894
rect 17593 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17735 5894
rect 9913 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10055 5502
rect 2233 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2375 5110
rect 17593 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17735 5110
rect 9913 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10055 4718
rect 2233 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2375 4326
rect 17593 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17735 4326
rect 9913 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10055 3934
rect 2233 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2375 3542
rect 17593 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17735 3542
rect 9913 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10055 3150
rect 2233 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2375 2758
rect 17593 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17735 2758
rect 8073 2590 8078 2618
rect 8106 2590 8694 2618
rect 8722 2590 8727 2618
rect 9913 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10055 2366
rect 8409 2030 8414 2058
rect 8442 2030 9198 2058
rect 9226 2030 9231 2058
rect 10425 2030 10430 2058
rect 10458 2030 11046 2058
rect 11074 2030 11079 2058
rect 2233 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2375 1974
rect 17593 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17735 1974
rect 11769 1806 11774 1834
rect 11802 1806 12782 1834
rect 12810 1806 12815 1834
rect 9913 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10055 1582
<< via3 >>
rect 2238 19194 2266 19222
rect 2290 19194 2318 19222
rect 2342 19194 2370 19222
rect 17598 19194 17626 19222
rect 17650 19194 17678 19222
rect 17702 19194 17730 19222
rect 9918 18802 9946 18830
rect 9970 18802 9998 18830
rect 10022 18802 10050 18830
rect 2238 18410 2266 18438
rect 2290 18410 2318 18438
rect 2342 18410 2370 18438
rect 17598 18410 17626 18438
rect 17650 18410 17678 18438
rect 17702 18410 17730 18438
rect 9918 18018 9946 18046
rect 9970 18018 9998 18046
rect 10022 18018 10050 18046
rect 2238 17626 2266 17654
rect 2290 17626 2318 17654
rect 2342 17626 2370 17654
rect 17598 17626 17626 17654
rect 17650 17626 17678 17654
rect 17702 17626 17730 17654
rect 9918 17234 9946 17262
rect 9970 17234 9998 17262
rect 10022 17234 10050 17262
rect 2238 16842 2266 16870
rect 2290 16842 2318 16870
rect 2342 16842 2370 16870
rect 17598 16842 17626 16870
rect 17650 16842 17678 16870
rect 17702 16842 17730 16870
rect 9918 16450 9946 16478
rect 9970 16450 9998 16478
rect 10022 16450 10050 16478
rect 2238 16058 2266 16086
rect 2290 16058 2318 16086
rect 2342 16058 2370 16086
rect 17598 16058 17626 16086
rect 17650 16058 17678 16086
rect 17702 16058 17730 16086
rect 9918 15666 9946 15694
rect 9970 15666 9998 15694
rect 10022 15666 10050 15694
rect 2238 15274 2266 15302
rect 2290 15274 2318 15302
rect 2342 15274 2370 15302
rect 17598 15274 17626 15302
rect 17650 15274 17678 15302
rect 17702 15274 17730 15302
rect 9918 14882 9946 14910
rect 9970 14882 9998 14910
rect 10022 14882 10050 14910
rect 2238 14490 2266 14518
rect 2290 14490 2318 14518
rect 2342 14490 2370 14518
rect 17598 14490 17626 14518
rect 17650 14490 17678 14518
rect 17702 14490 17730 14518
rect 9918 14098 9946 14126
rect 9970 14098 9998 14126
rect 10022 14098 10050 14126
rect 2238 13706 2266 13734
rect 2290 13706 2318 13734
rect 2342 13706 2370 13734
rect 17598 13706 17626 13734
rect 17650 13706 17678 13734
rect 17702 13706 17730 13734
rect 9918 13314 9946 13342
rect 9970 13314 9998 13342
rect 10022 13314 10050 13342
rect 2238 12922 2266 12950
rect 2290 12922 2318 12950
rect 2342 12922 2370 12950
rect 17598 12922 17626 12950
rect 17650 12922 17678 12950
rect 17702 12922 17730 12950
rect 9918 12530 9946 12558
rect 9970 12530 9998 12558
rect 10022 12530 10050 12558
rect 2238 12138 2266 12166
rect 2290 12138 2318 12166
rect 2342 12138 2370 12166
rect 17598 12138 17626 12166
rect 17650 12138 17678 12166
rect 17702 12138 17730 12166
rect 9918 11746 9946 11774
rect 9970 11746 9998 11774
rect 10022 11746 10050 11774
rect 2238 11354 2266 11382
rect 2290 11354 2318 11382
rect 2342 11354 2370 11382
rect 17598 11354 17626 11382
rect 17650 11354 17678 11382
rect 17702 11354 17730 11382
rect 9918 10962 9946 10990
rect 9970 10962 9998 10990
rect 10022 10962 10050 10990
rect 2238 10570 2266 10598
rect 2290 10570 2318 10598
rect 2342 10570 2370 10598
rect 17598 10570 17626 10598
rect 17650 10570 17678 10598
rect 17702 10570 17730 10598
rect 9918 10178 9946 10206
rect 9970 10178 9998 10206
rect 10022 10178 10050 10206
rect 2238 9786 2266 9814
rect 2290 9786 2318 9814
rect 2342 9786 2370 9814
rect 17598 9786 17626 9814
rect 17650 9786 17678 9814
rect 17702 9786 17730 9814
rect 9918 9394 9946 9422
rect 9970 9394 9998 9422
rect 10022 9394 10050 9422
rect 2238 9002 2266 9030
rect 2290 9002 2318 9030
rect 2342 9002 2370 9030
rect 17598 9002 17626 9030
rect 17650 9002 17678 9030
rect 17702 9002 17730 9030
rect 9918 8610 9946 8638
rect 9970 8610 9998 8638
rect 10022 8610 10050 8638
rect 2238 8218 2266 8246
rect 2290 8218 2318 8246
rect 2342 8218 2370 8246
rect 17598 8218 17626 8246
rect 17650 8218 17678 8246
rect 17702 8218 17730 8246
rect 9918 7826 9946 7854
rect 9970 7826 9998 7854
rect 10022 7826 10050 7854
rect 2238 7434 2266 7462
rect 2290 7434 2318 7462
rect 2342 7434 2370 7462
rect 17598 7434 17626 7462
rect 17650 7434 17678 7462
rect 17702 7434 17730 7462
rect 9918 7042 9946 7070
rect 9970 7042 9998 7070
rect 10022 7042 10050 7070
rect 2238 6650 2266 6678
rect 2290 6650 2318 6678
rect 2342 6650 2370 6678
rect 17598 6650 17626 6678
rect 17650 6650 17678 6678
rect 17702 6650 17730 6678
rect 9918 6258 9946 6286
rect 9970 6258 9998 6286
rect 10022 6258 10050 6286
rect 2238 5866 2266 5894
rect 2290 5866 2318 5894
rect 2342 5866 2370 5894
rect 17598 5866 17626 5894
rect 17650 5866 17678 5894
rect 17702 5866 17730 5894
rect 9918 5474 9946 5502
rect 9970 5474 9998 5502
rect 10022 5474 10050 5502
rect 2238 5082 2266 5110
rect 2290 5082 2318 5110
rect 2342 5082 2370 5110
rect 17598 5082 17626 5110
rect 17650 5082 17678 5110
rect 17702 5082 17730 5110
rect 9918 4690 9946 4718
rect 9970 4690 9998 4718
rect 10022 4690 10050 4718
rect 2238 4298 2266 4326
rect 2290 4298 2318 4326
rect 2342 4298 2370 4326
rect 17598 4298 17626 4326
rect 17650 4298 17678 4326
rect 17702 4298 17730 4326
rect 9918 3906 9946 3934
rect 9970 3906 9998 3934
rect 10022 3906 10050 3934
rect 2238 3514 2266 3542
rect 2290 3514 2318 3542
rect 2342 3514 2370 3542
rect 17598 3514 17626 3542
rect 17650 3514 17678 3542
rect 17702 3514 17730 3542
rect 9918 3122 9946 3150
rect 9970 3122 9998 3150
rect 10022 3122 10050 3150
rect 2238 2730 2266 2758
rect 2290 2730 2318 2758
rect 2342 2730 2370 2758
rect 17598 2730 17626 2758
rect 17650 2730 17678 2758
rect 17702 2730 17730 2758
rect 9918 2338 9946 2366
rect 9970 2338 9998 2366
rect 10022 2338 10050 2366
rect 2238 1946 2266 1974
rect 2290 1946 2318 1974
rect 2342 1946 2370 1974
rect 17598 1946 17626 1974
rect 17650 1946 17678 1974
rect 17702 1946 17730 1974
rect 9918 1554 9946 1582
rect 9970 1554 9998 1582
rect 10022 1554 10050 1582
<< metal4 >>
rect 2224 19222 2384 19238
rect 2224 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2384 19222
rect 2224 18438 2384 19194
rect 2224 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2384 18438
rect 2224 17654 2384 18410
rect 2224 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2384 17654
rect 2224 16870 2384 17626
rect 2224 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2384 16870
rect 2224 16086 2384 16842
rect 2224 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2384 16086
rect 2224 15302 2384 16058
rect 2224 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2384 15302
rect 2224 14518 2384 15274
rect 2224 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2384 14518
rect 2224 13734 2384 14490
rect 2224 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2384 13734
rect 2224 12950 2384 13706
rect 2224 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2384 12950
rect 2224 12166 2384 12922
rect 2224 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2384 12166
rect 2224 11382 2384 12138
rect 2224 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2384 11382
rect 2224 10598 2384 11354
rect 2224 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2384 10598
rect 2224 9814 2384 10570
rect 2224 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2384 9814
rect 2224 9030 2384 9786
rect 2224 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2384 9030
rect 2224 8246 2384 9002
rect 2224 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2384 8246
rect 2224 7462 2384 8218
rect 2224 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2384 7462
rect 2224 6678 2384 7434
rect 2224 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2384 6678
rect 2224 5894 2384 6650
rect 2224 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2384 5894
rect 2224 5110 2384 5866
rect 2224 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2384 5110
rect 2224 4326 2384 5082
rect 2224 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2384 4326
rect 2224 3542 2384 4298
rect 2224 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2384 3542
rect 2224 2758 2384 3514
rect 2224 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2384 2758
rect 2224 1974 2384 2730
rect 2224 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2384 1974
rect 2224 1538 2384 1946
rect 9904 18830 10064 19238
rect 9904 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10064 18830
rect 9904 18046 10064 18802
rect 9904 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10064 18046
rect 9904 17262 10064 18018
rect 9904 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10064 17262
rect 9904 16478 10064 17234
rect 9904 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10064 16478
rect 9904 15694 10064 16450
rect 9904 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10064 15694
rect 9904 14910 10064 15666
rect 9904 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10064 14910
rect 9904 14126 10064 14882
rect 9904 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10064 14126
rect 9904 13342 10064 14098
rect 9904 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10064 13342
rect 9904 12558 10064 13314
rect 9904 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10064 12558
rect 9904 11774 10064 12530
rect 9904 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10064 11774
rect 9904 10990 10064 11746
rect 9904 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10064 10990
rect 9904 10206 10064 10962
rect 9904 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10064 10206
rect 9904 9422 10064 10178
rect 9904 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10064 9422
rect 9904 8638 10064 9394
rect 9904 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10064 8638
rect 9904 7854 10064 8610
rect 9904 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10064 7854
rect 9904 7070 10064 7826
rect 9904 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10064 7070
rect 9904 6286 10064 7042
rect 9904 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10064 6286
rect 9904 5502 10064 6258
rect 9904 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10064 5502
rect 9904 4718 10064 5474
rect 9904 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10064 4718
rect 9904 3934 10064 4690
rect 9904 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10064 3934
rect 9904 3150 10064 3906
rect 9904 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10064 3150
rect 9904 2366 10064 3122
rect 9904 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10064 2366
rect 9904 1582 10064 2338
rect 9904 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10064 1582
rect 9904 1538 10064 1554
rect 17584 19222 17744 19238
rect 17584 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17744 19222
rect 17584 18438 17744 19194
rect 17584 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17744 18438
rect 17584 17654 17744 18410
rect 17584 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17744 17654
rect 17584 16870 17744 17626
rect 17584 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17744 16870
rect 17584 16086 17744 16842
rect 17584 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17744 16086
rect 17584 15302 17744 16058
rect 17584 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17744 15302
rect 17584 14518 17744 15274
rect 17584 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17744 14518
rect 17584 13734 17744 14490
rect 17584 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17744 13734
rect 17584 12950 17744 13706
rect 17584 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17744 12950
rect 17584 12166 17744 12922
rect 17584 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17744 12166
rect 17584 11382 17744 12138
rect 17584 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17744 11382
rect 17584 10598 17744 11354
rect 17584 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17744 10598
rect 17584 9814 17744 10570
rect 17584 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17744 9814
rect 17584 9030 17744 9786
rect 17584 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17744 9030
rect 17584 8246 17744 9002
rect 17584 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17744 8246
rect 17584 7462 17744 8218
rect 17584 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17744 7462
rect 17584 6678 17744 7434
rect 17584 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17744 6678
rect 17584 5894 17744 6650
rect 17584 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17744 5894
rect 17584 5110 17744 5866
rect 17584 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17744 5110
rect 17584 4326 17744 5082
rect 17584 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17744 4326
rect 17584 3542 17744 4298
rect 17584 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17744 3542
rect 17584 2758 17744 3514
rect 17584 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17744 2758
rect 17584 1974 17744 2730
rect 17584 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17744 1974
rect 17584 1538 17744 1946
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _104_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7672 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _105_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7840 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _106_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _107_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9072 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _108_
timestamp 1698175906
transform 1 0 10024 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _109_
timestamp 1698175906
transform 1 0 10920 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _110_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10920 0 1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _111_
timestamp 1698175906
transform -1 0 11256 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _112_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9912 0 1 10976
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _113_
timestamp 1698175906
transform -1 0 9632 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _114_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9296 0 -1 12544
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _115_
timestamp 1698175906
transform 1 0 8288 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _116_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8960 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _117_
timestamp 1698175906
transform -1 0 10360 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _118_
timestamp 1698175906
transform -1 0 9576 0 -1 13328
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _119_
timestamp 1698175906
transform -1 0 11648 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _120_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10584 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _121_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7392 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _122_
timestamp 1698175906
transform 1 0 8960 0 -1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _123_
timestamp 1698175906
transform 1 0 10584 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _124_
timestamp 1698175906
transform -1 0 8512 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _125_
timestamp 1698175906
transform 1 0 9296 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _126_
timestamp 1698175906
transform -1 0 10808 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _127_
timestamp 1698175906
transform 1 0 11704 0 1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _128_
timestamp 1698175906
transform -1 0 12432 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _129_
timestamp 1698175906
transform 1 0 11536 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _130_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11032 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _131_
timestamp 1698175906
transform 1 0 5768 0 -1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _132_
timestamp 1698175906
transform 1 0 9408 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _133_
timestamp 1698175906
transform -1 0 9352 0 -1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _134_
timestamp 1698175906
transform -1 0 8960 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _135_
timestamp 1698175906
transform 1 0 7952 0 -1 10976
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _136_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 8176 0 -1 9408
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _137_
timestamp 1698175906
transform -1 0 6944 0 1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _138_
timestamp 1698175906
transform -1 0 11424 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _139_
timestamp 1698175906
transform 1 0 11256 0 1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _140_
timestamp 1698175906
transform -1 0 11704 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _141_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8960 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _142_
timestamp 1698175906
transform -1 0 8400 0 -1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _143_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 8400 0 1 10192
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _144_
timestamp 1698175906
transform -1 0 7672 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _145_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7560 0 -1 8624
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _146_
timestamp 1698175906
transform 1 0 8288 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _147_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _148_
timestamp 1698175906
transform -1 0 9632 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _149_
timestamp 1698175906
transform 1 0 9520 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _150_
timestamp 1698175906
transform 1 0 9296 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _151_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 8960 0 1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _152_
timestamp 1698175906
transform 1 0 10192 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _153_
timestamp 1698175906
transform -1 0 11032 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _154_
timestamp 1698175906
transform -1 0 11760 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _155_
timestamp 1698175906
transform -1 0 6944 0 1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _156_
timestamp 1698175906
transform 1 0 6720 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _157_
timestamp 1698175906
transform -1 0 8960 0 1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _158_
timestamp 1698175906
transform -1 0 8288 0 -1 12544
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _159_
timestamp 1698175906
transform 1 0 7952 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _160_
timestamp 1698175906
transform -1 0 8624 0 1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _161_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 8288 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _162_
timestamp 1698175906
transform -1 0 8960 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _163_
timestamp 1698175906
transform 1 0 8232 0 -1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _164_
timestamp 1698175906
transform 1 0 12488 0 1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _165_
timestamp 1698175906
transform 1 0 12544 0 -1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _166_
timestamp 1698175906
transform -1 0 9240 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _167_
timestamp 1698175906
transform -1 0 10080 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _168_
timestamp 1698175906
transform 1 0 10192 0 -1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _169_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10584 0 1 7840
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _170_
timestamp 1698175906
transform 1 0 9576 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _171_
timestamp 1698175906
transform -1 0 8624 0 1 8624
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _172_
timestamp 1698175906
transform -1 0 7224 0 -1 8624
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _173_
timestamp 1698175906
transform 1 0 7224 0 -1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _174_
timestamp 1698175906
transform 1 0 11872 0 1 7840
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _175_
timestamp 1698175906
transform -1 0 11368 0 -1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _176_
timestamp 1698175906
transform 1 0 10584 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _177_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11312 0 1 7840
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _178_
timestamp 1698175906
transform 1 0 11424 0 -1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _179_
timestamp 1698175906
transform 1 0 7840 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _180_
timestamp 1698175906
transform 1 0 10584 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _181_
timestamp 1698175906
transform 1 0 12544 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _182_
timestamp 1698175906
transform 1 0 10808 0 1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _183_
timestamp 1698175906
transform -1 0 10472 0 1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _184_
timestamp 1698175906
transform 1 0 13328 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _185_
timestamp 1698175906
transform 1 0 9856 0 -1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _186_
timestamp 1698175906
transform 1 0 13104 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _187_
timestamp 1698175906
transform 1 0 13104 0 1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _188_
timestamp 1698175906
transform 1 0 13328 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _189_
timestamp 1698175906
transform -1 0 8064 0 -1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai221_1  _190_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 7784 0 -1 10192
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _191_
timestamp 1698175906
transform -1 0 6328 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _192_
timestamp 1698175906
transform 1 0 13720 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _193_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 -1 11760
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _194_
timestamp 1698175906
transform 1 0 12824 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _195_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 14392 0 1 8624
box -43 -43 883 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _196_
timestamp 1698175906
transform 1 0 14504 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _197_
timestamp 1698175906
transform -1 0 15288 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _198_
timestamp 1698175906
transform -1 0 12040 0 1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _199_
timestamp 1698175906
transform -1 0 13216 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _200_
timestamp 1698175906
transform 1 0 11760 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__and4_1  _201_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11032 0 -1 9408
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _202_
timestamp 1698175906
transform 1 0 13832 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _203_
timestamp 1698175906
transform -1 0 13832 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _204_
timestamp 1698175906
transform 1 0 10752 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _205_
timestamp 1698175906
transform 1 0 11256 0 -1 10976
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _206_
timestamp 1698175906
transform 1 0 13664 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _207_
timestamp 1698175906
transform -1 0 13496 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _208_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7728 0 1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _209_
timestamp 1698175906
transform 1 0 9744 0 -1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _210_
timestamp 1698175906
transform 1 0 11424 0 1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _211_
timestamp 1698175906
transform 1 0 6104 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _212_
timestamp 1698175906
transform 1 0 5768 0 -1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _213_
timestamp 1698175906
transform 1 0 5656 0 -1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _214_
timestamp 1698175906
transform -1 0 12432 0 -1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _215_
timestamp 1698175906
transform 1 0 6664 0 1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _216_
timestamp 1698175906
transform 1 0 8176 0 1 6272
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _217_
timestamp 1698175906
transform 1 0 9520 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _218_
timestamp 1698175906
transform -1 0 6720 0 -1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _219_
timestamp 1698175906
transform 1 0 7056 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _220_
timestamp 1698175906
transform 1 0 6888 0 -1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _221_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12544 0 -1 13328
box -43 -43 1779 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _222_
timestamp 1698175906
transform 1 0 9128 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _223_
timestamp 1698175906
transform -1 0 7056 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _224_
timestamp 1698175906
transform 1 0 11256 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _225_
timestamp 1698175906
transform 1 0 10080 0 -1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _226_
timestamp 1698175906
transform 1 0 12712 0 -1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _227_
timestamp 1698175906
transform -1 0 6888 0 -1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _228_
timestamp 1698175906
transform 1 0 12768 0 1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _229_
timestamp 1698175906
transform -1 0 15232 0 -1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _230_
timestamp 1698175906
transform 1 0 11480 0 1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _231_
timestamp 1698175906
transform 1 0 13272 0 -1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _232_
timestamp 1698175906
transform 1 0 12880 0 -1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _235_
timestamp 1698175906
transform 1 0 13776 0 1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _236_
timestamp 1698175906
transform 1 0 13328 0 1 13328
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _237_
timestamp 1698175906
transform 1 0 13328 0 1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__208__CLK dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9744 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__209__CLK
timestamp 1698175906
transform -1 0 11872 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__210__CLK
timestamp 1698175906
transform 1 0 13160 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__211__CLK
timestamp 1698175906
transform 1 0 8400 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__212__CLK
timestamp 1698175906
transform 1 0 7504 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__213__CLK
timestamp 1698175906
transform 1 0 7392 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__214__CLK
timestamp 1698175906
transform 1 0 12656 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__215__CLK
timestamp 1698175906
transform 1 0 8400 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__216__CLK
timestamp 1698175906
transform 1 0 9912 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__217__CLK
timestamp 1698175906
transform 1 0 9408 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__218__CLK
timestamp 1698175906
transform 1 0 7280 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__219__CLK
timestamp 1698175906
transform 1 0 9072 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__220__CLK
timestamp 1698175906
transform 1 0 8736 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__221__CLK
timestamp 1698175906
transform -1 0 14504 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__222__CLK
timestamp 1698175906
transform 1 0 9016 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__223__CLK
timestamp 1698175906
transform 1 0 7168 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__224__CLK
timestamp 1698175906
transform 1 0 12992 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__225__CLK
timestamp 1698175906
transform 1 0 11816 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__226__CLK
timestamp 1698175906
transform 1 0 14448 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__227__CLK
timestamp 1698175906
transform 1 0 7000 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__228__CLK
timestamp 1698175906
transform 1 0 14616 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__229__CLK
timestamp 1698175906
transform 1 0 13496 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__230__CLK
timestamp 1698175906
transform 1 0 13104 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__231__CLK
timestamp 1698175906
transform 1 0 15008 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__232__CLK
timestamp 1698175906
transform 1 0 14616 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform 1 0 9520 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9632 0 -1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 10472 0 1 9408
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 11592 0 1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 2688 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 4592 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 6496 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8400 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_172
timestamp 1698175906
transform 1 0 10304 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_176
timestamp 1698175906
transform 1 0 10528 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_232
timestamp 1698175906
transform 1 0 13664 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_236
timestamp 1698175906
transform 1 0 13888 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_0_240 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 14112 0 1 1568
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_256
timestamp 1698175906
transform 1 0 15008 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_258 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15120 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_263 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15400 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_271
timestamp 1698175906
transform 1 0 15848 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 16016 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 17920 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 19824 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 20048 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348
timestamp 1698175906
transform 1 0 20160 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 4368 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 4704 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 8288 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_168
timestamp 1698175906
transform 1 0 10080 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_172
timestamp 1698175906
transform 1 0 10304 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_174
timestamp 1698175906
transform 1 0 10416 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_201
timestamp 1698175906
transform 1 0 11928 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698175906
transform 1 0 12376 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_212
timestamp 1698175906
transform 1 0 12544 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_276
timestamp 1698175906
transform 1 0 16128 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 16464 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 20048 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 20160 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 784 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 2576 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 2744 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 6328 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_107
timestamp 1698175906
transform 1 0 6664 0 1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_123
timestamp 1698175906
transform 1 0 7560 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_131
timestamp 1698175906
transform 1 0 8008 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_159
timestamp 1698175906
transform 1 0 9576 0 1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698175906
transform 1 0 10584 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 14168 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 14504 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 18088 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 18424 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 784 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 4368 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 4704 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 8288 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 8624 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 12208 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 12544 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 16128 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 16464 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 20048 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 20160 0 -1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 784 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 2576 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 2744 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 6328 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 6664 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 10248 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 10584 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 14168 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 14504 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 18088 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 18424 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 784 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 4368 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 4704 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 8288 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 8624 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 12208 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 12544 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 16128 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 16464 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 20048 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 20160 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 784 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 2576 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 2744 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 6328 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 6664 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 10248 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 10584 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 14168 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 14504 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 18088 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 18424 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 784 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 4368 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 4704 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 8288 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 8624 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 12208 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 12544 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 16128 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 16464 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 20048 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 20160 0 -1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 784 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 2576 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 2744 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 6328 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 6664 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 10248 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 10584 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 14168 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 14504 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 18088 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 18424 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 784 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 4368 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 4704 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 8288 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 8624 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 12208 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 12544 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 16128 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 16464 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 20048 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 20160 0 -1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 784 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 2576 0 1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 2744 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 6328 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 6664 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 10248 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 10584 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 14168 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 14504 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 18088 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 18424 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 784 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 4368 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 4704 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 8288 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 8624 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 12208 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 12544 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 16128 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 16464 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 20048 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 20160 0 -1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 784 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 2576 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 2744 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 6328 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_107
timestamp 1698175906
transform 1 0 6664 0 1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_123
timestamp 1698175906
transform 1 0 7560 0 1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_131
timestamp 1698175906
transform 1 0 8008 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_133
timestamp 1698175906
transform 1 0 8120 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_163
timestamp 1698175906
transform 1 0 9800 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_167
timestamp 1698175906
transform 1 0 10024 0 1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_177
timestamp 1698175906
transform 1 0 10584 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698175906
transform 1 0 14168 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 14504 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 18088 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 18424 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 784 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 4368 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_72
timestamp 1698175906
transform 1 0 4704 0 -1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_104
timestamp 1698175906
transform 1 0 6496 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_108
timestamp 1698175906
transform 1 0 6720 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_110
timestamp 1698175906
transform 1 0 6832 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_142
timestamp 1698175906
transform 1 0 8624 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_146
timestamp 1698175906
transform 1 0 8848 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_162
timestamp 1698175906
transform 1 0 9744 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_166
timestamp 1698175906
transform 1 0 9968 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_197
timestamp 1698175906
transform 1 0 11704 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_201
timestamp 1698175906
transform 1 0 11928 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_209
timestamp 1698175906
transform 1 0 12376 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_212
timestamp 1698175906
transform 1 0 12544 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_214
timestamp 1698175906
transform 1 0 12656 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_244
timestamp 1698175906
transform 1 0 14336 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_248
timestamp 1698175906
transform 1 0 14560 0 -1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 16464 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 20048 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 20160 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 784 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 2576 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 2744 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 6328 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_107
timestamp 1698175906
transform 1 0 6664 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_123
timestamp 1698175906
transform 1 0 7560 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_127
timestamp 1698175906
transform 1 0 7784 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_148
timestamp 1698175906
transform 1 0 8960 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_152
timestamp 1698175906
transform 1 0 9184 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_162
timestamp 1698175906
transform 1 0 9744 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_166
timestamp 1698175906
transform 1 0 9968 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_168
timestamp 1698175906
transform 1 0 10080 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_177
timestamp 1698175906
transform 1 0 10584 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_187
timestamp 1698175906
transform 1 0 11144 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_218
timestamp 1698175906
transform 1 0 12880 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_228
timestamp 1698175906
transform 1 0 13440 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_232
timestamp 1698175906
transform 1 0 13664 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_240
timestamp 1698175906
transform 1 0 14112 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_244
timestamp 1698175906
transform 1 0 14336 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 14504 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 18088 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_317
timestamp 1698175906
transform 1 0 18424 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_321
timestamp 1698175906
transform 1 0 18648 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 784 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 4368 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_72
timestamp 1698175906
transform 1 0 4704 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_80
timestamp 1698175906
transform 1 0 5152 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_84
timestamp 1698175906
transform 1 0 5376 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_114
timestamp 1698175906
transform 1 0 7056 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_118
timestamp 1698175906
transform 1 0 7280 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_134
timestamp 1698175906
transform 1 0 8176 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_138
timestamp 1698175906
transform 1 0 8400 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_142
timestamp 1698175906
transform 1 0 8624 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_146
timestamp 1698175906
transform 1 0 8848 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_148
timestamp 1698175906
transform 1 0 8960 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_180
timestamp 1698175906
transform 1 0 10752 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_188
timestamp 1698175906
transform 1 0 11200 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_198
timestamp 1698175906
transform 1 0 11760 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_206
timestamp 1698175906
transform 1 0 12208 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_212
timestamp 1698175906
transform 1 0 12544 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_220
timestamp 1698175906
transform 1 0 12992 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_224
timestamp 1698175906
transform 1 0 13216 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_234
timestamp 1698175906
transform 1 0 13776 0 -1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_266
timestamp 1698175906
transform 1 0 15568 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_274
timestamp 1698175906
transform 1 0 16016 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_278
timestamp 1698175906
transform 1 0 16240 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_282
timestamp 1698175906
transform 1 0 16464 0 -1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_314
timestamp 1698175906
transform 1 0 18256 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_322
timestamp 1698175906
transform 1 0 18704 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 784 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 2576 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 2744 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 6328 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_136
timestamp 1698175906
transform 1 0 8288 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_140
timestamp 1698175906
transform 1 0 8512 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_172
timestamp 1698175906
transform 1 0 10304 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_174
timestamp 1698175906
transform 1 0 10416 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_187
timestamp 1698175906
transform 1 0 11144 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_189
timestamp 1698175906
transform 1 0 11256 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_205
timestamp 1698175906
transform 1 0 12152 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_237
timestamp 1698175906
transform 1 0 13944 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 14504 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 18088 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_317
timestamp 1698175906
transform 1 0 18424 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_28
timestamp 1698175906
transform 1 0 2240 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_60
timestamp 1698175906
transform 1 0 4032 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_68
timestamp 1698175906
transform 1 0 4480 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_72
timestamp 1698175906
transform 1 0 4704 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_104
timestamp 1698175906
transform 1 0 6496 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_122
timestamp 1698175906
transform 1 0 7504 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_132
timestamp 1698175906
transform 1 0 8064 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_138
timestamp 1698175906
transform 1 0 8400 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_142
timestamp 1698175906
transform 1 0 8624 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_158
timestamp 1698175906
transform 1 0 9520 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_167
timestamp 1698175906
transform 1 0 10024 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_183
timestamp 1698175906
transform 1 0 10920 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_185
timestamp 1698175906
transform 1 0 11032 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_191
timestamp 1698175906
transform 1 0 11368 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_207
timestamp 1698175906
transform 1 0 12264 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1698175906
transform 1 0 12376 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_212
timestamp 1698175906
transform 1 0 12544 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_220
timestamp 1698175906
transform 1 0 12992 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_224
timestamp 1698175906
transform 1 0 13216 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_228
timestamp 1698175906
transform 1 0 13440 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_260
timestamp 1698175906
transform 1 0 15232 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_276
timestamp 1698175906
transform 1 0 16128 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_282
timestamp 1698175906
transform 1 0 16464 0 -1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_346
timestamp 1698175906
transform 1 0 20048 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_348
timestamp 1698175906
transform 1 0 20160 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698175906
transform 1 0 784 0 1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 2576 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698175906
transform 1 0 2744 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698175906
transform 1 0 6328 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_112
timestamp 1698175906
transform 1 0 6944 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_128
timestamp 1698175906
transform 1 0 7840 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_132
timestamp 1698175906
transform 1 0 8064 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_134
timestamp 1698175906
transform 1 0 8176 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_142
timestamp 1698175906
transform 1 0 8624 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_146
timestamp 1698175906
transform 1 0 8848 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_153
timestamp 1698175906
transform 1 0 9240 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_168
timestamp 1698175906
transform 1 0 10080 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_172
timestamp 1698175906
transform 1 0 10304 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_174
timestamp 1698175906
transform 1 0 10416 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_177
timestamp 1698175906
transform 1 0 10584 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_261
timestamp 1698175906
transform 1 0 15288 0 1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_293
timestamp 1698175906
transform 1 0 17080 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_309
timestamp 1698175906
transform 1 0 17976 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_313
timestamp 1698175906
transform 1 0 18200 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_317
timestamp 1698175906
transform 1 0 18424 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_321
timestamp 1698175906
transform 1 0 18648 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_28
timestamp 1698175906
transform 1 0 2240 0 -1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_60
timestamp 1698175906
transform 1 0 4032 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_68
timestamp 1698175906
transform 1 0 4480 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_72
timestamp 1698175906
transform 1 0 4704 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_76
timestamp 1698175906
transform 1 0 4928 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_78
timestamp 1698175906
transform 1 0 5040 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_116
timestamp 1698175906
transform 1 0 7168 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_120
timestamp 1698175906
transform 1 0 7392 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_124
timestamp 1698175906
transform 1 0 7616 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_126
timestamp 1698175906
transform 1 0 7728 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_134
timestamp 1698175906
transform 1 0 8176 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_155
timestamp 1698175906
transform 1 0 9352 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_157
timestamp 1698175906
transform 1 0 9464 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_169
timestamp 1698175906
transform 1 0 10136 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_175
timestamp 1698175906
transform 1 0 10472 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_196
timestamp 1698175906
transform 1 0 11648 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_206
timestamp 1698175906
transform 1 0 12208 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_212
timestamp 1698175906
transform 1 0 12544 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_220
timestamp 1698175906
transform 1 0 12992 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_224
timestamp 1698175906
transform 1 0 13216 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_254
timestamp 1698175906
transform 1 0 14896 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_258
timestamp 1698175906
transform 1 0 15120 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_274
timestamp 1698175906
transform 1 0 16016 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_278
timestamp 1698175906
transform 1 0 16240 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_282
timestamp 1698175906
transform 1 0 16464 0 -1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_314
timestamp 1698175906
transform 1 0 18256 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_322
timestamp 1698175906
transform 1 0 18704 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 784 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 2576 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_37
timestamp 1698175906
transform 1 0 2744 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_69
timestamp 1698175906
transform 1 0 4536 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_85
timestamp 1698175906
transform 1 0 5432 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_93
timestamp 1698175906
transform 1 0 5880 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698175906
transform 1 0 6328 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_112
timestamp 1698175906
transform 1 0 6944 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_116
timestamp 1698175906
transform 1 0 7168 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_118
timestamp 1698175906
transform 1 0 7280 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_183
timestamp 1698175906
transform 1 0 10920 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_185
timestamp 1698175906
transform 1 0 11032 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_203
timestamp 1698175906
transform 1 0 12040 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_211
timestamp 1698175906
transform 1 0 12488 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_224
timestamp 1698175906
transform 1 0 13216 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_228
timestamp 1698175906
transform 1 0 13440 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_243
timestamp 1698175906
transform 1 0 14280 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698175906
transform 1 0 14504 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698175906
transform 1 0 18088 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_317
timestamp 1698175906
transform 1 0 18424 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_321
timestamp 1698175906
transform 1 0 18648 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698175906
transform 1 0 784 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698175906
transform 1 0 4368 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_72
timestamp 1698175906
transform 1 0 4704 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_80
timestamp 1698175906
transform 1 0 5152 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_111
timestamp 1698175906
transform 1 0 6888 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_132
timestamp 1698175906
transform 1 0 8064 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_153
timestamp 1698175906
transform 1 0 9240 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_157
timestamp 1698175906
transform 1 0 9464 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_212
timestamp 1698175906
transform 1 0 12544 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_220
timestamp 1698175906
transform 1 0 12992 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_224
timestamp 1698175906
transform 1 0 13216 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_240
timestamp 1698175906
transform 1 0 14112 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_272
timestamp 1698175906
transform 1 0 15904 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_282
timestamp 1698175906
transform 1 0 16464 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_346
timestamp 1698175906
transform 1 0 20048 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_348
timestamp 1698175906
transform 1 0 20160 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_28
timestamp 1698175906
transform 1 0 2240 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_32
timestamp 1698175906
transform 1 0 2464 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 2576 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698175906
transform 1 0 2744 0 1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698175906
transform 1 0 6328 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_107
timestamp 1698175906
transform 1 0 6664 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_123
timestamp 1698175906
transform 1 0 7560 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_125
timestamp 1698175906
transform 1 0 7672 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_138
timestamp 1698175906
transform 1 0 8400 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_146
timestamp 1698175906
transform 1 0 8848 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_164
timestamp 1698175906
transform 1 0 9856 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_166
timestamp 1698175906
transform 1 0 9968 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_173
timestamp 1698175906
transform 1 0 10360 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_177
timestamp 1698175906
transform 1 0 10584 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_194
timestamp 1698175906
transform 1 0 11536 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698175906
transform 1 0 14504 0 1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698175906
transform 1 0 18088 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_317
timestamp 1698175906
transform 1 0 18424 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698175906
transform 1 0 784 0 -1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698175906
transform 1 0 4368 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_72
timestamp 1698175906
transform 1 0 4704 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_88
timestamp 1698175906
transform 1 0 5600 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_118
timestamp 1698175906
transform 1 0 7280 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_122
timestamp 1698175906
transform 1 0 7504 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_188
timestamp 1698175906
transform 1 0 11200 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_199
timestamp 1698175906
transform 1 0 11816 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_207
timestamp 1698175906
transform 1 0 12264 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_209
timestamp 1698175906
transform 1 0 12376 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_212
timestamp 1698175906
transform 1 0 12544 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_216
timestamp 1698175906
transform 1 0 12768 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_247
timestamp 1698175906
transform 1 0 14504 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_251
timestamp 1698175906
transform 1 0 14728 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_267
timestamp 1698175906
transform 1 0 15624 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_275
timestamp 1698175906
transform 1 0 16072 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_279
timestamp 1698175906
transform 1 0 16296 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698175906
transform 1 0 16464 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_314
timestamp 1698175906
transform 1 0 18256 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_322
timestamp 1698175906
transform 1 0 18704 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698175906
transform 1 0 784 0 1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 2576 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698175906
transform 1 0 2744 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698175906
transform 1 0 6328 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_107
timestamp 1698175906
transform 1 0 6664 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_115
timestamp 1698175906
transform 1 0 7112 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_119
timestamp 1698175906
transform 1 0 7336 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_148
timestamp 1698175906
transform 1 0 8960 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_160
timestamp 1698175906
transform 1 0 9632 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_164
timestamp 1698175906
transform 1 0 9856 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_202
timestamp 1698175906
transform 1 0 11984 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_210
timestamp 1698175906
transform 1 0 12432 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_214
timestamp 1698175906
transform 1 0 12656 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_247
timestamp 1698175906
transform 1 0 14504 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_251
timestamp 1698175906
transform 1 0 14728 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_317
timestamp 1698175906
transform 1 0 18424 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698175906
transform 1 0 18648 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2
timestamp 1698175906
transform 1 0 784 0 -1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_66
timestamp 1698175906
transform 1 0 4368 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_72
timestamp 1698175906
transform 1 0 4704 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_88
timestamp 1698175906
transform 1 0 5600 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_90
timestamp 1698175906
transform 1 0 5712 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_120
timestamp 1698175906
transform 1 0 7392 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_124
timestamp 1698175906
transform 1 0 7616 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_152
timestamp 1698175906
transform 1 0 9184 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_160
timestamp 1698175906
transform 1 0 9632 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_164
timestamp 1698175906
transform 1 0 9856 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_166
timestamp 1698175906
transform 1 0 9968 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_212
timestamp 1698175906
transform 1 0 12544 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_216
timestamp 1698175906
transform 1 0 12768 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_229
timestamp 1698175906
transform 1 0 13496 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_241
timestamp 1698175906
transform 1 0 14168 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_273
timestamp 1698175906
transform 1 0 15960 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_277
timestamp 1698175906
transform 1 0 16184 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_279
timestamp 1698175906
transform 1 0 16296 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_282
timestamp 1698175906
transform 1 0 16464 0 -1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_346
timestamp 1698175906
transform 1 0 20048 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_348
timestamp 1698175906
transform 1 0 20160 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_2
timestamp 1698175906
transform 1 0 784 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 2576 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698175906
transform 1 0 2744 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698175906
transform 1 0 6328 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_107
timestamp 1698175906
transform 1 0 6664 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_123
timestamp 1698175906
transform 1 0 7560 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_131
timestamp 1698175906
transform 1 0 8008 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_163
timestamp 1698175906
transform 1 0 9800 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_171
timestamp 1698175906
transform 1 0 10248 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_185
timestamp 1698175906
transform 1 0 11032 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_217
timestamp 1698175906
transform 1 0 12824 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_233
timestamp 1698175906
transform 1 0 13720 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_241
timestamp 1698175906
transform 1 0 14168 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 14504 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 18088 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_317
timestamp 1698175906
transform 1 0 18424 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698175906
transform 1 0 784 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698175906
transform 1 0 4368 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_72
timestamp 1698175906
transform 1 0 4704 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_88
timestamp 1698175906
transform 1 0 5600 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_90
timestamp 1698175906
transform 1 0 5712 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_126
timestamp 1698175906
transform 1 0 7728 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_128
timestamp 1698175906
transform 1 0 7840 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_136
timestamp 1698175906
transform 1 0 8288 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_142
timestamp 1698175906
transform 1 0 8624 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_154
timestamp 1698175906
transform 1 0 9296 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_187
timestamp 1698175906
transform 1 0 11144 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_191
timestamp 1698175906
transform 1 0 11368 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_193
timestamp 1698175906
transform 1 0 11480 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_202
timestamp 1698175906
transform 1 0 11984 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_217
timestamp 1698175906
transform 1 0 12824 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_249
timestamp 1698175906
transform 1 0 14616 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_265
timestamp 1698175906
transform 1 0 15512 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_273
timestamp 1698175906
transform 1 0 15960 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_277
timestamp 1698175906
transform 1 0 16184 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_279
timestamp 1698175906
transform 1 0 16296 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_282
timestamp 1698175906
transform 1 0 16464 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_314
timestamp 1698175906
transform 1 0 18256 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_330
timestamp 1698175906
transform 1 0 19152 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_338
timestamp 1698175906
transform 1 0 19600 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_342
timestamp 1698175906
transform 1 0 19824 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_344
timestamp 1698175906
transform 1 0 19936 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698175906
transform 1 0 784 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 2576 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 2744 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 6328 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_107
timestamp 1698175906
transform 1 0 6664 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_123
timestamp 1698175906
transform 1 0 7560 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_125
timestamp 1698175906
transform 1 0 7672 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_160
timestamp 1698175906
transform 1 0 9632 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_164
timestamp 1698175906
transform 1 0 9856 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_168
timestamp 1698175906
transform 1 0 10080 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_185
timestamp 1698175906
transform 1 0 11032 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_189
timestamp 1698175906
transform 1 0 11256 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_191
timestamp 1698175906
transform 1 0 11368 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_221
timestamp 1698175906
transform 1 0 13048 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_225
timestamp 1698175906
transform 1 0 13272 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_232
timestamp 1698175906
transform 1 0 13664 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_240
timestamp 1698175906
transform 1 0 14112 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_244
timestamp 1698175906
transform 1 0 14336 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 14504 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 18088 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_317
timestamp 1698175906
transform 1 0 18424 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2
timestamp 1698175906
transform 1 0 784 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_66
timestamp 1698175906
transform 1 0 4368 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_72
timestamp 1698175906
transform 1 0 4704 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_104
timestamp 1698175906
transform 1 0 6496 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_120
timestamp 1698175906
transform 1 0 7392 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_128
timestamp 1698175906
transform 1 0 7840 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_135
timestamp 1698175906
transform 1 0 8232 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_139
timestamp 1698175906
transform 1 0 8456 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_142
timestamp 1698175906
transform 1 0 8624 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_150
timestamp 1698175906
transform 1 0 9072 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_152
timestamp 1698175906
transform 1 0 9184 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_159
timestamp 1698175906
transform 1 0 9576 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_161
timestamp 1698175906
transform 1 0 9688 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_196
timestamp 1698175906
transform 1 0 11648 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_200
timestamp 1698175906
transform 1 0 11872 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_204
timestamp 1698175906
transform 1 0 12096 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_243
timestamp 1698175906
transform 1 0 14280 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_247
timestamp 1698175906
transform 1 0 14504 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_279
timestamp 1698175906
transform 1 0 16296 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_282
timestamp 1698175906
transform 1 0 16464 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_314
timestamp 1698175906
transform 1 0 18256 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_322
timestamp 1698175906
transform 1 0 18704 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698175906
transform 1 0 784 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 2576 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 2744 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 6328 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_107
timestamp 1698175906
transform 1 0 6664 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_111
timestamp 1698175906
transform 1 0 6888 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_113
timestamp 1698175906
transform 1 0 7000 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_148
timestamp 1698175906
transform 1 0 8960 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_152
timestamp 1698175906
transform 1 0 9184 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_168
timestamp 1698175906
transform 1 0 10080 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_172
timestamp 1698175906
transform 1 0 10304 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_174
timestamp 1698175906
transform 1 0 10416 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_185
timestamp 1698175906
transform 1 0 11032 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_201
timestamp 1698175906
transform 1 0 11928 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_209
timestamp 1698175906
transform 1 0 12376 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_216
timestamp 1698175906
transform 1 0 12768 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_224
timestamp 1698175906
transform 1 0 13216 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_232
timestamp 1698175906
transform 1 0 13664 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_240
timestamp 1698175906
transform 1 0 14112 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_244
timestamp 1698175906
transform 1 0 14336 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 14504 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 18088 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_317
timestamp 1698175906
transform 1 0 18424 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_321
timestamp 1698175906
transform 1 0 18648 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 784 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 4368 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1698175906
transform 1 0 4704 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698175906
transform 1 0 8288 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_142
timestamp 1698175906
transform 1 0 8624 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_206
timestamp 1698175906
transform 1 0 12208 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698175906
transform 1 0 12544 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698175906
transform 1 0 16128 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_282
timestamp 1698175906
transform 1 0 16464 0 -1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_314
timestamp 1698175906
transform 1 0 18256 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_322
timestamp 1698175906
transform 1 0 18704 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 784 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 2576 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 2744 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 6328 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698175906
transform 1 0 6664 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698175906
transform 1 0 10248 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698175906
transform 1 0 10584 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698175906
transform 1 0 14168 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 14504 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 18088 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 18424 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 784 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 4368 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 4704 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 8288 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 8624 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 12208 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 12544 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 16128 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 16464 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 20048 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 20160 0 -1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 784 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 2576 0 1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 2744 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 6328 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 6664 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 10248 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 10584 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 14168 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 14504 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 18088 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 18424 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 784 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 4368 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 4704 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 8288 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 8624 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 12208 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 12544 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 16128 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 16464 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 20048 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 20160 0 -1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 784 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 2576 0 1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 2744 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 6328 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 6664 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 10248 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 10584 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 14168 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 14504 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 18088 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 18424 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 784 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 4368 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 4704 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 8288 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 8624 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 12208 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 12544 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 16128 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 16464 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 20048 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 20160 0 -1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 784 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 2576 0 1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 2744 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 6328 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 6664 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 10248 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 10584 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 14168 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 14504 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 18088 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 18424 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 784 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 4368 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 4704 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 8288 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 8624 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 12208 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 12544 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 16128 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 16464 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 20048 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 20160 0 -1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 784 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 2576 0 1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 2744 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 6328 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 6664 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 10248 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 10584 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 14168 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 14504 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 18088 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 18424 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 784 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 4368 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 4704 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 8288 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 8624 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 12208 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 12544 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 16128 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 16464 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 20048 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 20160 0 -1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 784 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 2576 0 1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 2744 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 6328 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698175906
transform 1 0 6664 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698175906
transform 1 0 10248 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698175906
transform 1 0 10584 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 14168 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 14504 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 18088 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 18424 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 784 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 4368 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 4704 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 8288 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_168
timestamp 1698175906
transform 1 0 10080 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_176
timestamp 1698175906
transform 1 0 10528 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_180
timestamp 1698175906
transform 1 0 10752 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_207
timestamp 1698175906
transform 1 0 12264 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 12376 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_212
timestamp 1698175906
transform 1 0 12544 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_276
timestamp 1698175906
transform 1 0 16128 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 16464 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 20048 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 20160 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 784 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 2688 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 4592 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 6496 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_138
timestamp 1698175906
transform 1 0 8400 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_142
timestamp 1698175906
transform 1 0 8624 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_172
timestamp 1698175906
transform 1 0 10304 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_176
timestamp 1698175906
transform 1 0 10528 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_206
timestamp 1698175906
transform 1 0 12208 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_210
timestamp 1698175906
transform 1 0 12432 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_240
timestamp 1698175906
transform 1 0 14112 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 16016 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 17920 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 19824 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 20048 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 20160 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita38_25 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 15400 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita38_26
timestamp 1698175906
transform 1 0 19992 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10472 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform 1 0 18760 0 -1 9408
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform 1 0 18760 0 -1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform -1 0 2240 0 -1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform 1 0 18760 0 1 7056
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform 1 0 18760 0 -1 14112
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform 1 0 18760 0 -1 7840
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform 1 0 18760 0 -1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform -1 0 2240 0 1 10192
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform 1 0 18760 0 1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform 1 0 18760 0 1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform 1 0 18760 0 1 9408
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform 1 0 18760 0 1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform 1 0 12208 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform -1 0 12096 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform 1 0 8624 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform 1 0 8624 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform -1 0 2240 0 -1 9408
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform 1 0 10808 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform 1 0 8736 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform 1 0 8120 0 1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform 1 0 12544 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform -1 0 12096 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698175906
transform -1 0 10192 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 20328 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 20328 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 20328 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 20328 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 20328 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 20328 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 20328 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 672 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 20328 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 672 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 20328 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 672 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 20328 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 672 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 20328 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 672 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 20328 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 672 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 20328 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 672 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 20328 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 672 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 20328 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 672 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 20328 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 672 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 20328 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 672 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 20328 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 672 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 20328 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 672 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 20328 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 672 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 20328 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 672 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 20328 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 672 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 20328 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 672 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 20328 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 672 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 20328 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 672 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 20328 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 672 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 20328 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 672 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 20328 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 672 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 20328 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 672 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 20328 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 672 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 20328 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 672 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 20328 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 672 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 20328 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 672 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 20328 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 672 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 20328 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 672 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 20328 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 672 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 20328 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 672 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 20328 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 672 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 20328 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 672 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 20328 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 672 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 20328 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 672 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 20328 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 672 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 20328 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 672 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 20328 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 672 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 20328 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 2576 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 4480 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 6384 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 8288 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 10192 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 12096 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 14000 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 15904 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 17808 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 19712 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 4592 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 8512 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 12432 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 16352 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 6552 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 10472 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 14392 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 18312 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 4592 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 8512 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 12432 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 16352 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 6552 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 10472 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 14392 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 18312 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 4592 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 8512 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 12432 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 16352 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 6552 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 10472 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 14392 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 18312 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 4592 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 8512 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 12432 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 16352 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 2632 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 6552 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 10472 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 14392 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 18312 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 4592 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 8512 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 12432 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 16352 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 2632 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 6552 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 10472 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 14392 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 18312 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 4592 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 8512 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 12432 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 16352 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 2632 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 6552 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 10472 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 14392 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 18312 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 4592 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 8512 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 12432 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 16352 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 2632 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 6552 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 10472 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 14392 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 18312 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 4592 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 8512 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 12432 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 16352 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 2632 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 6552 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 10472 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 14392 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 18312 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 4592 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 8512 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 12432 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 16352 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 2632 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 6552 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 10472 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 14392 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 18312 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 4592 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 8512 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 12432 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 16352 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 2632 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 6552 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 10472 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 14392 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 18312 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 4592 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 8512 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 12432 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 16352 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 2632 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 6552 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 10472 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 14392 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 18312 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 4592 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 8512 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 12432 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 16352 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 2632 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 6552 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 10472 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 14392 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 18312 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 4592 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 8512 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 12432 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 16352 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 2632 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 6552 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 10472 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 14392 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 18312 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 4592 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 8512 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 12432 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 16352 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 2632 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 6552 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 10472 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 14392 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 18312 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 4592 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 8512 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 12432 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 16352 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 2632 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 6552 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 10472 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 14392 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 18312 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 4592 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 8512 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 12432 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 16352 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 2632 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 6552 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 10472 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 14392 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 18312 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 4592 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 8512 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 12432 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 16352 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 2632 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 6552 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 10472 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 14392 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 18312 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 4592 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 8512 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 12432 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 16352 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 2632 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 6552 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 10472 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 14392 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 18312 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 4592 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 8512 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 12432 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 16352 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 2632 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 6552 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 10472 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 14392 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 18312 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 4592 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 8512 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 12432 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 16352 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 2632 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 6552 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 10472 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 14392 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 18312 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 4592 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 8512 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 12432 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 16352 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 2632 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 6552 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 10472 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 14392 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 18312 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 4592 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 8512 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 12432 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 16352 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 2576 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 4480 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 6384 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 8288 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 10192 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 12096 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 14000 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 15904 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 17808 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 19712 0 1 18816
box -43 -43 155 435
<< labels >>
flabel metal3 s 0 13440 400 13496 0 FreeSans 224 0 0 0 clk
port 0 nsew signal input
flabel metal2 s 15120 0 15176 400 0 FreeSans 224 90 0 0 segm[0]
port 1 nsew signal tristate
flabel metal2 s 10416 0 10472 400 0 FreeSans 224 90 0 0 segm[10]
port 2 nsew signal tristate
flabel metal3 s 20600 9072 21000 9128 0 FreeSans 224 0 0 0 segm[11]
port 3 nsew signal tristate
flabel metal3 s 20600 10752 21000 10808 0 FreeSans 224 0 0 0 segm[12]
port 4 nsew signal tristate
flabel metal3 s 0 8064 400 8120 0 FreeSans 224 0 0 0 segm[13]
port 5 nsew signal tristate
flabel metal3 s 20600 7056 21000 7112 0 FreeSans 224 0 0 0 segm[1]
port 6 nsew signal tristate
flabel metal3 s 20600 12096 21000 12152 0 FreeSans 224 0 0 0 segm[2]
port 7 nsew signal tristate
flabel metal3 s 20600 13440 21000 13496 0 FreeSans 224 0 0 0 segm[3]
port 8 nsew signal tristate
flabel metal3 s 20600 7392 21000 7448 0 FreeSans 224 0 0 0 segm[4]
port 9 nsew signal tristate
flabel metal3 s 20600 12768 21000 12824 0 FreeSans 224 0 0 0 segm[5]
port 10 nsew signal tristate
flabel metal3 s 0 10080 400 10136 0 FreeSans 224 0 0 0 segm[6]
port 11 nsew signal tristate
flabel metal3 s 20600 11088 21000 11144 0 FreeSans 224 0 0 0 segm[7]
port 12 nsew signal tristate
flabel metal3 s 20600 8736 21000 8792 0 FreeSans 224 0 0 0 segm[8]
port 13 nsew signal tristate
flabel metal3 s 20600 9408 21000 9464 0 FreeSans 224 0 0 0 segm[9]
port 14 nsew signal tristate
flabel metal3 s 20600 13104 21000 13160 0 FreeSans 224 0 0 0 sel[0]
port 15 nsew signal tristate
flabel metal2 s 11760 0 11816 400 0 FreeSans 224 90 0 0 sel[10]
port 16 nsew signal tristate
flabel metal2 s 11088 0 11144 400 0 FreeSans 224 90 0 0 sel[11]
port 17 nsew signal tristate
flabel metal2 s 8400 0 8456 400 0 FreeSans 224 90 0 0 sel[1]
port 18 nsew signal tristate
flabel metal2 s 8400 20600 8456 21000 0 FreeSans 224 90 0 0 sel[2]
port 19 nsew signal tristate
flabel metal3 s 0 9072 400 9128 0 FreeSans 224 0 0 0 sel[3]
port 20 nsew signal tristate
flabel metal2 s 10752 20600 10808 21000 0 FreeSans 224 90 0 0 sel[4]
port 21 nsew signal tristate
flabel metal2 s 9744 0 9800 400 0 FreeSans 224 90 0 0 sel[5]
port 22 nsew signal tristate
flabel metal2 s 8064 0 8120 400 0 FreeSans 224 90 0 0 sel[6]
port 23 nsew signal tristate
flabel metal2 s 12768 20600 12824 21000 0 FreeSans 224 90 0 0 sel[7]
port 24 nsew signal tristate
flabel metal2 s 11088 20600 11144 21000 0 FreeSans 224 90 0 0 sel[8]
port 25 nsew signal tristate
flabel metal2 s 9072 20600 9128 21000 0 FreeSans 224 90 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 2224 1538 2384 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 17584 1538 17744 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 9904 1538 10064 19238 0 FreeSans 640 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 10500 19208 10500 19208 0 vdd
rlabel metal1 10500 18816 10500 18816 0 vss
rlabel metal2 8764 12488 8764 12488 0 _000_
rlabel metal2 10724 13300 10724 13300 0 _001_
rlabel metal2 11676 12572 11676 12572 0 _002_
rlabel metal2 9156 12152 9156 12152 0 _003_
rlabel metal2 6244 12040 6244 12040 0 _004_
rlabel metal2 6804 9744 6804 9744 0 _005_
rlabel metal2 11564 11368 11564 11368 0 _006_
rlabel metal2 7812 8232 7812 8232 0 _007_
rlabel metal2 8680 6524 8680 6524 0 _008_
rlabel metal2 9996 12432 9996 12432 0 _009_
rlabel metal3 6552 9212 6552 9212 0 _010_
rlabel metal2 7532 13300 7532 13300 0 _011_
rlabel metal2 7364 7056 7364 7056 0 _012_
rlabel metal2 12796 12544 12796 12544 0 _013_
rlabel metal2 9660 7700 9660 7700 0 _014_
rlabel metal2 6580 8092 6580 8092 0 _015_
rlabel metal2 11732 7434 11732 7434 0 _016_
rlabel metal2 10556 6944 10556 6944 0 _017_
rlabel metal2 13216 6916 13216 6916 0 _018_
rlabel metal2 6188 9828 6188 9828 0 _019_
rlabel metal2 13216 11228 13216 11228 0 _020_
rlabel metal2 14840 8484 14840 8484 0 _021_
rlabel metal2 11956 9016 11956 9016 0 _022_
rlabel metal2 13720 9268 13720 9268 0 _023_
rlabel metal2 13356 11172 13356 11172 0 _024_
rlabel metal2 11480 9492 11480 9492 0 _025_
rlabel metal2 6804 9072 6804 9072 0 _026_
rlabel metal3 8400 13468 8400 13468 0 _027_
rlabel metal2 8036 12712 8036 12712 0 _028_
rlabel metal2 8428 7280 8428 7280 0 _029_
rlabel metal3 8540 9324 8540 9324 0 _030_
rlabel metal3 11452 10864 11452 10864 0 _031_
rlabel metal2 12740 13160 12740 13160 0 _032_
rlabel metal3 9436 8540 9436 8540 0 _033_
rlabel metal2 9660 8708 9660 8708 0 _034_
rlabel metal3 11676 9212 11676 9212 0 _035_
rlabel metal3 10360 8092 10360 8092 0 _036_
rlabel metal2 7364 8624 7364 8624 0 _037_
rlabel metal3 7140 8428 7140 8428 0 _038_
rlabel metal2 12012 8260 12012 8260 0 _039_
rlabel metal2 11508 7952 11508 7952 0 _040_
rlabel metal2 13636 7896 13636 7896 0 _041_
rlabel metal2 11592 7644 11592 7644 0 _042_
rlabel metal2 8036 11144 8036 11144 0 _043_
rlabel metal2 13804 9100 13804 9100 0 _044_
rlabel metal3 8932 9660 8932 9660 0 _045_
rlabel metal3 10668 7196 10668 7196 0 _046_
rlabel metal2 14000 10052 14000 10052 0 _047_
rlabel metal2 14084 8960 14084 8960 0 _048_
rlabel metal2 13496 7756 13496 7756 0 _049_
rlabel metal2 13384 7364 13384 7364 0 _050_
rlabel metal2 7672 10052 7672 10052 0 _051_
rlabel metal3 6720 9660 6720 9660 0 _052_
rlabel metal3 13468 11564 13468 11564 0 _053_
rlabel metal2 12908 11648 12908 11648 0 _054_
rlabel metal3 14476 8820 14476 8820 0 _055_
rlabel metal2 15148 8792 15148 8792 0 _056_
rlabel metal2 11788 9352 11788 9352 0 _057_
rlabel metal2 12124 9352 12124 9352 0 _058_
rlabel metal2 13636 9408 13636 9408 0 _059_
rlabel metal2 13972 9688 13972 9688 0 _060_
rlabel metal2 11508 10724 11508 10724 0 _061_
rlabel metal2 11732 11116 11732 11116 0 _062_
rlabel metal2 13804 10416 13804 10416 0 _063_
rlabel metal2 8764 11396 8764 11396 0 _064_
rlabel metal2 7364 10444 7364 10444 0 _065_
rlabel metal3 9660 11172 9660 11172 0 _066_
rlabel metal3 10668 7952 10668 7952 0 _067_
rlabel metal2 11480 9604 11480 9604 0 _068_
rlabel metal2 10752 10500 10752 10500 0 _069_
rlabel metal3 10500 11172 10500 11172 0 _070_
rlabel metal2 8988 11368 8988 11368 0 _071_
rlabel metal2 9212 12516 9212 12516 0 _072_
rlabel metal3 8708 10780 8708 10780 0 _073_
rlabel metal2 10836 10640 10836 10640 0 _074_
rlabel metal2 10752 13524 10752 13524 0 _075_
rlabel metal2 12572 13454 12572 13454 0 _076_
rlabel metal2 11200 13524 11200 13524 0 _077_
rlabel metal3 8540 10836 8540 10836 0 _078_
rlabel metal2 9268 9632 9268 9632 0 _079_
rlabel metal2 11340 10248 11340 10248 0 _080_
rlabel metal2 9464 11172 9464 11172 0 _081_
rlabel metal2 9856 8708 9856 8708 0 _082_
rlabel metal2 11116 8988 11116 8988 0 _083_
rlabel metal2 11620 12516 11620 12516 0 _084_
rlabel metal2 11956 12740 11956 12740 0 _085_
rlabel metal2 5908 12208 5908 12208 0 _086_
rlabel metal2 9800 10444 9800 10444 0 _087_
rlabel metal3 6888 8540 6888 8540 0 _088_
rlabel metal2 8764 10836 8764 10836 0 _089_
rlabel metal2 8708 11676 8708 11676 0 _090_
rlabel metal2 6888 9548 6888 9548 0 _091_
rlabel metal2 11172 9464 11172 9464 0 _092_
rlabel metal2 11508 10178 11508 10178 0 _093_
rlabel metal3 11032 10724 11032 10724 0 _094_
rlabel metal2 8064 8428 8064 8428 0 _095_
rlabel metal2 7980 9800 7980 9800 0 _096_
rlabel metal2 7868 7364 7868 7364 0 _097_
rlabel metal2 8652 9548 8652 9548 0 _098_
rlabel metal3 8428 7364 8428 7364 0 _099_
rlabel metal3 8960 7308 8960 7308 0 _100_
rlabel metal2 13748 10822 13748 10822 0 _101_
rlabel metal3 9156 7196 9156 7196 0 _102_
rlabel metal2 10528 12740 10528 12740 0 _103_
rlabel metal3 1239 13468 1239 13468 0 clk
rlabel metal2 11760 10052 11760 10052 0 clknet_0_clk
rlabel metal2 5908 11256 5908 11256 0 clknet_1_0__leaf_clk
rlabel metal2 14476 12964 14476 12964 0 clknet_1_1__leaf_clk
rlabel metal2 7756 12152 7756 12152 0 dut38.count\[0\]
rlabel metal2 7308 11340 7308 11340 0 dut38.count\[1\]
rlabel metal2 7196 10920 7196 10920 0 dut38.count\[2\]
rlabel metal2 8036 10612 8036 10612 0 dut38.count\[3\]
rlabel metal2 10556 3178 10556 3178 0 net1
rlabel metal2 14308 11200 14308 11200 0 net10
rlabel metal2 13692 8428 13692 8428 0 net11
rlabel metal3 15960 9576 15960 9576 0 net12
rlabel metal2 18956 13104 18956 13104 0 net13
rlabel metal3 12544 7308 12544 7308 0 net14
rlabel metal2 11620 6776 11620 6776 0 net15
rlabel metal2 8596 2156 8596 2156 0 net16
rlabel metal2 8708 13580 8708 13580 0 net17
rlabel metal3 3178 9212 3178 9212 0 net18
rlabel metal2 10948 16030 10948 16030 0 net19
rlabel metal2 14084 9352 14084 9352 0 net2
rlabel metal3 9268 6524 9268 6524 0 net20
rlabel metal2 8204 3374 8204 3374 0 net21
rlabel metal2 12852 17486 12852 17486 0 net22
rlabel metal2 11788 16226 11788 16226 0 net23
rlabel metal2 9660 19012 9660 19012 0 net24
rlabel metal2 15148 1015 15148 1015 0 net25
rlabel metal2 20132 12264 20132 12264 0 net26
rlabel metal3 14168 10724 14168 10724 0 net3
rlabel metal2 5516 8008 5516 8008 0 net4
rlabel metal3 18844 7196 18844 7196 0 net5
rlabel metal2 13580 13552 13580 13552 0 net6
rlabel metal2 13916 7224 13916 7224 0 net7
rlabel metal2 13468 12908 13468 12908 0 net8
rlabel metal3 3752 10388 3752 10388 0 net9
rlabel metal2 10444 1211 10444 1211 0 segm[10]
rlabel metal3 20321 9100 20321 9100 0 segm[11]
rlabel metal2 20020 10752 20020 10752 0 segm[12]
rlabel metal3 679 8092 679 8092 0 segm[13]
rlabel metal2 20020 7196 20020 7196 0 segm[1]
rlabel metal2 19964 13664 19964 13664 0 segm[3]
rlabel metal2 20020 7504 20020 7504 0 segm[4]
rlabel metal2 20020 12908 20020 12908 0 segm[5]
rlabel metal3 679 10108 679 10108 0 segm[6]
rlabel metal2 20020 11172 20020 11172 0 segm[7]
rlabel metal2 20020 8820 20020 8820 0 segm[8]
rlabel metal2 20020 9548 20020 9548 0 segm[9]
rlabel metal2 20020 13356 20020 13356 0 sel[0]
rlabel metal2 11788 1099 11788 1099 0 sel[10]
rlabel metal2 11116 1043 11116 1043 0 sel[11]
rlabel metal2 8428 1211 8428 1211 0 sel[1]
rlabel metal2 8428 19677 8428 19677 0 sel[2]
rlabel metal3 679 9100 679 9100 0 sel[3]
rlabel metal2 10780 19677 10780 19677 0 sel[4]
rlabel metal2 9772 1043 9772 1043 0 sel[5]
rlabel metal2 8092 1491 8092 1491 0 sel[6]
rlabel metal2 12796 20573 12796 20573 0 sel[7]
rlabel metal2 11116 19845 11116 19845 0 sel[8]
rlabel metal2 9100 19845 9100 19845 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 21000 21000
<< end >>
