magic
tech gf180mcuD
magscale 1 5
timestamp 1699641881
<< metal1 >>
rect 672 19221 20328 19238
rect 672 19195 2239 19221
rect 2265 19195 2291 19221
rect 2317 19195 2343 19221
rect 2369 19195 17599 19221
rect 17625 19195 17651 19221
rect 17677 19195 17703 19221
rect 17729 19195 20328 19221
rect 672 19178 20328 19195
rect 9311 19137 9337 19143
rect 9311 19105 9337 19111
rect 11215 19137 11241 19143
rect 11215 19105 11241 19111
rect 13063 19137 13089 19143
rect 13063 19105 13089 19111
rect 8801 18999 8807 19025
rect 8833 18999 8839 19025
rect 10817 18999 10823 19025
rect 10849 18999 10855 19025
rect 12665 18999 12671 19025
rect 12697 18999 12703 19025
rect 14239 18969 14265 18975
rect 14239 18937 14265 18943
rect 672 18829 20328 18846
rect 672 18803 9919 18829
rect 9945 18803 9971 18829
rect 9997 18803 10023 18829
rect 10049 18803 20328 18829
rect 672 18786 20328 18803
rect 9927 18745 9953 18751
rect 9927 18713 9953 18719
rect 11383 18745 11409 18751
rect 11383 18713 11409 18719
rect 13399 18745 13425 18751
rect 13399 18713 13425 18719
rect 9417 18607 9423 18633
rect 9449 18607 9455 18633
rect 11097 18607 11103 18633
rect 11129 18607 11135 18633
rect 12945 18607 12951 18633
rect 12977 18607 12983 18633
rect 672 18437 20328 18454
rect 672 18411 2239 18437
rect 2265 18411 2291 18437
rect 2317 18411 2343 18437
rect 2369 18411 17599 18437
rect 17625 18411 17651 18437
rect 17677 18411 17703 18437
rect 17729 18411 20328 18437
rect 672 18394 20328 18411
rect 9031 18353 9057 18359
rect 9031 18321 9057 18327
rect 8521 18215 8527 18241
rect 8553 18215 8559 18241
rect 672 18045 20328 18062
rect 672 18019 9919 18045
rect 9945 18019 9971 18045
rect 9997 18019 10023 18045
rect 10049 18019 20328 18045
rect 672 18002 20328 18019
rect 672 17653 20328 17670
rect 672 17627 2239 17653
rect 2265 17627 2291 17653
rect 2317 17627 2343 17653
rect 2369 17627 17599 17653
rect 17625 17627 17651 17653
rect 17677 17627 17703 17653
rect 17729 17627 20328 17653
rect 672 17610 20328 17627
rect 672 17261 20328 17278
rect 672 17235 9919 17261
rect 9945 17235 9971 17261
rect 9997 17235 10023 17261
rect 10049 17235 20328 17261
rect 672 17218 20328 17235
rect 672 16869 20328 16886
rect 672 16843 2239 16869
rect 2265 16843 2291 16869
rect 2317 16843 2343 16869
rect 2369 16843 17599 16869
rect 17625 16843 17651 16869
rect 17677 16843 17703 16869
rect 17729 16843 20328 16869
rect 672 16826 20328 16843
rect 672 16477 20328 16494
rect 672 16451 9919 16477
rect 9945 16451 9971 16477
rect 9997 16451 10023 16477
rect 10049 16451 20328 16477
rect 672 16434 20328 16451
rect 672 16085 20328 16102
rect 672 16059 2239 16085
rect 2265 16059 2291 16085
rect 2317 16059 2343 16085
rect 2369 16059 17599 16085
rect 17625 16059 17651 16085
rect 17677 16059 17703 16085
rect 17729 16059 20328 16085
rect 672 16042 20328 16059
rect 672 15693 20328 15710
rect 672 15667 9919 15693
rect 9945 15667 9971 15693
rect 9997 15667 10023 15693
rect 10049 15667 20328 15693
rect 672 15650 20328 15667
rect 672 15301 20328 15318
rect 672 15275 2239 15301
rect 2265 15275 2291 15301
rect 2317 15275 2343 15301
rect 2369 15275 17599 15301
rect 17625 15275 17651 15301
rect 17677 15275 17703 15301
rect 17729 15275 20328 15301
rect 672 15258 20328 15275
rect 672 14909 20328 14926
rect 672 14883 9919 14909
rect 9945 14883 9971 14909
rect 9997 14883 10023 14909
rect 10049 14883 20328 14909
rect 672 14866 20328 14883
rect 672 14517 20328 14534
rect 672 14491 2239 14517
rect 2265 14491 2291 14517
rect 2317 14491 2343 14517
rect 2369 14491 17599 14517
rect 17625 14491 17651 14517
rect 17677 14491 17703 14517
rect 17729 14491 20328 14517
rect 672 14474 20328 14491
rect 672 14125 20328 14142
rect 672 14099 9919 14125
rect 9945 14099 9971 14125
rect 9997 14099 10023 14125
rect 10049 14099 20328 14125
rect 672 14082 20328 14099
rect 8247 14041 8273 14047
rect 8247 14009 8273 14015
rect 12671 14041 12697 14047
rect 12671 14009 12697 14015
rect 8135 13929 8161 13935
rect 8135 13897 8161 13903
rect 8303 13929 8329 13935
rect 12615 13929 12641 13935
rect 9249 13903 9255 13929
rect 9281 13903 9287 13929
rect 10929 13903 10935 13929
rect 10961 13903 10967 13929
rect 8303 13897 8329 13903
rect 12615 13897 12641 13903
rect 13007 13929 13033 13935
rect 13007 13897 13033 13903
rect 8807 13873 8833 13879
rect 8807 13841 8833 13847
rect 9143 13873 9169 13879
rect 9641 13847 9647 13873
rect 9673 13847 9679 13873
rect 10705 13847 10711 13873
rect 10737 13847 10743 13873
rect 11265 13847 11271 13873
rect 11297 13847 11303 13873
rect 12329 13847 12335 13873
rect 12361 13847 12367 13873
rect 9143 13841 9169 13847
rect 12671 13817 12697 13823
rect 12671 13785 12697 13791
rect 672 13733 20328 13750
rect 672 13707 2239 13733
rect 2265 13707 2291 13733
rect 2317 13707 2343 13733
rect 2369 13707 17599 13733
rect 17625 13707 17651 13733
rect 17677 13707 17703 13733
rect 17729 13707 20328 13733
rect 672 13690 20328 13707
rect 10711 13593 10737 13599
rect 13175 13593 13201 13599
rect 8745 13567 8751 13593
rect 8777 13567 8783 13593
rect 10369 13567 10375 13593
rect 10401 13567 10407 13593
rect 12945 13567 12951 13593
rect 12977 13567 12983 13593
rect 10711 13561 10737 13567
rect 13175 13561 13201 13567
rect 11047 13537 11073 13543
rect 7289 13511 7295 13537
rect 7321 13511 7327 13537
rect 8969 13511 8975 13537
rect 9001 13511 9007 13537
rect 10929 13511 10935 13537
rect 10961 13511 10967 13537
rect 11489 13511 11495 13537
rect 11521 13511 11527 13537
rect 11047 13505 11073 13511
rect 10655 13481 10681 13487
rect 7681 13455 7687 13481
rect 7713 13455 7719 13481
rect 9305 13455 9311 13481
rect 9337 13455 9343 13481
rect 10655 13449 10681 13455
rect 10767 13481 10793 13487
rect 10767 13449 10793 13455
rect 11159 13481 11185 13487
rect 11159 13449 11185 13455
rect 11215 13481 11241 13487
rect 11881 13455 11887 13481
rect 11913 13455 11919 13481
rect 11215 13449 11241 13455
rect 672 13341 20328 13358
rect 672 13315 9919 13341
rect 9945 13315 9971 13341
rect 9997 13315 10023 13341
rect 10049 13315 20328 13341
rect 672 13298 20328 13315
rect 9087 13257 9113 13263
rect 10711 13257 10737 13263
rect 9641 13231 9647 13257
rect 9673 13231 9679 13257
rect 9087 13225 9113 13231
rect 10711 13225 10737 13231
rect 11719 13257 11745 13263
rect 11719 13225 11745 13231
rect 12223 13257 12249 13263
rect 12223 13225 12249 13231
rect 12559 13257 12585 13263
rect 12559 13225 12585 13231
rect 9143 13201 9169 13207
rect 11775 13201 11801 13207
rect 10873 13175 10879 13201
rect 10905 13175 10911 13201
rect 9143 13169 9169 13175
rect 11775 13169 11801 13175
rect 12167 13201 12193 13207
rect 12167 13169 12193 13175
rect 12335 13201 12361 13207
rect 12335 13169 12361 13175
rect 12671 13201 12697 13207
rect 12671 13169 12697 13175
rect 11663 13145 11689 13151
rect 6897 13119 6903 13145
rect 6929 13119 6935 13145
rect 9753 13119 9759 13145
rect 9785 13119 9791 13145
rect 11663 13113 11689 13119
rect 11999 13145 12025 13151
rect 11999 13113 12025 13119
rect 12727 13145 12753 13151
rect 12727 13113 12753 13119
rect 8863 13089 8889 13095
rect 7233 13063 7239 13089
rect 7265 13063 7271 13089
rect 8297 13063 8303 13089
rect 8329 13063 8335 13089
rect 8863 13057 8889 13063
rect 9087 13033 9113 13039
rect 9087 13001 9113 13007
rect 672 12949 20328 12966
rect 672 12923 2239 12949
rect 2265 12923 2291 12949
rect 2317 12923 2343 12949
rect 2369 12923 17599 12949
rect 17625 12923 17651 12949
rect 17677 12923 17703 12949
rect 17729 12923 20328 12949
rect 672 12906 20328 12923
rect 8807 12809 8833 12815
rect 8807 12777 8833 12783
rect 7631 12753 7657 12759
rect 7631 12721 7657 12727
rect 7799 12753 7825 12759
rect 7799 12721 7825 12727
rect 9087 12753 9113 12759
rect 9087 12721 9113 12727
rect 7743 12641 7769 12647
rect 7743 12609 7769 12615
rect 8415 12641 8441 12647
rect 8415 12609 8441 12615
rect 8751 12641 8777 12647
rect 8751 12609 8777 12615
rect 8863 12641 8889 12647
rect 8863 12609 8889 12615
rect 672 12557 20328 12574
rect 672 12531 9919 12557
rect 9945 12531 9971 12557
rect 9997 12531 10023 12557
rect 10049 12531 20328 12557
rect 672 12514 20328 12531
rect 12615 12361 12641 12367
rect 12615 12329 12641 12335
rect 12783 12361 12809 12367
rect 12783 12329 12809 12335
rect 12895 12361 12921 12367
rect 18937 12335 18943 12361
rect 18969 12335 18975 12361
rect 12895 12329 12921 12335
rect 12839 12305 12865 12311
rect 12839 12273 12865 12279
rect 20007 12249 20033 12255
rect 20007 12217 20033 12223
rect 672 12165 20328 12182
rect 672 12139 2239 12165
rect 2265 12139 2291 12165
rect 2317 12139 2343 12165
rect 2369 12139 17599 12165
rect 17625 12139 17651 12165
rect 17677 12139 17703 12165
rect 17729 12139 20328 12165
rect 672 12122 20328 12139
rect 9479 12081 9505 12087
rect 9479 12049 9505 12055
rect 967 12025 993 12031
rect 11327 12025 11353 12031
rect 9361 11999 9367 12025
rect 9393 11999 9399 12025
rect 11041 11999 11047 12025
rect 11073 11999 11079 12025
rect 967 11993 993 11999
rect 11327 11993 11353 11999
rect 11887 12025 11913 12031
rect 20007 12025 20033 12031
rect 13673 11999 13679 12025
rect 13705 11999 13711 12025
rect 11887 11993 11913 11999
rect 20007 11993 20033 11999
rect 9815 11969 9841 11975
rect 2137 11943 2143 11969
rect 2169 11943 2175 11969
rect 6785 11943 6791 11969
rect 6817 11943 6823 11969
rect 7961 11943 7967 11969
rect 7993 11943 7999 11969
rect 9815 11937 9841 11943
rect 9983 11969 10009 11975
rect 9983 11937 10009 11943
rect 10823 11969 10849 11975
rect 10823 11937 10849 11943
rect 10991 11969 11017 11975
rect 10991 11937 11017 11943
rect 11551 11969 11577 11975
rect 11551 11937 11577 11943
rect 11831 11969 11857 11975
rect 12217 11943 12223 11969
rect 12249 11943 12255 11969
rect 13897 11943 13903 11969
rect 13929 11943 13935 11969
rect 18825 11943 18831 11969
rect 18857 11943 18863 11969
rect 11831 11937 11857 11943
rect 8297 11887 8303 11913
rect 8329 11887 8335 11913
rect 12609 11887 12615 11913
rect 12641 11887 12647 11913
rect 6903 11857 6929 11863
rect 6903 11825 6929 11831
rect 9535 11857 9561 11863
rect 9535 11825 9561 11831
rect 9647 11857 9673 11863
rect 9647 11825 9673 11831
rect 10879 11857 10905 11863
rect 10879 11825 10905 11831
rect 11047 11857 11073 11863
rect 11047 11825 11073 11831
rect 11607 11857 11633 11863
rect 11607 11825 11633 11831
rect 11719 11857 11745 11863
rect 14239 11857 14265 11863
rect 14009 11831 14015 11857
rect 14041 11831 14047 11857
rect 11719 11825 11745 11831
rect 14239 11825 14265 11831
rect 672 11773 20328 11790
rect 672 11747 9919 11773
rect 9945 11747 9971 11773
rect 9997 11747 10023 11773
rect 10049 11747 20328 11773
rect 672 11730 20328 11747
rect 8135 11689 8161 11695
rect 8135 11657 8161 11663
rect 12055 11689 12081 11695
rect 12055 11657 12081 11663
rect 12111 11689 12137 11695
rect 12111 11657 12137 11663
rect 12167 11689 12193 11695
rect 12167 11657 12193 11663
rect 8023 11633 8049 11639
rect 7065 11607 7071 11633
rect 7097 11607 7103 11633
rect 8023 11601 8049 11607
rect 9143 11633 9169 11639
rect 9143 11601 9169 11607
rect 12279 11633 12305 11639
rect 13001 11607 13007 11633
rect 13033 11607 13039 11633
rect 12279 11601 12305 11607
rect 7631 11577 7657 11583
rect 7401 11551 7407 11577
rect 7433 11551 7439 11577
rect 7631 11545 7657 11551
rect 7743 11577 7769 11583
rect 7743 11545 7769 11551
rect 7967 11577 7993 11583
rect 7967 11545 7993 11551
rect 8191 11577 8217 11583
rect 8191 11545 8217 11551
rect 9031 11577 9057 11583
rect 9031 11545 9057 11551
rect 9367 11577 9393 11583
rect 11327 11577 11353 11583
rect 11209 11551 11215 11577
rect 11241 11551 11247 11577
rect 9367 11545 9393 11551
rect 11327 11545 11353 11551
rect 11551 11577 11577 11583
rect 11551 11545 11577 11551
rect 11663 11577 11689 11583
rect 12335 11577 12361 11583
rect 14295 11577 14321 11583
rect 11825 11551 11831 11577
rect 11857 11551 11863 11577
rect 11937 11551 11943 11577
rect 11969 11551 11975 11577
rect 12609 11551 12615 11577
rect 12641 11551 12647 11577
rect 18825 11551 18831 11577
rect 18857 11551 18863 11577
rect 11663 11545 11689 11551
rect 12335 11545 12361 11551
rect 14295 11545 14321 11551
rect 7687 11521 7713 11527
rect 11607 11521 11633 11527
rect 6001 11495 6007 11521
rect 6033 11495 6039 11521
rect 9753 11495 9759 11521
rect 9785 11495 9791 11521
rect 10817 11495 10823 11521
rect 10849 11495 10855 11521
rect 14065 11495 14071 11521
rect 14097 11495 14103 11521
rect 7687 11489 7713 11495
rect 11607 11489 11633 11495
rect 8975 11465 9001 11471
rect 8975 11433 9001 11439
rect 9255 11465 9281 11471
rect 9255 11433 9281 11439
rect 20007 11465 20033 11471
rect 20007 11433 20033 11439
rect 672 11381 20328 11398
rect 672 11355 2239 11381
rect 2265 11355 2291 11381
rect 2317 11355 2343 11381
rect 2369 11355 17599 11381
rect 17625 11355 17651 11381
rect 17677 11355 17703 11381
rect 17729 11355 20328 11381
rect 672 11338 20328 11355
rect 7239 11297 7265 11303
rect 7065 11271 7071 11297
rect 7097 11271 7103 11297
rect 7239 11265 7265 11271
rect 9031 11297 9057 11303
rect 9031 11265 9057 11271
rect 12391 11297 12417 11303
rect 12391 11265 12417 11271
rect 7799 11241 7825 11247
rect 7799 11209 7825 11215
rect 9255 11241 9281 11247
rect 9255 11209 9281 11215
rect 20007 11241 20033 11247
rect 20007 11209 20033 11215
rect 7351 11185 7377 11191
rect 7351 11153 7377 11159
rect 7967 11185 7993 11191
rect 7967 11153 7993 11159
rect 9143 11185 9169 11191
rect 9143 11153 9169 11159
rect 9311 11185 9337 11191
rect 9311 11153 9337 11159
rect 10655 11185 10681 11191
rect 10655 11153 10681 11159
rect 12279 11185 12305 11191
rect 12279 11153 12305 11159
rect 13119 11185 13145 11191
rect 18825 11159 18831 11185
rect 18857 11159 18863 11185
rect 13119 11153 13145 11159
rect 8079 11129 8105 11135
rect 8079 11097 8105 11103
rect 8975 11129 9001 11135
rect 8975 11097 9001 11103
rect 9479 11129 9505 11135
rect 9871 11129 9897 11135
rect 12559 11129 12585 11135
rect 9697 11103 9703 11129
rect 9729 11103 9735 11129
rect 10817 11103 10823 11129
rect 10849 11103 10855 11129
rect 11153 11103 11159 11129
rect 11185 11103 11191 11129
rect 9479 11097 9505 11103
rect 9871 11097 9897 11103
rect 12559 11097 12585 11103
rect 13231 11129 13257 11135
rect 13231 11097 13257 11103
rect 13287 11129 13313 11135
rect 13287 11097 13313 11103
rect 14239 11129 14265 11135
rect 14239 11097 14265 11103
rect 6903 11073 6929 11079
rect 6903 11041 6929 11047
rect 7575 11073 7601 11079
rect 12447 11073 12473 11079
rect 10873 11047 10879 11073
rect 10905 11047 10911 11073
rect 7575 11041 7601 11047
rect 12447 11041 12473 11047
rect 14071 11073 14097 11079
rect 14071 11041 14097 11047
rect 14743 11073 14769 11079
rect 14905 11047 14911 11073
rect 14937 11047 14943 11073
rect 14743 11041 14769 11047
rect 672 10989 20328 11006
rect 672 10963 9919 10989
rect 9945 10963 9971 10989
rect 9997 10963 10023 10989
rect 10049 10963 20328 10989
rect 672 10946 20328 10963
rect 8023 10905 8049 10911
rect 11663 10905 11689 10911
rect 9473 10879 9479 10905
rect 9505 10879 9511 10905
rect 8023 10873 8049 10879
rect 11663 10873 11689 10879
rect 13175 10905 13201 10911
rect 13175 10873 13201 10879
rect 9927 10849 9953 10855
rect 10599 10849 10625 10855
rect 10425 10823 10431 10849
rect 10457 10823 10463 10849
rect 13337 10823 13343 10849
rect 13369 10823 13375 10849
rect 14065 10823 14071 10849
rect 14097 10823 14103 10849
rect 9927 10817 9953 10823
rect 10599 10817 10625 10823
rect 7855 10793 7881 10799
rect 5609 10767 5615 10793
rect 5641 10767 5647 10793
rect 7457 10767 7463 10793
rect 7489 10767 7495 10793
rect 7855 10761 7881 10767
rect 9311 10793 9337 10799
rect 11439 10793 11465 10799
rect 10201 10767 10207 10793
rect 10233 10767 10239 10793
rect 10705 10767 10711 10793
rect 10737 10767 10743 10793
rect 9311 10761 9337 10767
rect 11439 10761 11465 10767
rect 11719 10793 11745 10799
rect 11719 10761 11745 10767
rect 11775 10793 11801 10799
rect 11775 10761 11801 10767
rect 11887 10793 11913 10799
rect 11887 10761 11913 10767
rect 12111 10793 12137 10799
rect 12111 10761 12137 10767
rect 12167 10793 12193 10799
rect 13449 10767 13455 10793
rect 13481 10767 13487 10793
rect 13673 10767 13679 10793
rect 13705 10767 13711 10793
rect 18825 10767 18831 10793
rect 18857 10767 18863 10793
rect 12167 10761 12193 10767
rect 7183 10737 7209 10743
rect 9647 10737 9673 10743
rect 5945 10711 5951 10737
rect 5977 10711 5983 10737
rect 7009 10711 7015 10737
rect 7041 10711 7047 10737
rect 7569 10711 7575 10737
rect 7601 10711 7607 10737
rect 7183 10705 7209 10711
rect 9647 10705 9673 10711
rect 11999 10737 12025 10743
rect 20007 10737 20033 10743
rect 15129 10711 15135 10737
rect 15161 10711 15167 10737
rect 11999 10705 12025 10711
rect 20007 10705 20033 10711
rect 10375 10681 10401 10687
rect 10375 10649 10401 10655
rect 672 10597 20328 10614
rect 672 10571 2239 10597
rect 2265 10571 2291 10597
rect 2317 10571 2343 10597
rect 2369 10571 17599 10597
rect 17625 10571 17651 10597
rect 17677 10571 17703 10597
rect 17729 10571 20328 10597
rect 672 10554 20328 10571
rect 14575 10513 14601 10519
rect 14575 10481 14601 10487
rect 11271 10457 11297 10463
rect 14743 10457 14769 10463
rect 7513 10431 7519 10457
rect 7545 10431 7551 10457
rect 7905 10431 7911 10457
rect 7937 10431 7943 10457
rect 10873 10431 10879 10457
rect 10905 10431 10911 10457
rect 13169 10431 13175 10457
rect 13201 10431 13207 10457
rect 15017 10431 15023 10457
rect 15049 10431 15055 10457
rect 11271 10425 11297 10431
rect 14743 10425 14769 10431
rect 6399 10401 6425 10407
rect 15191 10401 15217 10407
rect 7009 10375 7015 10401
rect 7041 10375 7047 10401
rect 7345 10375 7351 10401
rect 7377 10375 7383 10401
rect 10033 10375 10039 10401
rect 10065 10375 10071 10401
rect 10649 10375 10655 10401
rect 10681 10375 10687 10401
rect 11657 10375 11663 10401
rect 11689 10375 11695 10401
rect 6399 10369 6425 10375
rect 15191 10369 15217 10375
rect 15303 10401 15329 10407
rect 15303 10369 15329 10375
rect 6231 10345 6257 10351
rect 6231 10313 6257 10319
rect 11047 10345 11073 10351
rect 11047 10313 11073 10319
rect 11159 10345 11185 10351
rect 11159 10313 11185 10319
rect 11327 10345 11353 10351
rect 11327 10313 11353 10319
rect 14855 10345 14881 10351
rect 14855 10313 14881 10319
rect 10767 10289 10793 10295
rect 7121 10263 7127 10289
rect 7153 10263 7159 10289
rect 10767 10257 10793 10263
rect 10879 10289 10905 10295
rect 10879 10257 10905 10263
rect 672 10205 20328 10222
rect 672 10179 9919 10205
rect 9945 10179 9971 10205
rect 9997 10179 10023 10205
rect 10049 10179 20328 10205
rect 672 10162 20328 10179
rect 12559 10121 12585 10127
rect 9361 10095 9367 10121
rect 9393 10095 9399 10121
rect 12559 10089 12585 10095
rect 8359 10065 8385 10071
rect 9535 10065 9561 10071
rect 12671 10065 12697 10071
rect 8689 10039 8695 10065
rect 8721 10039 8727 10065
rect 9417 10039 9423 10065
rect 9449 10039 9455 10065
rect 11657 10039 11663 10065
rect 11689 10039 11695 10065
rect 8359 10033 8385 10039
rect 9535 10033 9561 10039
rect 12671 10033 12697 10039
rect 15023 10065 15049 10071
rect 15023 10033 15049 10039
rect 12727 10009 12753 10015
rect 8073 9983 8079 10009
rect 8105 9983 8111 10009
rect 8801 9983 8807 10009
rect 8833 9983 8839 10009
rect 9193 9983 9199 10009
rect 9225 9983 9231 10009
rect 9697 9983 9703 10009
rect 9729 9983 9735 10009
rect 13337 9983 13343 10009
rect 13369 9983 13375 10009
rect 18825 9983 18831 10009
rect 18857 9983 18863 10009
rect 12727 9977 12753 9983
rect 8017 9927 8023 9953
rect 8049 9927 8055 9953
rect 13729 9927 13735 9953
rect 13761 9927 13767 9953
rect 14793 9927 14799 9953
rect 14825 9927 14831 9953
rect 9311 9897 9337 9903
rect 9311 9865 9337 9871
rect 20007 9897 20033 9903
rect 20007 9865 20033 9871
rect 672 9813 20328 9830
rect 672 9787 2239 9813
rect 2265 9787 2291 9813
rect 2317 9787 2343 9813
rect 2369 9787 17599 9813
rect 17625 9787 17651 9813
rect 17677 9787 17703 9813
rect 17729 9787 20328 9813
rect 672 9770 20328 9787
rect 9143 9673 9169 9679
rect 8801 9647 8807 9673
rect 8833 9647 8839 9673
rect 9143 9641 9169 9647
rect 9423 9673 9449 9679
rect 9423 9641 9449 9647
rect 10655 9673 10681 9679
rect 12559 9673 12585 9679
rect 11265 9647 11271 9673
rect 11297 9647 11303 9673
rect 12329 9647 12335 9673
rect 12361 9647 12367 9673
rect 10655 9641 10681 9647
rect 12559 9641 12585 9647
rect 13623 9673 13649 9679
rect 13623 9641 13649 9647
rect 20007 9673 20033 9679
rect 20007 9641 20033 9647
rect 8975 9617 9001 9623
rect 13511 9617 13537 9623
rect 8465 9591 8471 9617
rect 8497 9591 8503 9617
rect 9641 9591 9647 9617
rect 9673 9591 9679 9617
rect 9809 9591 9815 9617
rect 9841 9591 9847 9617
rect 10145 9591 10151 9617
rect 10177 9591 10183 9617
rect 10929 9591 10935 9617
rect 10961 9591 10967 9617
rect 8975 9585 9001 9591
rect 13511 9585 13537 9591
rect 13735 9617 13761 9623
rect 13735 9585 13761 9591
rect 14071 9617 14097 9623
rect 14071 9585 14097 9591
rect 14239 9617 14265 9623
rect 18825 9591 18831 9617
rect 18857 9591 18863 9617
rect 14239 9585 14265 9591
rect 8023 9561 8049 9567
rect 8023 9529 8049 9535
rect 8191 9561 8217 9567
rect 8191 9529 8217 9535
rect 9479 9561 9505 9567
rect 13231 9561 13257 9567
rect 10257 9535 10263 9561
rect 10289 9535 10295 9561
rect 9479 9529 9505 9535
rect 13231 9529 13257 9535
rect 13847 9561 13873 9567
rect 13847 9529 13873 9535
rect 14183 9561 14209 9567
rect 14183 9529 14209 9535
rect 8583 9505 8609 9511
rect 8583 9473 8609 9479
rect 10711 9505 10737 9511
rect 10711 9473 10737 9479
rect 13287 9505 13313 9511
rect 13287 9473 13313 9479
rect 13399 9505 13425 9511
rect 13399 9473 13425 9479
rect 672 9421 20328 9438
rect 672 9395 9919 9421
rect 9945 9395 9971 9421
rect 9997 9395 10023 9421
rect 10049 9395 20328 9421
rect 672 9378 20328 9395
rect 10823 9337 10849 9343
rect 9081 9311 9087 9337
rect 9113 9311 9119 9337
rect 10823 9305 10849 9311
rect 10935 9337 10961 9343
rect 11209 9311 11215 9337
rect 11241 9311 11247 9337
rect 11713 9311 11719 9337
rect 11745 9311 11751 9337
rect 10935 9305 10961 9311
rect 7855 9281 7881 9287
rect 7855 9249 7881 9255
rect 7911 9281 7937 9287
rect 7911 9249 7937 9255
rect 9703 9281 9729 9287
rect 9703 9249 9729 9255
rect 10039 9281 10065 9287
rect 10039 9249 10065 9255
rect 10711 9281 10737 9287
rect 10711 9249 10737 9255
rect 7743 9225 7769 9231
rect 6225 9199 6231 9225
rect 6257 9199 6263 9225
rect 6561 9199 6567 9225
rect 6593 9199 6599 9225
rect 7743 9193 7769 9199
rect 8135 9225 8161 9231
rect 8135 9193 8161 9199
rect 8807 9225 8833 9231
rect 8807 9193 8833 9199
rect 8919 9225 8945 9231
rect 8919 9193 8945 9199
rect 9535 9225 9561 9231
rect 9535 9193 9561 9199
rect 10151 9225 10177 9231
rect 10151 9193 10177 9199
rect 10655 9225 10681 9231
rect 10655 9193 10681 9199
rect 11047 9225 11073 9231
rect 11551 9225 11577 9231
rect 11321 9199 11327 9225
rect 11353 9199 11359 9225
rect 12889 9199 12895 9225
rect 12921 9199 12927 9225
rect 18825 9199 18831 9225
rect 18857 9199 18863 9225
rect 11047 9193 11073 9199
rect 11551 9193 11577 9199
rect 10599 9169 10625 9175
rect 14575 9169 14601 9175
rect 7625 9143 7631 9169
rect 7657 9143 7663 9169
rect 13281 9143 13287 9169
rect 13313 9143 13319 9169
rect 14345 9143 14351 9169
rect 14377 9143 14383 9169
rect 10599 9137 10625 9143
rect 14575 9137 14601 9143
rect 10263 9113 10289 9119
rect 10263 9081 10289 9087
rect 10375 9113 10401 9119
rect 10375 9081 10401 9087
rect 20007 9113 20033 9119
rect 20007 9081 20033 9087
rect 672 9029 20328 9046
rect 672 9003 2239 9029
rect 2265 9003 2291 9029
rect 2317 9003 2343 9029
rect 2369 9003 17599 9029
rect 17625 9003 17651 9029
rect 17677 9003 17703 9029
rect 17729 9003 20328 9029
rect 672 8986 20328 9003
rect 9759 8945 9785 8951
rect 9759 8913 9785 8919
rect 9199 8889 9225 8895
rect 9305 8863 9311 8889
rect 9337 8863 9343 8889
rect 9199 8857 9225 8863
rect 7407 8833 7433 8839
rect 7967 8833 7993 8839
rect 7737 8807 7743 8833
rect 7769 8807 7775 8833
rect 7407 8801 7433 8807
rect 7967 8801 7993 8807
rect 8135 8833 8161 8839
rect 8135 8801 8161 8807
rect 9031 8833 9057 8839
rect 10263 8833 10289 8839
rect 9921 8807 9927 8833
rect 9953 8807 9959 8833
rect 9031 8801 9057 8807
rect 10263 8801 10289 8807
rect 10655 8833 10681 8839
rect 10655 8801 10681 8807
rect 13343 8833 13369 8839
rect 13343 8801 13369 8807
rect 13455 8833 13481 8839
rect 13455 8801 13481 8807
rect 13567 8833 13593 8839
rect 13567 8801 13593 8807
rect 6903 8777 6929 8783
rect 6903 8745 6929 8751
rect 7239 8777 7265 8783
rect 7681 8751 7687 8777
rect 7713 8751 7719 8777
rect 8857 8751 8863 8777
rect 8889 8751 8895 8777
rect 7239 8745 7265 8751
rect 6735 8721 6761 8727
rect 6735 8689 6761 8695
rect 8079 8721 8105 8727
rect 8079 8689 8105 8695
rect 9815 8721 9841 8727
rect 13399 8721 13425 8727
rect 10089 8695 10095 8721
rect 10121 8695 10127 8721
rect 10817 8695 10823 8721
rect 10849 8695 10855 8721
rect 9815 8689 9841 8695
rect 13399 8689 13425 8695
rect 672 8637 20328 8654
rect 672 8611 9919 8637
rect 9945 8611 9971 8637
rect 9997 8611 10023 8637
rect 10049 8611 20328 8637
rect 672 8594 20328 8611
rect 7799 8553 7825 8559
rect 7799 8521 7825 8527
rect 9031 8553 9057 8559
rect 9031 8521 9057 8527
rect 9479 8553 9505 8559
rect 9479 8521 9505 8527
rect 6505 8471 6511 8497
rect 6537 8471 6543 8497
rect 9647 8441 9673 8447
rect 6169 8415 6175 8441
rect 6201 8415 6207 8441
rect 9361 8415 9367 8441
rect 9393 8415 9399 8441
rect 9647 8409 9673 8415
rect 9143 8385 9169 8391
rect 7569 8359 7575 8385
rect 7601 8359 7607 8385
rect 9143 8353 9169 8359
rect 8975 8329 9001 8335
rect 8975 8297 9001 8303
rect 9703 8329 9729 8335
rect 9703 8297 9729 8303
rect 672 8245 20328 8262
rect 672 8219 2239 8245
rect 2265 8219 2291 8245
rect 2317 8219 2343 8245
rect 2369 8219 17599 8245
rect 17625 8219 17651 8245
rect 17677 8219 17703 8245
rect 17729 8219 20328 8245
rect 672 8202 20328 8219
rect 967 8105 993 8111
rect 967 8073 993 8079
rect 20007 8105 20033 8111
rect 20007 8073 20033 8079
rect 8135 8049 8161 8055
rect 2137 8023 2143 8049
rect 2169 8023 2175 8049
rect 8135 8017 8161 8023
rect 8191 8049 8217 8055
rect 8191 8017 8217 8023
rect 9031 8049 9057 8055
rect 9031 8017 9057 8023
rect 10095 8049 10121 8055
rect 10095 8017 10121 8023
rect 11271 8049 11297 8055
rect 11271 8017 11297 8023
rect 11663 8049 11689 8055
rect 13679 8049 13705 8055
rect 13113 8023 13119 8049
rect 13145 8023 13151 8049
rect 13449 8023 13455 8049
rect 13481 8023 13487 8049
rect 11663 8017 11689 8023
rect 13679 8017 13705 8023
rect 13903 8049 13929 8055
rect 18937 8023 18943 8049
rect 18969 8023 18975 8049
rect 13903 8017 13929 8023
rect 7631 7993 7657 7999
rect 7631 7961 7657 7967
rect 7687 7993 7713 7999
rect 7687 7961 7713 7967
rect 7799 7993 7825 7999
rect 7799 7961 7825 7967
rect 7911 7993 7937 7999
rect 11439 7993 11465 7999
rect 10257 7967 10263 7993
rect 10289 7967 10295 7993
rect 7911 7961 7937 7967
rect 11439 7961 11465 7967
rect 11551 7993 11577 7999
rect 11551 7961 11577 7967
rect 11943 7993 11969 7999
rect 11943 7961 11969 7967
rect 13287 7993 13313 7999
rect 13287 7961 13313 7967
rect 14015 7993 14041 7999
rect 14015 7961 14041 7967
rect 8023 7937 8049 7943
rect 8023 7905 8049 7911
rect 8079 7937 8105 7943
rect 10655 7937 10681 7943
rect 11327 7937 11353 7943
rect 8857 7911 8863 7937
rect 8889 7911 8895 7937
rect 10817 7911 10823 7937
rect 10849 7911 10855 7937
rect 8079 7905 8105 7911
rect 10655 7905 10681 7911
rect 11327 7905 11353 7911
rect 11887 7937 11913 7943
rect 11887 7905 11913 7911
rect 11999 7937 12025 7943
rect 11999 7905 12025 7911
rect 13231 7937 13257 7943
rect 13231 7905 13257 7911
rect 13623 7937 13649 7943
rect 13623 7905 13649 7911
rect 13735 7937 13761 7943
rect 13735 7905 13761 7911
rect 13959 7937 13985 7943
rect 13959 7905 13985 7911
rect 672 7853 20328 7870
rect 672 7827 9919 7853
rect 9945 7827 9971 7853
rect 9997 7827 10023 7853
rect 10049 7827 20328 7853
rect 672 7810 20328 7827
rect 7743 7769 7769 7775
rect 7743 7737 7769 7743
rect 9143 7769 9169 7775
rect 10711 7769 10737 7775
rect 10145 7743 10151 7769
rect 10177 7743 10183 7769
rect 9143 7737 9169 7743
rect 10711 7737 10737 7743
rect 14687 7769 14713 7775
rect 14687 7737 14713 7743
rect 10319 7713 10345 7719
rect 14631 7713 14657 7719
rect 7121 7687 7127 7713
rect 7153 7687 7159 7713
rect 10425 7687 10431 7713
rect 10457 7687 10463 7713
rect 11265 7687 11271 7713
rect 11297 7687 11303 7713
rect 13393 7687 13399 7713
rect 13425 7687 13431 7713
rect 10319 7681 10345 7687
rect 14631 7681 14657 7687
rect 8919 7657 8945 7663
rect 7513 7631 7519 7657
rect 7545 7631 7551 7657
rect 8919 7625 8945 7631
rect 8975 7657 9001 7663
rect 8975 7625 9001 7631
rect 9087 7657 9113 7663
rect 9087 7625 9113 7631
rect 9367 7657 9393 7663
rect 12671 7657 12697 7663
rect 9417 7631 9423 7657
rect 9449 7631 9455 7657
rect 9641 7631 9647 7657
rect 9673 7631 9679 7657
rect 10033 7631 10039 7657
rect 10065 7631 10071 7657
rect 10705 7631 10711 7657
rect 10737 7631 10743 7657
rect 10929 7631 10935 7657
rect 10961 7631 10967 7657
rect 13001 7631 13007 7657
rect 13033 7631 13039 7657
rect 14793 7631 14799 7657
rect 14825 7631 14831 7657
rect 18825 7631 18831 7657
rect 18857 7631 18863 7657
rect 9367 7625 9393 7631
rect 12671 7625 12697 7631
rect 9031 7601 9057 7607
rect 6057 7575 6063 7601
rect 6089 7575 6095 7601
rect 9031 7569 9057 7575
rect 10543 7601 10569 7607
rect 15023 7601 15049 7607
rect 12329 7575 12335 7601
rect 12361 7575 12367 7601
rect 14457 7575 14463 7601
rect 14489 7575 14495 7601
rect 10543 7569 10569 7575
rect 15023 7569 15049 7575
rect 20007 7601 20033 7607
rect 20007 7569 20033 7575
rect 672 7461 20328 7478
rect 672 7435 2239 7461
rect 2265 7435 2291 7461
rect 2317 7435 2343 7461
rect 2369 7435 17599 7461
rect 17625 7435 17651 7461
rect 17677 7435 17703 7461
rect 17729 7435 20328 7461
rect 672 7418 20328 7435
rect 9815 7377 9841 7383
rect 9815 7345 9841 7351
rect 9927 7321 9953 7327
rect 11047 7321 11073 7327
rect 14631 7321 14657 7327
rect 7961 7295 7967 7321
rect 7993 7295 7999 7321
rect 9025 7295 9031 7321
rect 9057 7295 9063 7321
rect 10201 7295 10207 7321
rect 10233 7295 10239 7321
rect 13225 7295 13231 7321
rect 13257 7295 13263 7321
rect 14289 7295 14295 7321
rect 14321 7295 14327 7321
rect 9927 7289 9953 7295
rect 11047 7289 11073 7295
rect 14631 7289 14657 7295
rect 7687 7265 7713 7271
rect 10991 7265 11017 7271
rect 9417 7239 9423 7265
rect 9449 7239 9455 7265
rect 9697 7239 9703 7265
rect 9729 7239 9735 7265
rect 12889 7239 12895 7265
rect 12921 7239 12927 7265
rect 7687 7233 7713 7239
rect 10991 7233 11017 7239
rect 9591 7209 9617 7215
rect 9591 7177 9617 7183
rect 10039 7209 10065 7215
rect 10039 7177 10065 7183
rect 10263 7209 10289 7215
rect 10263 7177 10289 7183
rect 10375 7209 10401 7215
rect 10375 7177 10401 7183
rect 11215 7209 11241 7215
rect 11215 7177 11241 7183
rect 7743 7153 7769 7159
rect 7743 7121 7769 7127
rect 7855 7153 7881 7159
rect 11103 7153 11129 7159
rect 9753 7127 9759 7153
rect 9785 7127 9791 7153
rect 7855 7121 7881 7127
rect 11103 7121 11129 7127
rect 20119 7153 20145 7159
rect 20119 7121 20145 7127
rect 672 7069 20328 7086
rect 672 7043 9919 7069
rect 9945 7043 9971 7069
rect 9997 7043 10023 7069
rect 10049 7043 20328 7069
rect 672 7026 20328 7043
rect 8247 6985 8273 6991
rect 8247 6953 8273 6959
rect 8919 6985 8945 6991
rect 8919 6953 8945 6959
rect 9031 6985 9057 6991
rect 9031 6953 9057 6959
rect 9703 6985 9729 6991
rect 9703 6953 9729 6959
rect 12111 6985 12137 6991
rect 12111 6953 12137 6959
rect 8191 6929 8217 6935
rect 10817 6903 10823 6929
rect 10849 6903 10855 6929
rect 8191 6897 8217 6903
rect 9087 6873 9113 6879
rect 6617 6847 6623 6873
rect 6649 6847 6655 6873
rect 10481 6847 10487 6873
rect 10513 6847 10519 6873
rect 9087 6841 9113 6847
rect 9535 6817 9561 6823
rect 6953 6791 6959 6817
rect 6985 6791 6991 6817
rect 8017 6791 8023 6817
rect 8049 6791 8055 6817
rect 9535 6785 9561 6791
rect 9759 6817 9785 6823
rect 11881 6791 11887 6817
rect 11913 6791 11919 6817
rect 9759 6785 9785 6791
rect 8247 6761 8273 6767
rect 8247 6729 8273 6735
rect 672 6677 20328 6694
rect 672 6651 2239 6677
rect 2265 6651 2291 6677
rect 2317 6651 2343 6677
rect 2369 6651 17599 6677
rect 17625 6651 17651 6677
rect 17677 6651 17703 6677
rect 17729 6651 20328 6677
rect 672 6634 20328 6651
rect 8191 6537 8217 6543
rect 10375 6537 10401 6543
rect 9081 6511 9087 6537
rect 9113 6511 9119 6537
rect 10145 6511 10151 6537
rect 10177 6511 10183 6537
rect 8191 6505 8217 6511
rect 10375 6505 10401 6511
rect 8745 6455 8751 6481
rect 8777 6455 8783 6481
rect 672 6285 20328 6302
rect 672 6259 9919 6285
rect 9945 6259 9971 6285
rect 9997 6259 10023 6285
rect 10049 6259 20328 6285
rect 672 6242 20328 6259
rect 672 5893 20328 5910
rect 672 5867 2239 5893
rect 2265 5867 2291 5893
rect 2317 5867 2343 5893
rect 2369 5867 17599 5893
rect 17625 5867 17651 5893
rect 17677 5867 17703 5893
rect 17729 5867 20328 5893
rect 672 5850 20328 5867
rect 672 5501 20328 5518
rect 672 5475 9919 5501
rect 9945 5475 9971 5501
rect 9997 5475 10023 5501
rect 10049 5475 20328 5501
rect 672 5458 20328 5475
rect 672 5109 20328 5126
rect 672 5083 2239 5109
rect 2265 5083 2291 5109
rect 2317 5083 2343 5109
rect 2369 5083 17599 5109
rect 17625 5083 17651 5109
rect 17677 5083 17703 5109
rect 17729 5083 20328 5109
rect 672 5066 20328 5083
rect 672 4717 20328 4734
rect 672 4691 9919 4717
rect 9945 4691 9971 4717
rect 9997 4691 10023 4717
rect 10049 4691 20328 4717
rect 672 4674 20328 4691
rect 672 4325 20328 4342
rect 672 4299 2239 4325
rect 2265 4299 2291 4325
rect 2317 4299 2343 4325
rect 2369 4299 17599 4325
rect 17625 4299 17651 4325
rect 17677 4299 17703 4325
rect 17729 4299 20328 4325
rect 672 4282 20328 4299
rect 672 3933 20328 3950
rect 672 3907 9919 3933
rect 9945 3907 9971 3933
rect 9997 3907 10023 3933
rect 10049 3907 20328 3933
rect 672 3890 20328 3907
rect 672 3541 20328 3558
rect 672 3515 2239 3541
rect 2265 3515 2291 3541
rect 2317 3515 2343 3541
rect 2369 3515 17599 3541
rect 17625 3515 17651 3541
rect 17677 3515 17703 3541
rect 17729 3515 20328 3541
rect 672 3498 20328 3515
rect 672 3149 20328 3166
rect 672 3123 9919 3149
rect 9945 3123 9971 3149
rect 9997 3123 10023 3149
rect 10049 3123 20328 3149
rect 672 3106 20328 3123
rect 672 2757 20328 2774
rect 672 2731 2239 2757
rect 2265 2731 2291 2757
rect 2317 2731 2343 2757
rect 2369 2731 17599 2757
rect 17625 2731 17651 2757
rect 17677 2731 17703 2757
rect 17729 2731 20328 2757
rect 672 2714 20328 2731
rect 8695 2617 8721 2623
rect 8695 2585 8721 2591
rect 8185 2535 8191 2561
rect 8217 2535 8223 2561
rect 672 2365 20328 2382
rect 672 2339 9919 2365
rect 9945 2339 9971 2365
rect 9997 2339 10023 2365
rect 10049 2339 20328 2365
rect 672 2322 20328 2339
rect 9865 2143 9871 2169
rect 9897 2143 9903 2169
rect 10375 2057 10401 2063
rect 10375 2025 10401 2031
rect 672 1973 20328 1990
rect 672 1947 2239 1973
rect 2265 1947 2291 1973
rect 2317 1947 2343 1973
rect 2369 1947 17599 1973
rect 17625 1947 17651 1973
rect 17677 1947 17703 1973
rect 17729 1947 20328 1973
rect 672 1930 20328 1947
rect 9311 1833 9337 1839
rect 9311 1801 9337 1807
rect 12783 1833 12809 1839
rect 12783 1801 12809 1807
rect 8801 1751 8807 1777
rect 8833 1751 8839 1777
rect 11769 1751 11775 1777
rect 11801 1751 11807 1777
rect 12273 1751 12279 1777
rect 12305 1751 12311 1777
rect 11097 1695 11103 1721
rect 11129 1695 11135 1721
rect 672 1581 20328 1598
rect 672 1555 9919 1581
rect 9945 1555 9971 1581
rect 9997 1555 10023 1581
rect 10049 1555 20328 1581
rect 672 1538 20328 1555
<< via1 >>
rect 2239 19195 2265 19221
rect 2291 19195 2317 19221
rect 2343 19195 2369 19221
rect 17599 19195 17625 19221
rect 17651 19195 17677 19221
rect 17703 19195 17729 19221
rect 9311 19111 9337 19137
rect 11215 19111 11241 19137
rect 13063 19111 13089 19137
rect 8807 18999 8833 19025
rect 10823 18999 10849 19025
rect 12671 18999 12697 19025
rect 14239 18943 14265 18969
rect 9919 18803 9945 18829
rect 9971 18803 9997 18829
rect 10023 18803 10049 18829
rect 9927 18719 9953 18745
rect 11383 18719 11409 18745
rect 13399 18719 13425 18745
rect 9423 18607 9449 18633
rect 11103 18607 11129 18633
rect 12951 18607 12977 18633
rect 2239 18411 2265 18437
rect 2291 18411 2317 18437
rect 2343 18411 2369 18437
rect 17599 18411 17625 18437
rect 17651 18411 17677 18437
rect 17703 18411 17729 18437
rect 9031 18327 9057 18353
rect 8527 18215 8553 18241
rect 9919 18019 9945 18045
rect 9971 18019 9997 18045
rect 10023 18019 10049 18045
rect 2239 17627 2265 17653
rect 2291 17627 2317 17653
rect 2343 17627 2369 17653
rect 17599 17627 17625 17653
rect 17651 17627 17677 17653
rect 17703 17627 17729 17653
rect 9919 17235 9945 17261
rect 9971 17235 9997 17261
rect 10023 17235 10049 17261
rect 2239 16843 2265 16869
rect 2291 16843 2317 16869
rect 2343 16843 2369 16869
rect 17599 16843 17625 16869
rect 17651 16843 17677 16869
rect 17703 16843 17729 16869
rect 9919 16451 9945 16477
rect 9971 16451 9997 16477
rect 10023 16451 10049 16477
rect 2239 16059 2265 16085
rect 2291 16059 2317 16085
rect 2343 16059 2369 16085
rect 17599 16059 17625 16085
rect 17651 16059 17677 16085
rect 17703 16059 17729 16085
rect 9919 15667 9945 15693
rect 9971 15667 9997 15693
rect 10023 15667 10049 15693
rect 2239 15275 2265 15301
rect 2291 15275 2317 15301
rect 2343 15275 2369 15301
rect 17599 15275 17625 15301
rect 17651 15275 17677 15301
rect 17703 15275 17729 15301
rect 9919 14883 9945 14909
rect 9971 14883 9997 14909
rect 10023 14883 10049 14909
rect 2239 14491 2265 14517
rect 2291 14491 2317 14517
rect 2343 14491 2369 14517
rect 17599 14491 17625 14517
rect 17651 14491 17677 14517
rect 17703 14491 17729 14517
rect 9919 14099 9945 14125
rect 9971 14099 9997 14125
rect 10023 14099 10049 14125
rect 8247 14015 8273 14041
rect 12671 14015 12697 14041
rect 8135 13903 8161 13929
rect 8303 13903 8329 13929
rect 9255 13903 9281 13929
rect 10935 13903 10961 13929
rect 12615 13903 12641 13929
rect 13007 13903 13033 13929
rect 8807 13847 8833 13873
rect 9143 13847 9169 13873
rect 9647 13847 9673 13873
rect 10711 13847 10737 13873
rect 11271 13847 11297 13873
rect 12335 13847 12361 13873
rect 12671 13791 12697 13817
rect 2239 13707 2265 13733
rect 2291 13707 2317 13733
rect 2343 13707 2369 13733
rect 17599 13707 17625 13733
rect 17651 13707 17677 13733
rect 17703 13707 17729 13733
rect 8751 13567 8777 13593
rect 10375 13567 10401 13593
rect 10711 13567 10737 13593
rect 12951 13567 12977 13593
rect 13175 13567 13201 13593
rect 7295 13511 7321 13537
rect 8975 13511 9001 13537
rect 10935 13511 10961 13537
rect 11047 13511 11073 13537
rect 11495 13511 11521 13537
rect 7687 13455 7713 13481
rect 9311 13455 9337 13481
rect 10655 13455 10681 13481
rect 10767 13455 10793 13481
rect 11159 13455 11185 13481
rect 11215 13455 11241 13481
rect 11887 13455 11913 13481
rect 9919 13315 9945 13341
rect 9971 13315 9997 13341
rect 10023 13315 10049 13341
rect 9087 13231 9113 13257
rect 9647 13231 9673 13257
rect 10711 13231 10737 13257
rect 11719 13231 11745 13257
rect 12223 13231 12249 13257
rect 12559 13231 12585 13257
rect 9143 13175 9169 13201
rect 10879 13175 10905 13201
rect 11775 13175 11801 13201
rect 12167 13175 12193 13201
rect 12335 13175 12361 13201
rect 12671 13175 12697 13201
rect 6903 13119 6929 13145
rect 9759 13119 9785 13145
rect 11663 13119 11689 13145
rect 11999 13119 12025 13145
rect 12727 13119 12753 13145
rect 7239 13063 7265 13089
rect 8303 13063 8329 13089
rect 8863 13063 8889 13089
rect 9087 13007 9113 13033
rect 2239 12923 2265 12949
rect 2291 12923 2317 12949
rect 2343 12923 2369 12949
rect 17599 12923 17625 12949
rect 17651 12923 17677 12949
rect 17703 12923 17729 12949
rect 8807 12783 8833 12809
rect 7631 12727 7657 12753
rect 7799 12727 7825 12753
rect 9087 12727 9113 12753
rect 7743 12615 7769 12641
rect 8415 12615 8441 12641
rect 8751 12615 8777 12641
rect 8863 12615 8889 12641
rect 9919 12531 9945 12557
rect 9971 12531 9997 12557
rect 10023 12531 10049 12557
rect 12615 12335 12641 12361
rect 12783 12335 12809 12361
rect 12895 12335 12921 12361
rect 18943 12335 18969 12361
rect 12839 12279 12865 12305
rect 20007 12223 20033 12249
rect 2239 12139 2265 12165
rect 2291 12139 2317 12165
rect 2343 12139 2369 12165
rect 17599 12139 17625 12165
rect 17651 12139 17677 12165
rect 17703 12139 17729 12165
rect 9479 12055 9505 12081
rect 967 11999 993 12025
rect 9367 11999 9393 12025
rect 11047 11999 11073 12025
rect 11327 11999 11353 12025
rect 11887 11999 11913 12025
rect 13679 11999 13705 12025
rect 20007 11999 20033 12025
rect 2143 11943 2169 11969
rect 6791 11943 6817 11969
rect 7967 11943 7993 11969
rect 9815 11943 9841 11969
rect 9983 11943 10009 11969
rect 10823 11943 10849 11969
rect 10991 11943 11017 11969
rect 11551 11943 11577 11969
rect 11831 11943 11857 11969
rect 12223 11943 12249 11969
rect 13903 11943 13929 11969
rect 18831 11943 18857 11969
rect 8303 11887 8329 11913
rect 12615 11887 12641 11913
rect 6903 11831 6929 11857
rect 9535 11831 9561 11857
rect 9647 11831 9673 11857
rect 10879 11831 10905 11857
rect 11047 11831 11073 11857
rect 11607 11831 11633 11857
rect 11719 11831 11745 11857
rect 14015 11831 14041 11857
rect 14239 11831 14265 11857
rect 9919 11747 9945 11773
rect 9971 11747 9997 11773
rect 10023 11747 10049 11773
rect 8135 11663 8161 11689
rect 12055 11663 12081 11689
rect 12111 11663 12137 11689
rect 12167 11663 12193 11689
rect 7071 11607 7097 11633
rect 8023 11607 8049 11633
rect 9143 11607 9169 11633
rect 12279 11607 12305 11633
rect 13007 11607 13033 11633
rect 7407 11551 7433 11577
rect 7631 11551 7657 11577
rect 7743 11551 7769 11577
rect 7967 11551 7993 11577
rect 8191 11551 8217 11577
rect 9031 11551 9057 11577
rect 9367 11551 9393 11577
rect 11215 11551 11241 11577
rect 11327 11551 11353 11577
rect 11551 11551 11577 11577
rect 11663 11551 11689 11577
rect 11831 11551 11857 11577
rect 11943 11551 11969 11577
rect 12335 11551 12361 11577
rect 12615 11551 12641 11577
rect 14295 11551 14321 11577
rect 18831 11551 18857 11577
rect 6007 11495 6033 11521
rect 7687 11495 7713 11521
rect 9759 11495 9785 11521
rect 10823 11495 10849 11521
rect 11607 11495 11633 11521
rect 14071 11495 14097 11521
rect 8975 11439 9001 11465
rect 9255 11439 9281 11465
rect 20007 11439 20033 11465
rect 2239 11355 2265 11381
rect 2291 11355 2317 11381
rect 2343 11355 2369 11381
rect 17599 11355 17625 11381
rect 17651 11355 17677 11381
rect 17703 11355 17729 11381
rect 7071 11271 7097 11297
rect 7239 11271 7265 11297
rect 9031 11271 9057 11297
rect 12391 11271 12417 11297
rect 7799 11215 7825 11241
rect 9255 11215 9281 11241
rect 20007 11215 20033 11241
rect 7351 11159 7377 11185
rect 7967 11159 7993 11185
rect 9143 11159 9169 11185
rect 9311 11159 9337 11185
rect 10655 11159 10681 11185
rect 12279 11159 12305 11185
rect 13119 11159 13145 11185
rect 18831 11159 18857 11185
rect 8079 11103 8105 11129
rect 8975 11103 9001 11129
rect 9479 11103 9505 11129
rect 9703 11103 9729 11129
rect 9871 11103 9897 11129
rect 10823 11103 10849 11129
rect 11159 11103 11185 11129
rect 12559 11103 12585 11129
rect 13231 11103 13257 11129
rect 13287 11103 13313 11129
rect 14239 11103 14265 11129
rect 6903 11047 6929 11073
rect 7575 11047 7601 11073
rect 10879 11047 10905 11073
rect 12447 11047 12473 11073
rect 14071 11047 14097 11073
rect 14743 11047 14769 11073
rect 14911 11047 14937 11073
rect 9919 10963 9945 10989
rect 9971 10963 9997 10989
rect 10023 10963 10049 10989
rect 8023 10879 8049 10905
rect 9479 10879 9505 10905
rect 11663 10879 11689 10905
rect 13175 10879 13201 10905
rect 9927 10823 9953 10849
rect 10431 10823 10457 10849
rect 10599 10823 10625 10849
rect 13343 10823 13369 10849
rect 14071 10823 14097 10849
rect 5615 10767 5641 10793
rect 7463 10767 7489 10793
rect 7855 10767 7881 10793
rect 9311 10767 9337 10793
rect 10207 10767 10233 10793
rect 10711 10767 10737 10793
rect 11439 10767 11465 10793
rect 11719 10767 11745 10793
rect 11775 10767 11801 10793
rect 11887 10767 11913 10793
rect 12111 10767 12137 10793
rect 12167 10767 12193 10793
rect 13455 10767 13481 10793
rect 13679 10767 13705 10793
rect 18831 10767 18857 10793
rect 5951 10711 5977 10737
rect 7015 10711 7041 10737
rect 7183 10711 7209 10737
rect 7575 10711 7601 10737
rect 9647 10711 9673 10737
rect 11999 10711 12025 10737
rect 15135 10711 15161 10737
rect 20007 10711 20033 10737
rect 10375 10655 10401 10681
rect 2239 10571 2265 10597
rect 2291 10571 2317 10597
rect 2343 10571 2369 10597
rect 17599 10571 17625 10597
rect 17651 10571 17677 10597
rect 17703 10571 17729 10597
rect 14575 10487 14601 10513
rect 7519 10431 7545 10457
rect 7911 10431 7937 10457
rect 10879 10431 10905 10457
rect 11271 10431 11297 10457
rect 13175 10431 13201 10457
rect 14743 10431 14769 10457
rect 15023 10431 15049 10457
rect 6399 10375 6425 10401
rect 7015 10375 7041 10401
rect 7351 10375 7377 10401
rect 10039 10375 10065 10401
rect 10655 10375 10681 10401
rect 11663 10375 11689 10401
rect 15191 10375 15217 10401
rect 15303 10375 15329 10401
rect 6231 10319 6257 10345
rect 11047 10319 11073 10345
rect 11159 10319 11185 10345
rect 11327 10319 11353 10345
rect 14855 10319 14881 10345
rect 7127 10263 7153 10289
rect 10767 10263 10793 10289
rect 10879 10263 10905 10289
rect 9919 10179 9945 10205
rect 9971 10179 9997 10205
rect 10023 10179 10049 10205
rect 9367 10095 9393 10121
rect 12559 10095 12585 10121
rect 8359 10039 8385 10065
rect 8695 10039 8721 10065
rect 9423 10039 9449 10065
rect 9535 10039 9561 10065
rect 11663 10039 11689 10065
rect 12671 10039 12697 10065
rect 15023 10039 15049 10065
rect 8079 9983 8105 10009
rect 8807 9983 8833 10009
rect 9199 9983 9225 10009
rect 9703 9983 9729 10009
rect 12727 9983 12753 10009
rect 13343 9983 13369 10009
rect 18831 9983 18857 10009
rect 8023 9927 8049 9953
rect 13735 9927 13761 9953
rect 14799 9927 14825 9953
rect 9311 9871 9337 9897
rect 20007 9871 20033 9897
rect 2239 9787 2265 9813
rect 2291 9787 2317 9813
rect 2343 9787 2369 9813
rect 17599 9787 17625 9813
rect 17651 9787 17677 9813
rect 17703 9787 17729 9813
rect 8807 9647 8833 9673
rect 9143 9647 9169 9673
rect 9423 9647 9449 9673
rect 10655 9647 10681 9673
rect 11271 9647 11297 9673
rect 12335 9647 12361 9673
rect 12559 9647 12585 9673
rect 13623 9647 13649 9673
rect 20007 9647 20033 9673
rect 8471 9591 8497 9617
rect 8975 9591 9001 9617
rect 9647 9591 9673 9617
rect 9815 9591 9841 9617
rect 10151 9591 10177 9617
rect 10935 9591 10961 9617
rect 13511 9591 13537 9617
rect 13735 9591 13761 9617
rect 14071 9591 14097 9617
rect 14239 9591 14265 9617
rect 18831 9591 18857 9617
rect 8023 9535 8049 9561
rect 8191 9535 8217 9561
rect 9479 9535 9505 9561
rect 10263 9535 10289 9561
rect 13231 9535 13257 9561
rect 13847 9535 13873 9561
rect 14183 9535 14209 9561
rect 8583 9479 8609 9505
rect 10711 9479 10737 9505
rect 13287 9479 13313 9505
rect 13399 9479 13425 9505
rect 9919 9395 9945 9421
rect 9971 9395 9997 9421
rect 10023 9395 10049 9421
rect 9087 9311 9113 9337
rect 10823 9311 10849 9337
rect 10935 9311 10961 9337
rect 11215 9311 11241 9337
rect 11719 9311 11745 9337
rect 7855 9255 7881 9281
rect 7911 9255 7937 9281
rect 9703 9255 9729 9281
rect 10039 9255 10065 9281
rect 10711 9255 10737 9281
rect 6231 9199 6257 9225
rect 6567 9199 6593 9225
rect 7743 9199 7769 9225
rect 8135 9199 8161 9225
rect 8807 9199 8833 9225
rect 8919 9199 8945 9225
rect 9535 9199 9561 9225
rect 10151 9199 10177 9225
rect 10655 9199 10681 9225
rect 11047 9199 11073 9225
rect 11327 9199 11353 9225
rect 11551 9199 11577 9225
rect 12895 9199 12921 9225
rect 18831 9199 18857 9225
rect 7631 9143 7657 9169
rect 10599 9143 10625 9169
rect 13287 9143 13313 9169
rect 14351 9143 14377 9169
rect 14575 9143 14601 9169
rect 10263 9087 10289 9113
rect 10375 9087 10401 9113
rect 20007 9087 20033 9113
rect 2239 9003 2265 9029
rect 2291 9003 2317 9029
rect 2343 9003 2369 9029
rect 17599 9003 17625 9029
rect 17651 9003 17677 9029
rect 17703 9003 17729 9029
rect 9759 8919 9785 8945
rect 9199 8863 9225 8889
rect 9311 8863 9337 8889
rect 7407 8807 7433 8833
rect 7743 8807 7769 8833
rect 7967 8807 7993 8833
rect 8135 8807 8161 8833
rect 9031 8807 9057 8833
rect 9927 8807 9953 8833
rect 10263 8807 10289 8833
rect 10655 8807 10681 8833
rect 13343 8807 13369 8833
rect 13455 8807 13481 8833
rect 13567 8807 13593 8833
rect 6903 8751 6929 8777
rect 7239 8751 7265 8777
rect 7687 8751 7713 8777
rect 8863 8751 8889 8777
rect 6735 8695 6761 8721
rect 8079 8695 8105 8721
rect 9815 8695 9841 8721
rect 10095 8695 10121 8721
rect 10823 8695 10849 8721
rect 13399 8695 13425 8721
rect 9919 8611 9945 8637
rect 9971 8611 9997 8637
rect 10023 8611 10049 8637
rect 7799 8527 7825 8553
rect 9031 8527 9057 8553
rect 9479 8527 9505 8553
rect 6511 8471 6537 8497
rect 6175 8415 6201 8441
rect 9367 8415 9393 8441
rect 9647 8415 9673 8441
rect 7575 8359 7601 8385
rect 9143 8359 9169 8385
rect 8975 8303 9001 8329
rect 9703 8303 9729 8329
rect 2239 8219 2265 8245
rect 2291 8219 2317 8245
rect 2343 8219 2369 8245
rect 17599 8219 17625 8245
rect 17651 8219 17677 8245
rect 17703 8219 17729 8245
rect 967 8079 993 8105
rect 20007 8079 20033 8105
rect 2143 8023 2169 8049
rect 8135 8023 8161 8049
rect 8191 8023 8217 8049
rect 9031 8023 9057 8049
rect 10095 8023 10121 8049
rect 11271 8023 11297 8049
rect 11663 8023 11689 8049
rect 13119 8023 13145 8049
rect 13455 8023 13481 8049
rect 13679 8023 13705 8049
rect 13903 8023 13929 8049
rect 18943 8023 18969 8049
rect 7631 7967 7657 7993
rect 7687 7967 7713 7993
rect 7799 7967 7825 7993
rect 7911 7967 7937 7993
rect 10263 7967 10289 7993
rect 11439 7967 11465 7993
rect 11551 7967 11577 7993
rect 11943 7967 11969 7993
rect 13287 7967 13313 7993
rect 14015 7967 14041 7993
rect 8023 7911 8049 7937
rect 8079 7911 8105 7937
rect 8863 7911 8889 7937
rect 10655 7911 10681 7937
rect 10823 7911 10849 7937
rect 11327 7911 11353 7937
rect 11887 7911 11913 7937
rect 11999 7911 12025 7937
rect 13231 7911 13257 7937
rect 13623 7911 13649 7937
rect 13735 7911 13761 7937
rect 13959 7911 13985 7937
rect 9919 7827 9945 7853
rect 9971 7827 9997 7853
rect 10023 7827 10049 7853
rect 7743 7743 7769 7769
rect 9143 7743 9169 7769
rect 10151 7743 10177 7769
rect 10711 7743 10737 7769
rect 14687 7743 14713 7769
rect 7127 7687 7153 7713
rect 10319 7687 10345 7713
rect 10431 7687 10457 7713
rect 11271 7687 11297 7713
rect 13399 7687 13425 7713
rect 14631 7687 14657 7713
rect 7519 7631 7545 7657
rect 8919 7631 8945 7657
rect 8975 7631 9001 7657
rect 9087 7631 9113 7657
rect 9367 7631 9393 7657
rect 9423 7631 9449 7657
rect 9647 7631 9673 7657
rect 10039 7631 10065 7657
rect 10711 7631 10737 7657
rect 10935 7631 10961 7657
rect 12671 7631 12697 7657
rect 13007 7631 13033 7657
rect 14799 7631 14825 7657
rect 18831 7631 18857 7657
rect 6063 7575 6089 7601
rect 9031 7575 9057 7601
rect 10543 7575 10569 7601
rect 12335 7575 12361 7601
rect 14463 7575 14489 7601
rect 15023 7575 15049 7601
rect 20007 7575 20033 7601
rect 2239 7435 2265 7461
rect 2291 7435 2317 7461
rect 2343 7435 2369 7461
rect 17599 7435 17625 7461
rect 17651 7435 17677 7461
rect 17703 7435 17729 7461
rect 9815 7351 9841 7377
rect 7967 7295 7993 7321
rect 9031 7295 9057 7321
rect 9927 7295 9953 7321
rect 10207 7295 10233 7321
rect 11047 7295 11073 7321
rect 13231 7295 13257 7321
rect 14295 7295 14321 7321
rect 14631 7295 14657 7321
rect 7687 7239 7713 7265
rect 9423 7239 9449 7265
rect 9703 7239 9729 7265
rect 10991 7239 11017 7265
rect 12895 7239 12921 7265
rect 9591 7183 9617 7209
rect 10039 7183 10065 7209
rect 10263 7183 10289 7209
rect 10375 7183 10401 7209
rect 11215 7183 11241 7209
rect 7743 7127 7769 7153
rect 7855 7127 7881 7153
rect 9759 7127 9785 7153
rect 11103 7127 11129 7153
rect 20119 7127 20145 7153
rect 9919 7043 9945 7069
rect 9971 7043 9997 7069
rect 10023 7043 10049 7069
rect 8247 6959 8273 6985
rect 8919 6959 8945 6985
rect 9031 6959 9057 6985
rect 9703 6959 9729 6985
rect 12111 6959 12137 6985
rect 8191 6903 8217 6929
rect 10823 6903 10849 6929
rect 6623 6847 6649 6873
rect 9087 6847 9113 6873
rect 10487 6847 10513 6873
rect 6959 6791 6985 6817
rect 8023 6791 8049 6817
rect 9535 6791 9561 6817
rect 9759 6791 9785 6817
rect 11887 6791 11913 6817
rect 8247 6735 8273 6761
rect 2239 6651 2265 6677
rect 2291 6651 2317 6677
rect 2343 6651 2369 6677
rect 17599 6651 17625 6677
rect 17651 6651 17677 6677
rect 17703 6651 17729 6677
rect 8191 6511 8217 6537
rect 9087 6511 9113 6537
rect 10151 6511 10177 6537
rect 10375 6511 10401 6537
rect 8751 6455 8777 6481
rect 9919 6259 9945 6285
rect 9971 6259 9997 6285
rect 10023 6259 10049 6285
rect 2239 5867 2265 5893
rect 2291 5867 2317 5893
rect 2343 5867 2369 5893
rect 17599 5867 17625 5893
rect 17651 5867 17677 5893
rect 17703 5867 17729 5893
rect 9919 5475 9945 5501
rect 9971 5475 9997 5501
rect 10023 5475 10049 5501
rect 2239 5083 2265 5109
rect 2291 5083 2317 5109
rect 2343 5083 2369 5109
rect 17599 5083 17625 5109
rect 17651 5083 17677 5109
rect 17703 5083 17729 5109
rect 9919 4691 9945 4717
rect 9971 4691 9997 4717
rect 10023 4691 10049 4717
rect 2239 4299 2265 4325
rect 2291 4299 2317 4325
rect 2343 4299 2369 4325
rect 17599 4299 17625 4325
rect 17651 4299 17677 4325
rect 17703 4299 17729 4325
rect 9919 3907 9945 3933
rect 9971 3907 9997 3933
rect 10023 3907 10049 3933
rect 2239 3515 2265 3541
rect 2291 3515 2317 3541
rect 2343 3515 2369 3541
rect 17599 3515 17625 3541
rect 17651 3515 17677 3541
rect 17703 3515 17729 3541
rect 9919 3123 9945 3149
rect 9971 3123 9997 3149
rect 10023 3123 10049 3149
rect 2239 2731 2265 2757
rect 2291 2731 2317 2757
rect 2343 2731 2369 2757
rect 17599 2731 17625 2757
rect 17651 2731 17677 2757
rect 17703 2731 17729 2757
rect 8695 2591 8721 2617
rect 8191 2535 8217 2561
rect 9919 2339 9945 2365
rect 9971 2339 9997 2365
rect 10023 2339 10049 2365
rect 9871 2143 9897 2169
rect 10375 2031 10401 2057
rect 2239 1947 2265 1973
rect 2291 1947 2317 1973
rect 2343 1947 2369 1973
rect 17599 1947 17625 1973
rect 17651 1947 17677 1973
rect 17703 1947 17729 1973
rect 9311 1807 9337 1833
rect 12783 1807 12809 1833
rect 8807 1751 8833 1777
rect 11775 1751 11801 1777
rect 12279 1751 12305 1777
rect 11103 1695 11129 1721
rect 9919 1555 9945 1581
rect 9971 1555 9997 1581
rect 10023 1555 10049 1581
<< metal2 >>
rect 8400 20600 8456 21000
rect 9072 20600 9128 21000
rect 9408 20600 9464 21000
rect 10752 20600 10808 21000
rect 11088 20600 11144 21000
rect 12432 20600 12488 21000
rect 12768 20600 12824 21000
rect 14112 20600 14168 21000
rect 2238 19222 2370 19227
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2238 19189 2370 19194
rect 2238 18438 2370 18443
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2238 18405 2370 18410
rect 8414 18354 8442 20600
rect 9086 19138 9114 20600
rect 9310 19138 9338 19143
rect 9086 19137 9338 19138
rect 9086 19111 9311 19137
rect 9337 19111 9338 19137
rect 9086 19110 9338 19111
rect 9310 19105 9338 19110
rect 8414 18321 8442 18326
rect 8806 19025 8834 19031
rect 8806 18999 8807 19025
rect 8833 18999 8834 19025
rect 8526 18242 8554 18247
rect 8246 18241 8554 18242
rect 8246 18215 8527 18241
rect 8553 18215 8554 18241
rect 8246 18214 8554 18215
rect 2238 17654 2370 17659
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2238 17621 2370 17626
rect 2238 16870 2370 16875
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2238 16837 2370 16842
rect 2238 16086 2370 16091
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2238 16053 2370 16058
rect 2238 15302 2370 15307
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2238 15269 2370 15274
rect 2238 14518 2370 14523
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2238 14485 2370 14490
rect 8246 14041 8274 18214
rect 8526 18209 8554 18214
rect 8806 17654 8834 18999
rect 9422 18746 9450 20600
rect 9918 18830 10050 18835
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 9918 18797 10050 18802
rect 9422 18713 9450 18718
rect 9926 18746 9954 18751
rect 9926 18699 9954 18718
rect 10766 18746 10794 20600
rect 11102 19138 11130 20600
rect 11214 19138 11242 19143
rect 11102 19137 11242 19138
rect 11102 19111 11215 19137
rect 11241 19111 11242 19137
rect 11102 19110 11242 19111
rect 11214 19105 11242 19110
rect 12446 19138 12474 20600
rect 12446 19105 12474 19110
rect 10766 18713 10794 18718
rect 10822 19025 10850 19031
rect 10822 18999 10823 19025
rect 10849 18999 10850 19025
rect 9422 18633 9450 18639
rect 9422 18607 9423 18633
rect 9449 18607 9450 18633
rect 9030 18354 9058 18359
rect 9030 18307 9058 18326
rect 8246 14015 8247 14041
rect 8273 14015 8274 14041
rect 8134 13930 8162 13935
rect 7798 13929 8162 13930
rect 7798 13903 8135 13929
rect 8161 13903 8162 13929
rect 7798 13902 8162 13903
rect 2238 13734 2370 13739
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2238 13701 2370 13706
rect 7294 13538 7322 13543
rect 7182 13537 7322 13538
rect 7182 13511 7295 13537
rect 7321 13511 7322 13537
rect 7182 13510 7322 13511
rect 2086 13482 2114 13487
rect 966 12025 994 12031
rect 966 11999 967 12025
rect 993 11999 994 12025
rect 966 11802 994 11999
rect 966 11769 994 11774
rect 2086 9506 2114 13454
rect 6902 13146 6930 13151
rect 7182 13146 7210 13510
rect 7294 13505 7322 13510
rect 6902 13145 7210 13146
rect 6902 13119 6903 13145
rect 6929 13119 7210 13145
rect 6902 13118 7210 13119
rect 7686 13481 7714 13487
rect 7686 13455 7687 13481
rect 7713 13455 7714 13481
rect 2238 12950 2370 12955
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2238 12917 2370 12922
rect 2238 12166 2370 12171
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2238 12133 2370 12138
rect 2142 11970 2170 11975
rect 2142 11923 2170 11942
rect 6006 11970 6034 11975
rect 6006 11690 6034 11942
rect 6006 11521 6034 11662
rect 6006 11495 6007 11521
rect 6033 11495 6034 11521
rect 6006 11489 6034 11495
rect 6790 11969 6818 11975
rect 6790 11943 6791 11969
rect 6817 11943 6818 11969
rect 6790 11466 6818 11943
rect 6902 11970 6930 13118
rect 7238 13090 7266 13095
rect 7238 13043 7266 13062
rect 7630 13090 7658 13095
rect 7630 12753 7658 13062
rect 7686 12810 7714 13455
rect 7686 12777 7714 12782
rect 7630 12727 7631 12753
rect 7657 12727 7658 12753
rect 7630 12721 7658 12727
rect 7798 12753 7826 13902
rect 8134 13897 8162 13902
rect 8246 13090 8274 14015
rect 8750 17626 8834 17654
rect 8302 13929 8330 13935
rect 8302 13903 8303 13929
rect 8329 13903 8330 13929
rect 8302 13258 8330 13903
rect 8750 13593 8778 17626
rect 9422 15974 9450 18607
rect 9918 18046 10050 18051
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 9918 18013 10050 18018
rect 9918 17262 10050 17267
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 9918 17229 10050 17234
rect 9918 16478 10050 16483
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 9918 16445 10050 16450
rect 9366 15946 9450 15974
rect 9254 13929 9282 13935
rect 9254 13903 9255 13929
rect 9281 13903 9282 13929
rect 8806 13874 8834 13879
rect 9142 13874 9170 13879
rect 9254 13874 9282 13903
rect 8806 13873 8890 13874
rect 8806 13847 8807 13873
rect 8833 13847 8890 13873
rect 8806 13846 8890 13847
rect 8806 13841 8834 13846
rect 8750 13567 8751 13593
rect 8777 13567 8778 13593
rect 8750 13426 8778 13567
rect 8862 13538 8890 13846
rect 9142 13873 9282 13874
rect 9142 13847 9143 13873
rect 9169 13847 9282 13873
rect 9142 13846 9282 13847
rect 8974 13538 9002 13543
rect 9142 13538 9170 13846
rect 8862 13537 9170 13538
rect 8862 13511 8975 13537
rect 9001 13511 9170 13537
rect 8862 13510 9170 13511
rect 8974 13505 9002 13510
rect 9030 13454 9058 13510
rect 8750 13393 8778 13398
rect 8918 13426 9058 13454
rect 9310 13482 9338 13487
rect 9310 13435 9338 13454
rect 9086 13426 9114 13431
rect 8302 13225 8330 13230
rect 8302 13090 8330 13095
rect 8246 13089 8330 13090
rect 8246 13063 8303 13089
rect 8329 13063 8330 13089
rect 8246 13062 8330 13063
rect 8302 13057 8330 13062
rect 8862 13090 8890 13095
rect 8918 13090 8946 13426
rect 9086 13257 9114 13398
rect 9086 13231 9087 13257
rect 9113 13231 9114 13257
rect 9086 13225 9114 13231
rect 9142 13258 9170 13263
rect 9142 13201 9170 13230
rect 9142 13175 9143 13201
rect 9169 13175 9170 13201
rect 9142 13169 9170 13175
rect 8862 13089 8946 13090
rect 8862 13063 8863 13089
rect 8889 13063 8946 13089
rect 8862 13062 8946 13063
rect 8862 13057 8890 13062
rect 8806 12810 8834 12815
rect 8806 12763 8834 12782
rect 7798 12727 7799 12753
rect 7825 12727 7826 12753
rect 7798 12721 7826 12727
rect 7742 12642 7770 12647
rect 7742 12641 7882 12642
rect 7742 12615 7743 12641
rect 7769 12615 7882 12641
rect 7742 12614 7882 12615
rect 7742 12609 7770 12614
rect 6902 11937 6930 11942
rect 7574 11970 7602 11975
rect 6902 11858 6930 11863
rect 6902 11857 7098 11858
rect 6902 11831 6903 11857
rect 6929 11831 7098 11857
rect 6902 11830 7098 11831
rect 6902 11825 6930 11830
rect 7070 11633 7098 11830
rect 7070 11607 7071 11633
rect 7097 11607 7098 11633
rect 7070 11601 7098 11607
rect 7406 11578 7434 11583
rect 7238 11522 7266 11527
rect 6790 11438 7098 11466
rect 2238 11382 2370 11387
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2238 11349 2370 11354
rect 7070 11297 7098 11438
rect 7070 11271 7071 11297
rect 7097 11271 7098 11297
rect 7070 11265 7098 11271
rect 7238 11297 7266 11494
rect 7238 11271 7239 11297
rect 7265 11271 7266 11297
rect 7238 11265 7266 11271
rect 7350 11466 7378 11471
rect 7350 11185 7378 11438
rect 7350 11159 7351 11185
rect 7377 11159 7378 11185
rect 5614 11074 5642 11079
rect 5614 10793 5642 11046
rect 6902 11074 6930 11079
rect 6902 11027 6930 11046
rect 7350 10962 7378 11159
rect 7406 11074 7434 11550
rect 7574 11578 7602 11942
rect 7574 11545 7602 11550
rect 7630 11577 7658 11583
rect 7630 11551 7631 11577
rect 7657 11551 7658 11577
rect 7630 11186 7658 11551
rect 7742 11577 7770 11583
rect 7742 11551 7743 11577
rect 7769 11551 7770 11577
rect 7686 11522 7714 11527
rect 7686 11475 7714 11494
rect 7630 11153 7658 11158
rect 7406 11041 7434 11046
rect 7574 11074 7602 11079
rect 7574 11027 7602 11046
rect 7350 10934 7434 10962
rect 5614 10767 5615 10793
rect 5641 10767 5642 10793
rect 5614 10761 5642 10767
rect 7014 10794 7042 10799
rect 5950 10738 5978 10743
rect 6398 10738 6426 10743
rect 5950 10737 6258 10738
rect 5950 10711 5951 10737
rect 5977 10711 6258 10737
rect 5950 10710 6258 10711
rect 5950 10705 5978 10710
rect 2238 10598 2370 10603
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2238 10565 2370 10570
rect 6230 10345 6258 10710
rect 6398 10401 6426 10710
rect 6398 10375 6399 10401
rect 6425 10375 6426 10401
rect 6398 10369 6426 10375
rect 7014 10737 7042 10766
rect 7014 10711 7015 10737
rect 7041 10711 7042 10737
rect 7014 10401 7042 10711
rect 7182 10738 7210 10743
rect 7182 10691 7210 10710
rect 7014 10375 7015 10401
rect 7041 10375 7042 10401
rect 7014 10369 7042 10375
rect 7350 10401 7378 10407
rect 7350 10375 7351 10401
rect 7377 10375 7378 10401
rect 6230 10319 6231 10345
rect 6257 10319 6258 10345
rect 6230 10313 6258 10319
rect 7126 10290 7154 10295
rect 7350 10290 7378 10375
rect 7126 10289 7378 10290
rect 7126 10263 7127 10289
rect 7153 10263 7378 10289
rect 7126 10262 7378 10263
rect 7126 10257 7154 10262
rect 2238 9814 2370 9819
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2238 9781 2370 9786
rect 7350 9562 7378 10262
rect 7350 9529 7378 9534
rect 2086 9473 2114 9478
rect 6230 9225 6258 9231
rect 6230 9199 6231 9225
rect 6257 9199 6258 9225
rect 6230 9170 6258 9199
rect 6566 9226 6594 9231
rect 6566 9179 6594 9198
rect 2238 9030 2370 9035
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2238 8997 2370 9002
rect 6174 8442 6202 8447
rect 6230 8442 6258 9142
rect 7406 8833 7434 10934
rect 7462 10793 7490 10799
rect 7462 10767 7463 10793
rect 7489 10767 7490 10793
rect 7462 10738 7490 10767
rect 7574 10738 7602 10743
rect 7462 10705 7490 10710
rect 7518 10737 7602 10738
rect 7518 10711 7575 10737
rect 7601 10711 7602 10737
rect 7518 10710 7602 10711
rect 7518 10457 7546 10710
rect 7574 10705 7602 10710
rect 7742 10738 7770 11551
rect 7798 11241 7826 11247
rect 7798 11215 7799 11241
rect 7825 11215 7826 11241
rect 7798 11186 7826 11215
rect 7798 11153 7826 11158
rect 7854 11018 7882 12614
rect 8414 12641 8442 12647
rect 8414 12615 8415 12641
rect 8441 12615 8442 12641
rect 7966 11970 7994 11975
rect 7966 11923 7994 11942
rect 8414 11970 8442 12615
rect 8750 12641 8778 12647
rect 8862 12642 8890 12647
rect 8750 12615 8751 12641
rect 8777 12615 8778 12641
rect 8750 12082 8778 12615
rect 8750 12049 8778 12054
rect 8806 12641 8890 12642
rect 8806 12615 8863 12641
rect 8889 12615 8890 12641
rect 8806 12614 8890 12615
rect 8414 11937 8442 11942
rect 8302 11913 8330 11919
rect 8302 11887 8303 11913
rect 8329 11887 8330 11913
rect 8134 11690 8162 11695
rect 8134 11643 8162 11662
rect 8022 11633 8050 11639
rect 8022 11607 8023 11633
rect 8049 11607 8050 11633
rect 7966 11578 7994 11583
rect 8022 11578 8050 11607
rect 8302 11634 8330 11887
rect 8302 11601 8330 11606
rect 7966 11577 8050 11578
rect 7966 11551 7967 11577
rect 7993 11551 8050 11577
rect 7966 11550 8050 11551
rect 8190 11577 8218 11583
rect 8190 11551 8191 11577
rect 8217 11551 8218 11577
rect 7966 11545 7994 11550
rect 7966 11185 7994 11191
rect 7966 11159 7967 11185
rect 7993 11159 7994 11185
rect 7854 10985 7882 10990
rect 7910 11074 7938 11079
rect 7854 10794 7882 10799
rect 7854 10747 7882 10766
rect 7742 10705 7770 10710
rect 7518 10431 7519 10457
rect 7545 10431 7546 10457
rect 7518 10010 7546 10431
rect 7910 10458 7938 11046
rect 7966 10626 7994 11159
rect 8078 11130 8106 11135
rect 8022 11102 8078 11130
rect 8022 10905 8050 11102
rect 8078 11083 8106 11102
rect 8022 10879 8023 10905
rect 8049 10879 8050 10905
rect 8022 10873 8050 10879
rect 8190 10626 8218 11551
rect 8806 11466 8834 12614
rect 8862 12609 8890 12614
rect 8862 11970 8890 11975
rect 8918 11970 8946 13062
rect 9086 13033 9114 13039
rect 9086 13007 9087 13033
rect 9113 13007 9114 13033
rect 9086 12753 9114 13007
rect 9086 12727 9087 12753
rect 9113 12727 9114 12753
rect 9086 12721 9114 12727
rect 9366 12026 9394 15946
rect 9918 15694 10050 15699
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 9918 15661 10050 15666
rect 9918 14910 10050 14915
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 9918 14877 10050 14882
rect 9918 14126 10050 14131
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 9918 14093 10050 14098
rect 9646 13873 9674 13879
rect 9646 13847 9647 13873
rect 9673 13847 9674 13873
rect 9646 13594 9674 13847
rect 10710 13874 10738 13879
rect 10710 13827 10738 13846
rect 9646 13561 9674 13566
rect 10374 13594 10402 13599
rect 10710 13594 10738 13599
rect 10374 13593 10626 13594
rect 10374 13567 10375 13593
rect 10401 13567 10626 13593
rect 10374 13566 10626 13567
rect 10374 13561 10402 13566
rect 9534 13482 9562 13487
rect 9478 12082 9506 12087
rect 9478 12035 9506 12054
rect 8890 11942 8946 11970
rect 9310 12025 9394 12026
rect 9310 11999 9367 12025
rect 9393 11999 9394 12025
rect 9310 11998 9394 11999
rect 8862 11937 8890 11942
rect 9086 11858 9114 11863
rect 9030 11578 9058 11583
rect 8918 11577 9058 11578
rect 8918 11551 9031 11577
rect 9057 11551 9058 11577
rect 8918 11550 9058 11551
rect 8862 11466 8890 11471
rect 8806 11438 8862 11466
rect 8862 11433 8890 11438
rect 8918 11298 8946 11550
rect 9030 11545 9058 11550
rect 8974 11465 9002 11471
rect 8974 11439 8975 11465
rect 9001 11439 9002 11465
rect 8974 11410 9002 11439
rect 8974 11377 9002 11382
rect 9030 11298 9058 11303
rect 8918 11270 9030 11298
rect 9030 11251 9058 11270
rect 9086 11186 9114 11830
rect 9142 11634 9170 11639
rect 9142 11587 9170 11606
rect 9254 11466 9282 11471
rect 9254 11419 9282 11438
rect 9142 11410 9170 11415
rect 9170 11382 9226 11410
rect 9142 11377 9170 11382
rect 9198 11242 9226 11382
rect 9254 11242 9282 11247
rect 9198 11241 9282 11242
rect 9198 11215 9255 11241
rect 9281 11215 9282 11241
rect 9198 11214 9282 11215
rect 9254 11209 9282 11214
rect 9142 11186 9170 11191
rect 9086 11185 9170 11186
rect 9086 11159 9143 11185
rect 9169 11159 9170 11185
rect 9086 11158 9170 11159
rect 8974 11130 9002 11135
rect 8974 11083 9002 11102
rect 7966 10598 8218 10626
rect 7910 10457 8162 10458
rect 7910 10431 7911 10457
rect 7937 10431 8162 10457
rect 7910 10430 8162 10431
rect 7910 10425 7938 10430
rect 7518 9977 7546 9982
rect 8078 10009 8106 10015
rect 8078 9983 8079 10009
rect 8105 9983 8106 10009
rect 8022 9953 8050 9959
rect 8022 9927 8023 9953
rect 8049 9927 8050 9953
rect 8022 9561 8050 9927
rect 8022 9535 8023 9561
rect 8049 9535 8050 9561
rect 7910 9394 7938 9399
rect 7630 9338 7658 9343
rect 7630 9169 7658 9310
rect 7854 9281 7882 9287
rect 7854 9255 7855 9281
rect 7881 9255 7882 9281
rect 7742 9226 7770 9231
rect 7742 9179 7770 9198
rect 7630 9143 7631 9169
rect 7657 9143 7658 9169
rect 7630 9137 7658 9143
rect 7798 9170 7826 9175
rect 7406 8807 7407 8833
rect 7433 8807 7434 8833
rect 6902 8778 6930 8783
rect 7238 8778 7266 8783
rect 6902 8777 7266 8778
rect 6902 8751 6903 8777
rect 6929 8751 7239 8777
rect 7265 8751 7266 8777
rect 6902 8750 7266 8751
rect 6902 8745 6930 8750
rect 7238 8745 7266 8750
rect 7406 8778 7434 8807
rect 7406 8745 7434 8750
rect 7630 8890 7658 8895
rect 6734 8722 6762 8727
rect 6510 8721 6762 8722
rect 6510 8695 6735 8721
rect 6761 8695 6762 8721
rect 6510 8694 6762 8695
rect 6510 8497 6538 8694
rect 6734 8689 6762 8694
rect 6510 8471 6511 8497
rect 6537 8471 6538 8497
rect 6510 8465 6538 8471
rect 6174 8441 6258 8442
rect 6174 8415 6175 8441
rect 6201 8415 6258 8441
rect 6174 8414 6258 8415
rect 6174 8409 6202 8414
rect 7574 8386 7602 8391
rect 7630 8386 7658 8862
rect 7742 8834 7770 8839
rect 7742 8787 7770 8806
rect 7574 8385 7658 8386
rect 7574 8359 7575 8385
rect 7601 8359 7658 8385
rect 7574 8358 7658 8359
rect 7686 8777 7714 8783
rect 7686 8751 7687 8777
rect 7713 8751 7714 8777
rect 7574 8353 7602 8358
rect 7686 8330 7714 8751
rect 7798 8554 7826 9142
rect 7854 8834 7882 9255
rect 7910 9281 7938 9366
rect 8022 9338 8050 9535
rect 8022 9305 8050 9310
rect 7910 9255 7911 9281
rect 7937 9255 7938 9281
rect 7910 9249 7938 9255
rect 8078 9226 8106 9983
rect 8078 8890 8106 9198
rect 8134 9225 8162 10430
rect 8190 10066 8218 10598
rect 8190 10033 8218 10038
rect 8246 10682 8274 10687
rect 8190 9618 8218 9623
rect 8190 9561 8218 9590
rect 8190 9535 8191 9561
rect 8217 9535 8218 9561
rect 8190 9529 8218 9535
rect 8134 9199 8135 9225
rect 8161 9199 8162 9225
rect 8134 9170 8162 9199
rect 8134 9137 8162 9142
rect 8246 9058 8274 10654
rect 8358 10346 8386 10351
rect 8358 10065 8386 10318
rect 8358 10039 8359 10065
rect 8385 10039 8386 10065
rect 8358 10033 8386 10039
rect 8694 10066 8722 10071
rect 8694 10019 8722 10038
rect 8806 10009 8834 10015
rect 8806 9983 8807 10009
rect 8833 9983 8834 10009
rect 8806 9730 8834 9983
rect 8806 9702 8946 9730
rect 8806 9673 8834 9702
rect 8806 9647 8807 9673
rect 8833 9647 8834 9673
rect 8470 9618 8498 9623
rect 8470 9571 8498 9590
rect 8806 9618 8834 9647
rect 8806 9585 8834 9590
rect 8078 8857 8106 8862
rect 8134 9030 8274 9058
rect 8582 9505 8610 9511
rect 8582 9479 8583 9505
rect 8609 9479 8610 9505
rect 7966 8834 7994 8839
rect 7854 8833 7994 8834
rect 7854 8807 7967 8833
rect 7993 8807 7994 8833
rect 7854 8806 7994 8807
rect 7966 8801 7994 8806
rect 8134 8834 8162 9030
rect 8582 8890 8610 9479
rect 8806 9226 8834 9231
rect 8806 9179 8834 9198
rect 8918 9225 8946 9702
rect 8974 9618 9002 9623
rect 8974 9571 9002 9590
rect 9086 9337 9114 11158
rect 9142 11153 9170 11158
rect 9310 11185 9338 11998
rect 9366 11993 9394 11998
rect 9534 11857 9562 13454
rect 9918 13342 10050 13347
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 9918 13309 10050 13314
rect 9646 13258 9674 13263
rect 9646 13211 9674 13230
rect 9758 13146 9786 13151
rect 9758 13099 9786 13118
rect 10094 13146 10122 13151
rect 9918 12558 10050 12563
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 9918 12525 10050 12530
rect 9814 12082 9842 12087
rect 9814 11969 9842 12054
rect 9814 11943 9815 11969
rect 9841 11943 9842 11969
rect 9534 11831 9535 11857
rect 9561 11831 9562 11857
rect 9366 11802 9394 11807
rect 9366 11577 9394 11774
rect 9366 11551 9367 11577
rect 9393 11551 9394 11577
rect 9366 11545 9394 11551
rect 9534 11242 9562 11831
rect 9310 11159 9311 11185
rect 9337 11159 9338 11185
rect 9310 11153 9338 11159
rect 9366 11214 9562 11242
rect 9646 11857 9674 11863
rect 9646 11831 9647 11857
rect 9673 11831 9674 11857
rect 9646 11578 9674 11831
rect 9814 11802 9842 11943
rect 9982 11970 10010 11975
rect 9982 11923 10010 11942
rect 10094 11858 10122 13118
rect 10094 11825 10122 11830
rect 9198 11130 9226 11135
rect 9198 10738 9226 11102
rect 9310 10793 9338 10799
rect 9310 10767 9311 10793
rect 9337 10767 9338 10793
rect 9310 10738 9338 10767
rect 9198 10710 9338 10738
rect 9086 9311 9087 9337
rect 9113 9311 9114 9337
rect 9086 9305 9114 9311
rect 9142 10458 9170 10463
rect 9142 9673 9170 10430
rect 9198 10009 9226 10710
rect 9366 10682 9394 11214
rect 9478 11130 9506 11135
rect 9478 11129 9562 11130
rect 9478 11103 9479 11129
rect 9505 11103 9562 11129
rect 9478 11102 9562 11103
rect 9478 11097 9506 11102
rect 9478 10962 9506 10967
rect 9478 10905 9506 10934
rect 9478 10879 9479 10905
rect 9505 10879 9506 10905
rect 9478 10873 9506 10879
rect 9198 9983 9199 10009
rect 9225 9983 9226 10009
rect 9198 9977 9226 9983
rect 9254 10654 9394 10682
rect 9422 10850 9450 10855
rect 9142 9647 9143 9673
rect 9169 9647 9170 9673
rect 8918 9199 8919 9225
rect 8945 9199 8946 9225
rect 8918 9193 8946 9199
rect 9030 9226 9058 9231
rect 8582 8857 8610 8862
rect 8974 8890 9002 8895
rect 8134 8787 8162 8806
rect 8862 8778 8890 8783
rect 8862 8731 8890 8750
rect 7686 8297 7714 8302
rect 7742 8553 7826 8554
rect 7742 8527 7799 8553
rect 7825 8527 7826 8553
rect 7742 8526 7826 8527
rect 2238 8246 2370 8251
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2238 8213 2370 8218
rect 966 8105 994 8111
rect 966 8079 967 8105
rect 993 8079 994 8105
rect 966 7770 994 8079
rect 7630 8106 7658 8111
rect 2142 8050 2170 8055
rect 2142 8003 2170 8022
rect 6062 8050 6090 8055
rect 966 7737 994 7742
rect 6062 7601 6090 8022
rect 7630 7993 7658 8078
rect 7630 7967 7631 7993
rect 7657 7967 7658 7993
rect 7126 7938 7154 7943
rect 7126 7713 7154 7910
rect 7126 7687 7127 7713
rect 7153 7687 7154 7713
rect 7126 7681 7154 7687
rect 7630 7714 7658 7967
rect 7686 8050 7714 8055
rect 7686 7993 7714 8022
rect 7686 7967 7687 7993
rect 7713 7967 7714 7993
rect 7686 7961 7714 7967
rect 7742 7770 7770 8526
rect 7798 8521 7826 8526
rect 8078 8721 8106 8727
rect 8078 8695 8079 8721
rect 8105 8695 8106 8721
rect 8078 8106 8106 8695
rect 8078 8073 8106 8078
rect 8134 8722 8162 8727
rect 8134 8049 8162 8694
rect 8974 8442 9002 8862
rect 9030 8833 9058 9198
rect 9030 8807 9031 8833
rect 9057 8807 9058 8833
rect 9030 8553 9058 8807
rect 9030 8527 9031 8553
rect 9057 8527 9058 8553
rect 9030 8521 9058 8527
rect 9142 8498 9170 9647
rect 9254 9002 9282 10654
rect 9366 10121 9394 10127
rect 9366 10095 9367 10121
rect 9393 10095 9394 10121
rect 9310 9897 9338 9903
rect 9310 9871 9311 9897
rect 9337 9871 9338 9897
rect 9310 9226 9338 9871
rect 9366 9338 9394 10095
rect 9422 10065 9450 10822
rect 9534 10458 9562 11102
rect 9646 10962 9674 11550
rect 9702 11774 9814 11802
rect 9702 11129 9730 11774
rect 9814 11769 9842 11774
rect 9918 11774 10050 11779
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 9918 11741 10050 11746
rect 9758 11690 9786 11695
rect 9758 11521 9786 11662
rect 9758 11495 9759 11521
rect 9785 11495 9786 11521
rect 9758 11489 9786 11495
rect 9870 11130 9898 11135
rect 9702 11103 9703 11129
rect 9729 11103 9730 11129
rect 9702 11097 9730 11103
rect 9758 11102 9870 11130
rect 9646 10929 9674 10934
rect 9534 10425 9562 10430
rect 9646 10738 9674 10743
rect 9646 10290 9674 10710
rect 9646 10257 9674 10262
rect 9422 10039 9423 10065
rect 9449 10039 9450 10065
rect 9422 10033 9450 10039
rect 9534 10066 9562 10071
rect 9534 10019 9562 10038
rect 9702 10010 9730 10015
rect 9590 10009 9730 10010
rect 9590 9983 9703 10009
rect 9729 9983 9730 10009
rect 9590 9982 9730 9983
rect 9590 9730 9618 9982
rect 9702 9977 9730 9982
rect 9422 9702 9618 9730
rect 9422 9673 9450 9702
rect 9422 9647 9423 9673
rect 9449 9647 9450 9673
rect 9422 9506 9450 9647
rect 9646 9618 9674 9623
rect 9758 9618 9786 11102
rect 9870 11083 9898 11102
rect 9918 10990 10050 10995
rect 9814 10962 9842 10967
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 9918 10957 10050 10962
rect 10430 10962 10458 13566
rect 10598 13258 10626 13566
rect 10710 13547 10738 13566
rect 10654 13481 10682 13487
rect 10654 13455 10655 13481
rect 10681 13455 10682 13481
rect 10654 13426 10682 13455
rect 10766 13482 10794 13487
rect 10766 13435 10794 13454
rect 10654 13393 10682 13398
rect 10710 13258 10738 13263
rect 10598 13257 10738 13258
rect 10598 13231 10711 13257
rect 10737 13231 10738 13257
rect 10598 13230 10738 13231
rect 10710 13225 10738 13230
rect 10822 11969 10850 18999
rect 12670 19025 12698 19031
rect 12670 18999 12671 19025
rect 12697 18999 12698 19025
rect 11382 18746 11410 18751
rect 11382 18699 11410 18718
rect 11102 18633 11130 18639
rect 11102 18607 11103 18633
rect 11129 18607 11130 18633
rect 10934 13930 10962 13935
rect 10934 13883 10962 13902
rect 11102 13874 11130 18607
rect 12670 14042 12698 18999
rect 12782 18746 12810 20600
rect 13062 19138 13090 19143
rect 13062 19091 13090 19110
rect 14126 18970 14154 20600
rect 17598 19222 17730 19227
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17598 19189 17730 19194
rect 14238 18970 14266 18975
rect 14126 18969 14266 18970
rect 14126 18943 14239 18969
rect 14265 18943 14266 18969
rect 14126 18942 14266 18943
rect 14238 18937 14266 18942
rect 12782 18713 12810 18718
rect 13398 18746 13426 18751
rect 13398 18699 13426 18718
rect 12334 14041 12698 14042
rect 12334 14015 12671 14041
rect 12697 14015 12698 14041
rect 12334 14014 12698 14015
rect 11494 13930 11522 13935
rect 11130 13846 11186 13874
rect 11102 13841 11130 13846
rect 10934 13538 10962 13543
rect 11046 13538 11074 13543
rect 10934 13537 11074 13538
rect 10934 13511 10935 13537
rect 10961 13511 11047 13537
rect 11073 13511 11074 13537
rect 10934 13510 11074 13511
rect 10934 13505 10962 13510
rect 11046 13505 11074 13510
rect 11158 13481 11186 13846
rect 11270 13873 11298 13879
rect 11270 13847 11271 13873
rect 11297 13847 11298 13873
rect 11158 13455 11159 13481
rect 11185 13455 11186 13481
rect 11158 13449 11186 13455
rect 11214 13481 11242 13487
rect 11214 13455 11215 13481
rect 11241 13455 11242 13481
rect 10878 13202 10906 13207
rect 10878 12362 10906 13174
rect 11214 13146 11242 13455
rect 11270 13258 11298 13847
rect 11494 13538 11522 13902
rect 12334 13873 12362 14014
rect 12670 14009 12698 14014
rect 12950 18633 12978 18639
rect 12950 18607 12951 18633
rect 12977 18607 12978 18633
rect 12334 13847 12335 13873
rect 12361 13847 12362 13873
rect 12334 13841 12362 13847
rect 12614 13929 12642 13935
rect 12614 13903 12615 13929
rect 12641 13903 12642 13929
rect 11270 13225 11298 13230
rect 11326 13537 11522 13538
rect 11326 13511 11495 13537
rect 11521 13511 11522 13537
rect 11326 13510 11522 13511
rect 11214 13113 11242 13118
rect 10878 12334 11018 12362
rect 10822 11943 10823 11969
rect 10849 11943 10850 11969
rect 10822 11690 10850 11943
rect 10990 11969 11018 12334
rect 11046 12026 11074 12031
rect 11326 12026 11354 13510
rect 11494 13505 11522 13510
rect 11998 13818 12026 13823
rect 11886 13481 11914 13487
rect 11886 13455 11887 13481
rect 11913 13455 11914 13481
rect 11662 13426 11690 13431
rect 11662 13145 11690 13398
rect 11886 13314 11914 13455
rect 11886 13281 11914 13286
rect 11718 13258 11746 13263
rect 11718 13211 11746 13230
rect 11662 13119 11663 13145
rect 11689 13119 11690 13145
rect 11046 12025 11186 12026
rect 11046 11999 11047 12025
rect 11073 11999 11186 12025
rect 11046 11998 11186 11999
rect 11046 11993 11074 11998
rect 10990 11943 10991 11969
rect 11017 11943 11018 11969
rect 10990 11937 11018 11943
rect 10878 11858 10906 11863
rect 10878 11811 10906 11830
rect 11046 11857 11074 11863
rect 11046 11831 11047 11857
rect 11073 11831 11074 11857
rect 10822 11657 10850 11662
rect 10878 11634 10906 11639
rect 10822 11522 10850 11527
rect 10822 11475 10850 11494
rect 10654 11185 10682 11191
rect 10654 11159 10655 11185
rect 10681 11159 10682 11185
rect 10654 11130 10682 11159
rect 10654 11097 10682 11102
rect 10822 11129 10850 11135
rect 10822 11103 10823 11129
rect 10849 11103 10850 11129
rect 10766 10962 10794 10967
rect 9814 10066 9842 10934
rect 10430 10934 10738 10962
rect 9926 10850 9954 10855
rect 9926 10803 9954 10822
rect 10430 10849 10458 10934
rect 10430 10823 10431 10849
rect 10457 10823 10458 10849
rect 10430 10817 10458 10823
rect 10598 10850 10626 10855
rect 10206 10793 10234 10799
rect 10206 10767 10207 10793
rect 10233 10767 10234 10793
rect 10038 10402 10066 10407
rect 10038 10355 10066 10374
rect 10150 10290 10178 10295
rect 9918 10206 10050 10211
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 9918 10173 10050 10178
rect 9814 10038 10010 10066
rect 9646 9617 9786 9618
rect 9646 9591 9647 9617
rect 9673 9591 9786 9617
rect 9646 9590 9786 9591
rect 9814 9954 9842 9959
rect 9814 9617 9842 9926
rect 9814 9591 9815 9617
rect 9841 9591 9842 9617
rect 9422 9473 9450 9478
rect 9478 9561 9506 9567
rect 9478 9535 9479 9561
rect 9505 9535 9506 9561
rect 9478 9450 9506 9535
rect 9478 9417 9506 9422
rect 9366 9310 9618 9338
rect 9310 9193 9338 9198
rect 9534 9225 9562 9231
rect 9534 9199 9535 9225
rect 9561 9199 9562 9225
rect 9366 9170 9394 9175
rect 9254 8969 9282 8974
rect 9310 9058 9338 9063
rect 9198 8890 9226 8895
rect 9310 8890 9338 9030
rect 9198 8843 9226 8862
rect 9254 8889 9338 8890
rect 9254 8863 9311 8889
rect 9337 8863 9338 8889
rect 9254 8862 9338 8863
rect 9086 8470 9170 8498
rect 8974 8414 9058 8442
rect 8134 8023 8135 8049
rect 8161 8023 8162 8049
rect 8134 8017 8162 8023
rect 8190 8330 8218 8335
rect 8190 8049 8218 8302
rect 8974 8330 9002 8335
rect 8974 8283 9002 8302
rect 8190 8023 8191 8049
rect 8217 8023 8218 8049
rect 8190 8017 8218 8023
rect 9030 8049 9058 8414
rect 9030 8023 9031 8049
rect 9057 8023 9058 8049
rect 9030 8017 9058 8023
rect 7798 7994 7826 7999
rect 7910 7994 7938 7999
rect 7798 7993 7938 7994
rect 7798 7967 7799 7993
rect 7825 7967 7911 7993
rect 7937 7967 7938 7993
rect 7798 7966 7938 7967
rect 7798 7961 7826 7966
rect 7910 7961 7938 7966
rect 8022 7937 8050 7943
rect 8022 7911 8023 7937
rect 8049 7911 8050 7937
rect 7742 7769 7826 7770
rect 7742 7743 7743 7769
rect 7769 7743 7826 7769
rect 7742 7742 7826 7743
rect 7686 7714 7714 7719
rect 7630 7686 7686 7714
rect 7686 7681 7714 7686
rect 7518 7657 7546 7663
rect 7518 7631 7519 7657
rect 7545 7631 7546 7657
rect 6734 7602 6762 7607
rect 6062 7575 6063 7601
rect 6089 7575 6090 7601
rect 6062 7569 6090 7575
rect 6622 7574 6734 7602
rect 2238 7462 2370 7467
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2238 7429 2370 7434
rect 6622 6873 6650 7574
rect 6734 7569 6762 7574
rect 7518 7602 7546 7631
rect 7742 7602 7770 7742
rect 7546 7574 7770 7602
rect 7518 7555 7546 7574
rect 7686 7490 7714 7495
rect 7686 7265 7714 7462
rect 7686 7239 7687 7265
rect 7713 7239 7714 7265
rect 7686 7233 7714 7239
rect 6622 6847 6623 6873
rect 6649 6847 6650 6873
rect 6622 6841 6650 6847
rect 7742 7153 7770 7159
rect 7742 7127 7743 7153
rect 7769 7127 7770 7153
rect 6958 6817 6986 6823
rect 6958 6791 6959 6817
rect 6985 6791 6986 6817
rect 6958 6762 6986 6791
rect 6958 6729 6986 6734
rect 2238 6678 2370 6683
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2238 6645 2370 6650
rect 7742 6426 7770 7127
rect 7798 6538 7826 7742
rect 8022 7574 8050 7911
rect 8078 7938 8106 7943
rect 8078 7891 8106 7910
rect 8862 7937 8890 7943
rect 8862 7911 8863 7937
rect 8889 7911 8890 7937
rect 8246 7658 8274 7663
rect 8246 7574 8274 7630
rect 8022 7546 8274 7574
rect 7966 7322 7994 7327
rect 7966 7275 7994 7294
rect 7854 7154 7882 7159
rect 7854 7153 8218 7154
rect 7854 7127 7855 7153
rect 7881 7127 8218 7153
rect 7854 7126 8218 7127
rect 7854 7121 7882 7126
rect 8190 6929 8218 7126
rect 8246 6985 8274 7546
rect 8862 7602 8890 7911
rect 9086 7770 9114 8470
rect 9254 8442 9282 8862
rect 9310 8857 9338 8862
rect 9142 8414 9282 8442
rect 9366 8442 9394 9142
rect 9534 9114 9562 9199
rect 9478 9002 9506 9007
rect 9478 8722 9506 8974
rect 9478 8689 9506 8694
rect 9478 8554 9506 8559
rect 9534 8554 9562 9086
rect 9590 8834 9618 9310
rect 9646 9058 9674 9590
rect 9814 9506 9842 9591
rect 9982 9506 10010 10038
rect 10150 9617 10178 10262
rect 10150 9591 10151 9617
rect 10177 9591 10178 9617
rect 10150 9585 10178 9591
rect 10206 9618 10234 10767
rect 10374 10682 10402 10687
rect 10374 10635 10402 10654
rect 9982 9478 10122 9506
rect 9814 9473 9842 9478
rect 9918 9422 10050 9427
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 9918 9389 10050 9394
rect 9702 9281 9730 9287
rect 9702 9255 9703 9281
rect 9729 9255 9730 9281
rect 9702 9226 9730 9255
rect 10038 9282 10066 9287
rect 10038 9235 10066 9254
rect 9730 9198 9786 9226
rect 9702 9193 9730 9198
rect 9646 9025 9674 9030
rect 9758 8945 9786 9198
rect 9758 8919 9759 8945
rect 9785 8919 9786 8945
rect 9758 8913 9786 8919
rect 10094 8946 10122 9478
rect 10150 9226 10178 9231
rect 10206 9226 10234 9590
rect 10598 9674 10626 10822
rect 10710 10793 10738 10934
rect 10710 10767 10711 10793
rect 10737 10767 10738 10793
rect 10710 10761 10738 10767
rect 10654 10458 10682 10463
rect 10654 10401 10682 10430
rect 10654 10375 10655 10401
rect 10681 10375 10682 10401
rect 10654 10369 10682 10375
rect 10766 10289 10794 10934
rect 10766 10263 10767 10289
rect 10793 10263 10794 10289
rect 10654 9674 10682 9679
rect 10598 9673 10682 9674
rect 10598 9647 10655 9673
rect 10681 9647 10682 9673
rect 10598 9646 10682 9647
rect 10262 9561 10290 9567
rect 10262 9535 10263 9561
rect 10289 9535 10290 9561
rect 10262 9338 10290 9535
rect 10290 9310 10346 9338
rect 10262 9305 10290 9310
rect 10150 9225 10234 9226
rect 10150 9199 10151 9225
rect 10177 9199 10234 9225
rect 10150 9198 10234 9199
rect 10150 9193 10178 9198
rect 10262 9114 10290 9119
rect 10262 9067 10290 9086
rect 10094 8918 10178 8946
rect 9926 8834 9954 8839
rect 9590 8806 9786 8834
rect 9478 8553 9562 8554
rect 9478 8527 9479 8553
rect 9505 8527 9562 8553
rect 9478 8526 9562 8527
rect 9478 8521 9506 8526
rect 9646 8442 9674 8447
rect 9366 8441 9674 8442
rect 9366 8415 9367 8441
rect 9393 8415 9647 8441
rect 9673 8415 9674 8441
rect 9366 8414 9674 8415
rect 9142 8385 9170 8414
rect 9366 8409 9394 8414
rect 9646 8409 9674 8414
rect 9142 8359 9143 8385
rect 9169 8359 9170 8385
rect 9142 8353 9170 8359
rect 9702 8330 9730 8335
rect 9142 7770 9170 7775
rect 9086 7769 9450 7770
rect 9086 7743 9143 7769
rect 9169 7743 9450 7769
rect 9086 7742 9450 7743
rect 9142 7737 9170 7742
rect 8246 6959 8247 6985
rect 8273 6959 8274 6985
rect 8246 6953 8274 6959
rect 8806 7322 8834 7327
rect 8806 6986 8834 7294
rect 8190 6903 8191 6929
rect 8217 6903 8218 6929
rect 8190 6897 8218 6903
rect 7798 6505 7826 6510
rect 8022 6817 8050 6823
rect 8022 6791 8023 6817
rect 8049 6791 8050 6817
rect 8022 6426 8050 6791
rect 8246 6762 8274 6767
rect 8246 6715 8274 6734
rect 8190 6538 8218 6543
rect 8190 6491 8218 6510
rect 8750 6538 8778 6543
rect 8750 6481 8778 6510
rect 8750 6455 8751 6481
rect 8777 6455 8778 6481
rect 8750 6449 8778 6455
rect 7742 6398 8050 6426
rect 2238 5894 2370 5899
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2238 5861 2370 5866
rect 2238 5110 2370 5115
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2238 5077 2370 5082
rect 2238 4326 2370 4331
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2238 4293 2370 4298
rect 8022 4214 8050 6398
rect 8022 4186 8218 4214
rect 2238 3542 2370 3547
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2238 3509 2370 3514
rect 2238 2758 2370 2763
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2238 2725 2370 2730
rect 8078 2618 8106 2623
rect 2238 1974 2370 1979
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2238 1941 2370 1946
rect 8078 400 8106 2590
rect 8190 2561 8218 4186
rect 8694 2618 8722 2623
rect 8694 2571 8722 2590
rect 8190 2535 8191 2561
rect 8217 2535 8218 2561
rect 8190 2529 8218 2535
rect 8806 1777 8834 6958
rect 8862 6874 8890 7574
rect 8918 7657 8946 7663
rect 8918 7631 8919 7657
rect 8945 7631 8946 7657
rect 8918 6985 8946 7631
rect 8974 7658 9002 7663
rect 8974 7611 9002 7630
rect 9086 7657 9114 7663
rect 9086 7631 9087 7657
rect 9113 7631 9114 7657
rect 9030 7601 9058 7607
rect 9030 7575 9031 7601
rect 9057 7575 9058 7601
rect 9030 7321 9058 7575
rect 9086 7602 9114 7631
rect 9366 7658 9394 7663
rect 9366 7611 9394 7630
rect 9422 7657 9450 7742
rect 9422 7631 9423 7657
rect 9449 7631 9450 7657
rect 9422 7625 9450 7631
rect 9590 7658 9618 7663
rect 9086 7569 9114 7574
rect 9590 7434 9618 7630
rect 9646 7658 9674 7663
rect 9702 7658 9730 8302
rect 9646 7657 9730 7658
rect 9646 7631 9647 7657
rect 9673 7631 9730 7657
rect 9646 7630 9730 7631
rect 9646 7625 9674 7630
rect 9590 7406 9730 7434
rect 9030 7295 9031 7321
rect 9057 7295 9058 7321
rect 9030 7289 9058 7295
rect 9422 7265 9450 7271
rect 9422 7239 9423 7265
rect 9449 7239 9450 7265
rect 9142 7154 9170 7159
rect 8918 6959 8919 6985
rect 8945 6959 8946 6985
rect 8918 6953 8946 6959
rect 9030 6986 9058 6991
rect 9030 6939 9058 6958
rect 9086 6874 9114 6879
rect 8862 6873 9114 6874
rect 8862 6847 9087 6873
rect 9113 6847 9114 6873
rect 8862 6846 9114 6847
rect 9086 6841 9114 6846
rect 9086 6538 9114 6543
rect 9142 6538 9170 7126
rect 9422 6818 9450 7239
rect 9702 7265 9730 7406
rect 9758 7378 9786 8806
rect 9926 8787 9954 8806
rect 9814 8721 9842 8727
rect 9814 8695 9815 8721
rect 9841 8695 9842 8721
rect 9814 7602 9842 8695
rect 10094 8722 10122 8727
rect 10094 8675 10122 8694
rect 9918 8638 10050 8643
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 9918 8605 10050 8610
rect 10150 8386 10178 8918
rect 10262 8834 10290 8839
rect 10262 8787 10290 8806
rect 10150 8353 10178 8358
rect 10094 8330 10122 8335
rect 10094 8049 10122 8302
rect 10094 8023 10095 8049
rect 10121 8023 10122 8049
rect 10094 7938 10122 8023
rect 10262 7994 10290 7999
rect 10318 7994 10346 9310
rect 10598 9282 10626 9646
rect 10654 9641 10682 9646
rect 10598 9249 10626 9254
rect 10710 9505 10738 9511
rect 10710 9479 10711 9505
rect 10737 9479 10738 9505
rect 10710 9281 10738 9479
rect 10710 9255 10711 9281
rect 10737 9255 10738 9281
rect 10654 9226 10682 9231
rect 10654 9179 10682 9198
rect 10598 9170 10626 9175
rect 10598 9123 10626 9142
rect 10374 9113 10402 9119
rect 10374 9087 10375 9113
rect 10401 9087 10402 9113
rect 10374 8890 10402 9087
rect 10374 8857 10402 8862
rect 10654 8890 10682 8895
rect 10654 8833 10682 8862
rect 10654 8807 10655 8833
rect 10681 8807 10682 8833
rect 10654 8801 10682 8807
rect 10710 8834 10738 9255
rect 10710 8801 10738 8806
rect 10430 8386 10458 8391
rect 10262 7993 10402 7994
rect 10262 7967 10263 7993
rect 10289 7967 10402 7993
rect 10262 7966 10402 7967
rect 10262 7961 10290 7966
rect 9918 7854 10050 7859
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 9918 7821 10050 7826
rect 9814 7569 9842 7574
rect 9870 7714 9898 7719
rect 9814 7378 9842 7383
rect 9758 7377 9842 7378
rect 9758 7351 9815 7377
rect 9841 7351 9842 7377
rect 9758 7350 9842 7351
rect 9814 7345 9842 7350
rect 9702 7239 9703 7265
rect 9729 7239 9730 7265
rect 9702 7233 9730 7239
rect 9590 7210 9618 7215
rect 9870 7210 9898 7686
rect 10038 7658 10066 7663
rect 10094 7658 10122 7910
rect 10150 7770 10178 7775
rect 10318 7770 10346 7775
rect 10150 7769 10318 7770
rect 10150 7743 10151 7769
rect 10177 7743 10318 7769
rect 10150 7742 10318 7743
rect 10150 7737 10178 7742
rect 10318 7713 10346 7742
rect 10318 7687 10319 7713
rect 10345 7687 10346 7713
rect 10318 7681 10346 7687
rect 10038 7657 10122 7658
rect 10038 7631 10039 7657
rect 10065 7631 10122 7657
rect 10038 7630 10122 7631
rect 10038 7625 10066 7630
rect 10374 7574 10402 7966
rect 10430 7714 10458 8358
rect 10654 7938 10682 7943
rect 10766 7938 10794 10263
rect 10822 9506 10850 11103
rect 10878 11073 10906 11606
rect 10878 11047 10879 11073
rect 10905 11047 10906 11073
rect 10878 11041 10906 11047
rect 11046 10962 11074 11831
rect 11158 11466 11186 11998
rect 11214 11998 11326 12026
rect 11214 11577 11242 11998
rect 11326 11979 11354 11998
rect 11550 12082 11578 12087
rect 11550 11969 11578 12054
rect 11550 11943 11551 11969
rect 11577 11943 11578 11969
rect 11550 11937 11578 11943
rect 11606 11857 11634 11863
rect 11606 11831 11607 11857
rect 11633 11831 11634 11857
rect 11606 11690 11634 11831
rect 11662 11746 11690 13119
rect 11774 13202 11802 13207
rect 11774 11970 11802 13174
rect 11886 13146 11914 13151
rect 11886 12025 11914 13118
rect 11998 13145 12026 13790
rect 12166 13370 12194 13375
rect 12166 13201 12194 13342
rect 12614 13370 12642 13903
rect 12670 13818 12698 13823
rect 12670 13771 12698 13790
rect 12614 13337 12642 13342
rect 12950 13593 12978 18607
rect 17598 18438 17730 18443
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17598 18405 17730 18410
rect 17598 17654 17730 17659
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17598 17621 17730 17626
rect 17598 16870 17730 16875
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17598 16837 17730 16842
rect 17598 16086 17730 16091
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17598 16053 17730 16058
rect 17598 15302 17730 15307
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17598 15269 17730 15274
rect 17598 14518 17730 14523
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17598 14485 17730 14490
rect 13006 13930 13034 13935
rect 13034 13902 13202 13930
rect 13006 13883 13034 13902
rect 12950 13567 12951 13593
rect 12977 13567 12978 13593
rect 12558 13314 12586 13319
rect 12222 13258 12250 13263
rect 12222 13211 12250 13230
rect 12558 13257 12586 13286
rect 12558 13231 12559 13257
rect 12585 13231 12586 13257
rect 12558 13225 12586 13231
rect 12950 13258 12978 13567
rect 13174 13593 13202 13902
rect 17598 13734 17730 13739
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17598 13701 17730 13706
rect 13174 13567 13175 13593
rect 13201 13567 13202 13593
rect 13174 13561 13202 13567
rect 12950 13225 12978 13230
rect 12166 13175 12167 13201
rect 12193 13175 12194 13201
rect 12166 13169 12194 13175
rect 12334 13202 12362 13207
rect 12334 13155 12362 13174
rect 12670 13202 12698 13207
rect 12670 13155 12698 13174
rect 11998 13119 11999 13145
rect 12025 13119 12026 13145
rect 11998 13113 12026 13119
rect 12726 13146 12754 13151
rect 12726 13099 12754 13118
rect 17598 12950 17730 12955
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17598 12917 17730 12922
rect 11886 11999 11887 12025
rect 11913 11999 11914 12025
rect 11886 11993 11914 11999
rect 12110 12362 12138 12367
rect 11830 11970 11858 11975
rect 11774 11969 11858 11970
rect 11774 11943 11831 11969
rect 11857 11943 11858 11969
rect 11774 11942 11858 11943
rect 11830 11914 11858 11942
rect 11830 11886 12082 11914
rect 11718 11857 11746 11863
rect 11718 11831 11719 11857
rect 11745 11831 11746 11857
rect 11718 11802 11746 11831
rect 11718 11774 11858 11802
rect 11830 11746 11858 11774
rect 11662 11718 11802 11746
rect 11830 11718 11914 11746
rect 11606 11662 11746 11690
rect 11214 11551 11215 11577
rect 11241 11551 11242 11577
rect 11214 11545 11242 11551
rect 11326 11577 11354 11583
rect 11326 11551 11327 11577
rect 11353 11551 11354 11577
rect 11326 11466 11354 11551
rect 11550 11578 11578 11583
rect 11550 11531 11578 11550
rect 11662 11577 11690 11583
rect 11662 11551 11663 11577
rect 11689 11551 11690 11577
rect 11606 11522 11634 11527
rect 11606 11475 11634 11494
rect 11158 11438 11354 11466
rect 11662 11410 11690 11551
rect 11606 11382 11690 11410
rect 11158 11130 11186 11135
rect 11214 11130 11242 11135
rect 11158 11129 11214 11130
rect 11158 11103 11159 11129
rect 11185 11103 11214 11129
rect 11158 11102 11214 11103
rect 11158 11097 11186 11102
rect 11102 10962 11130 10967
rect 11046 10934 11102 10962
rect 11102 10929 11130 10934
rect 10878 10514 10906 10519
rect 10878 10457 10906 10486
rect 10878 10431 10879 10457
rect 10905 10431 10906 10457
rect 10878 10425 10906 10431
rect 11046 10346 11074 10351
rect 11046 10299 11074 10318
rect 11158 10345 11186 10351
rect 11158 10319 11159 10345
rect 11185 10319 11186 10345
rect 10878 10290 10906 10295
rect 10878 10243 10906 10262
rect 11158 10066 11186 10319
rect 11158 10033 11186 10038
rect 11214 9786 11242 11102
rect 11438 10794 11466 10799
rect 11606 10794 11634 11382
rect 11662 11298 11690 11303
rect 11662 10905 11690 11270
rect 11718 11074 11746 11662
rect 11774 11634 11802 11718
rect 11774 11601 11802 11606
rect 11830 11577 11858 11583
rect 11830 11551 11831 11577
rect 11857 11551 11858 11577
rect 11774 11074 11802 11079
rect 11718 11046 11774 11074
rect 11662 10879 11663 10905
rect 11689 10879 11690 10905
rect 11662 10873 11690 10879
rect 11438 10793 11634 10794
rect 11438 10767 11439 10793
rect 11465 10767 11634 10793
rect 11438 10766 11634 10767
rect 11718 10794 11746 10799
rect 11326 10682 11354 10687
rect 11270 10458 11298 10463
rect 11270 10411 11298 10430
rect 11326 10345 11354 10654
rect 11326 10319 11327 10345
rect 11353 10319 11354 10345
rect 10934 9618 10962 9623
rect 10934 9617 11018 9618
rect 10934 9591 10935 9617
rect 10961 9591 11018 9617
rect 10934 9590 11018 9591
rect 10934 9585 10962 9590
rect 10822 9337 10850 9478
rect 10822 9311 10823 9337
rect 10849 9311 10850 9337
rect 10822 9305 10850 9311
rect 10934 9338 10962 9343
rect 10934 9291 10962 9310
rect 10822 8722 10850 8727
rect 10822 8675 10850 8694
rect 10822 7938 10850 7943
rect 10766 7910 10822 7938
rect 10654 7891 10682 7910
rect 10822 7891 10850 7910
rect 10710 7770 10738 7775
rect 10710 7769 10850 7770
rect 10710 7743 10711 7769
rect 10737 7743 10850 7769
rect 10710 7742 10850 7743
rect 10710 7737 10738 7742
rect 10430 7667 10458 7686
rect 10262 7546 10402 7574
rect 10486 7658 10514 7663
rect 9926 7322 9954 7327
rect 10206 7322 10234 7327
rect 9926 7321 10234 7322
rect 9926 7295 9927 7321
rect 9953 7295 10207 7321
rect 10233 7295 10234 7321
rect 9926 7294 10234 7295
rect 9926 7289 9954 7294
rect 10206 7289 10234 7294
rect 10262 7266 10290 7546
rect 10038 7210 10066 7215
rect 9590 7209 9674 7210
rect 9590 7183 9591 7209
rect 9617 7183 9674 7209
rect 9590 7182 9674 7183
rect 9870 7209 10066 7210
rect 9870 7183 10039 7209
rect 10065 7183 10066 7209
rect 9870 7182 10066 7183
rect 9590 7177 9618 7182
rect 9646 6986 9674 7182
rect 10038 7177 10066 7182
rect 10262 7209 10290 7238
rect 10262 7183 10263 7209
rect 10289 7183 10290 7209
rect 10262 7177 10290 7183
rect 10374 7210 10402 7215
rect 10374 7163 10402 7182
rect 9758 7154 9786 7159
rect 9758 7107 9786 7126
rect 9918 7070 10050 7075
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 9918 7037 10050 7042
rect 9702 6986 9730 6991
rect 9646 6985 9730 6986
rect 9646 6959 9703 6985
rect 9729 6959 9730 6985
rect 9646 6958 9730 6959
rect 9702 6953 9730 6958
rect 10486 6873 10514 7630
rect 10710 7657 10738 7663
rect 10710 7631 10711 7657
rect 10737 7631 10738 7657
rect 10542 7602 10570 7621
rect 10542 7569 10570 7574
rect 10710 7322 10738 7631
rect 10710 7289 10738 7294
rect 10822 6929 10850 7742
rect 10934 7658 10962 7663
rect 10990 7658 11018 9590
rect 11214 9337 11242 9758
rect 11270 10122 11298 10127
rect 11270 9673 11298 10094
rect 11270 9647 11271 9673
rect 11297 9647 11298 9673
rect 11270 9641 11298 9647
rect 11326 9338 11354 10319
rect 11438 10346 11466 10766
rect 11718 10747 11746 10766
rect 11774 10793 11802 11046
rect 11830 10962 11858 11551
rect 11886 11578 11914 11718
rect 12054 11689 12082 11886
rect 12054 11663 12055 11689
rect 12081 11663 12082 11689
rect 12054 11657 12082 11663
rect 12110 11689 12138 12334
rect 12614 12361 12642 12367
rect 12614 12335 12615 12361
rect 12641 12335 12642 12361
rect 12614 12082 12642 12335
rect 12614 12049 12642 12054
rect 12782 12361 12810 12367
rect 12782 12335 12783 12361
rect 12809 12335 12810 12361
rect 12222 12026 12250 12031
rect 12222 11969 12250 11998
rect 12222 11943 12223 11969
rect 12249 11943 12250 11969
rect 12222 11937 12250 11943
rect 12558 12026 12586 12031
rect 12110 11663 12111 11689
rect 12137 11663 12138 11689
rect 12110 11657 12138 11663
rect 12166 11914 12194 11919
rect 12166 11689 12194 11886
rect 12558 11746 12586 11998
rect 12614 11914 12642 11919
rect 12614 11867 12642 11886
rect 12558 11718 12642 11746
rect 12166 11663 12167 11689
rect 12193 11663 12194 11689
rect 12166 11657 12194 11663
rect 12278 11634 12306 11639
rect 12278 11587 12306 11606
rect 12558 11634 12586 11639
rect 11942 11578 11970 11583
rect 11886 11577 11970 11578
rect 11886 11551 11943 11577
rect 11969 11551 11970 11577
rect 11886 11550 11970 11551
rect 11942 11298 11970 11550
rect 12334 11577 12362 11583
rect 12334 11551 12335 11577
rect 12361 11551 12362 11577
rect 12334 11298 12362 11551
rect 12390 11298 12418 11303
rect 12334 11297 12418 11298
rect 12334 11271 12391 11297
rect 12417 11271 12418 11297
rect 12334 11270 12418 11271
rect 11942 11265 11970 11270
rect 12390 11265 12418 11270
rect 12278 11186 12306 11191
rect 12278 11139 12306 11158
rect 12558 11129 12586 11606
rect 12614 11578 12642 11718
rect 12614 11531 12642 11550
rect 12782 11522 12810 12335
rect 12894 12362 12922 12367
rect 12894 12315 12922 12334
rect 18942 12361 18970 12367
rect 18942 12335 18943 12361
rect 18969 12335 18970 12361
rect 12838 12305 12866 12311
rect 12838 12279 12839 12305
rect 12865 12279 12866 12305
rect 12838 11634 12866 12279
rect 17598 12166 17730 12171
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17598 12133 17730 12138
rect 13678 12026 13706 12031
rect 13006 11634 13034 11639
rect 12838 11633 13034 11634
rect 12838 11607 13007 11633
rect 13033 11607 13034 11633
rect 12838 11606 13034 11607
rect 13006 11601 13034 11606
rect 13678 11634 13706 11998
rect 13902 12026 13930 12031
rect 13902 11969 13930 11998
rect 13902 11943 13903 11969
rect 13929 11943 13930 11969
rect 13902 11937 13930 11943
rect 18830 11970 18858 11975
rect 18830 11923 18858 11942
rect 14014 11858 14042 11863
rect 14014 11811 14042 11830
rect 14238 11857 14266 11863
rect 14238 11831 14239 11857
rect 14265 11831 14266 11857
rect 14238 11802 14266 11831
rect 18942 11858 18970 12335
rect 20006 12249 20034 12255
rect 20006 12223 20007 12249
rect 20033 12223 20034 12249
rect 20006 12138 20034 12223
rect 20006 12105 20034 12110
rect 18942 11825 18970 11830
rect 20006 12025 20034 12031
rect 20006 11999 20007 12025
rect 20033 11999 20034 12025
rect 20006 11802 20034 11999
rect 14238 11774 14322 11802
rect 13678 11601 13706 11606
rect 13174 11578 13202 11583
rect 12782 11494 13146 11522
rect 13118 11185 13146 11494
rect 13118 11159 13119 11185
rect 13145 11159 13146 11185
rect 13118 11153 13146 11159
rect 12558 11103 12559 11129
rect 12585 11103 12586 11129
rect 12558 11097 12586 11103
rect 12446 11074 12474 11079
rect 12446 11027 12474 11046
rect 11830 10929 11858 10934
rect 13174 10905 13202 11550
rect 14294 11578 14322 11774
rect 20006 11769 20034 11774
rect 14294 11531 14322 11550
rect 18830 11578 18858 11583
rect 18830 11531 18858 11550
rect 13230 11522 13258 11527
rect 13230 11129 13258 11494
rect 14070 11522 14098 11527
rect 14070 11475 14098 11494
rect 20006 11466 20034 11471
rect 20006 11419 20034 11438
rect 17598 11382 17730 11387
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17598 11349 17730 11354
rect 20006 11241 20034 11247
rect 20006 11215 20007 11241
rect 20033 11215 20034 11241
rect 18830 11186 18858 11191
rect 18830 11139 18858 11158
rect 13230 11103 13231 11129
rect 13257 11103 13258 11129
rect 13230 11097 13258 11103
rect 13286 11130 13314 11135
rect 13286 11083 13314 11102
rect 14238 11129 14266 11135
rect 14238 11103 14239 11129
rect 14265 11103 14266 11129
rect 13174 10879 13175 10905
rect 13201 10879 13202 10905
rect 11774 10767 11775 10793
rect 11801 10767 11802 10793
rect 11438 10313 11466 10318
rect 11662 10402 11690 10407
rect 11662 10065 11690 10374
rect 11662 10039 11663 10065
rect 11689 10039 11690 10065
rect 11662 10033 11690 10039
rect 11214 9311 11215 9337
rect 11241 9311 11242 9337
rect 11214 9305 11242 9311
rect 11270 9310 11354 9338
rect 11718 9562 11746 9567
rect 11774 9562 11802 10767
rect 11886 10793 11914 10799
rect 11886 10767 11887 10793
rect 11913 10767 11914 10793
rect 11886 10514 11914 10767
rect 12110 10793 12138 10799
rect 12110 10767 12111 10793
rect 12137 10767 12138 10793
rect 11886 10481 11914 10486
rect 11998 10737 12026 10743
rect 11998 10711 11999 10737
rect 12025 10711 12026 10737
rect 11998 10122 12026 10711
rect 11998 10089 12026 10094
rect 12110 10066 12138 10767
rect 12166 10794 12194 10799
rect 12166 10747 12194 10766
rect 13174 10794 13202 10879
rect 14070 11073 14098 11079
rect 14070 11047 14071 11073
rect 14097 11047 14098 11073
rect 13342 10850 13370 10855
rect 13342 10849 13426 10850
rect 13342 10823 13343 10849
rect 13369 10823 13426 10849
rect 13342 10822 13426 10823
rect 13342 10817 13370 10822
rect 13174 10457 13202 10766
rect 13174 10431 13175 10457
rect 13201 10431 13202 10457
rect 12110 10033 12138 10038
rect 12558 10121 12586 10127
rect 12558 10095 12559 10121
rect 12585 10095 12586 10121
rect 12558 10066 12586 10095
rect 12558 10033 12586 10038
rect 12614 10122 12642 10127
rect 12334 10010 12362 10015
rect 12334 9673 12362 9982
rect 12334 9647 12335 9673
rect 12361 9647 12362 9673
rect 12334 9641 12362 9647
rect 12558 9674 12586 9679
rect 12614 9674 12642 10094
rect 12894 10122 12922 10127
rect 12670 10066 12698 10071
rect 12670 10019 12698 10038
rect 12558 9673 12642 9674
rect 12558 9647 12559 9673
rect 12585 9647 12642 9673
rect 12558 9646 12642 9647
rect 12726 10009 12754 10015
rect 12726 9983 12727 10009
rect 12753 9983 12754 10009
rect 12558 9641 12586 9646
rect 11746 9534 11802 9562
rect 11718 9337 11746 9534
rect 11718 9311 11719 9337
rect 11745 9311 11746 9337
rect 11046 9225 11074 9231
rect 11046 9199 11047 9225
rect 11073 9199 11074 9225
rect 11046 8722 11074 9199
rect 11046 8689 11074 8694
rect 11270 8049 11298 9310
rect 11718 9305 11746 9311
rect 11326 9226 11354 9231
rect 11550 9226 11578 9231
rect 11326 9225 11578 9226
rect 11326 9199 11327 9225
rect 11353 9199 11551 9225
rect 11577 9199 11578 9225
rect 11326 9198 11578 9199
rect 11326 9114 11354 9198
rect 11550 9193 11578 9198
rect 12726 9170 12754 9983
rect 12726 9137 12754 9142
rect 12894 9225 12922 10094
rect 13174 10122 13202 10431
rect 13174 10089 13202 10094
rect 13342 10122 13370 10127
rect 13342 10009 13370 10094
rect 13398 10094 13426 10822
rect 14070 10849 14098 11047
rect 14070 10823 14071 10849
rect 14097 10823 14098 10849
rect 14070 10817 14098 10823
rect 13454 10793 13482 10799
rect 13454 10767 13455 10793
rect 13481 10767 13482 10793
rect 13454 10458 13482 10767
rect 13678 10794 13706 10799
rect 13678 10747 13706 10766
rect 14238 10514 14266 11103
rect 20006 11130 20034 11215
rect 20006 11097 20034 11102
rect 14742 11073 14770 11079
rect 14742 11047 14743 11073
rect 14769 11047 14770 11073
rect 14742 10738 14770 11047
rect 14910 11074 14938 11079
rect 14910 11027 14938 11046
rect 18830 10793 18858 10799
rect 18830 10767 18831 10793
rect 18857 10767 18858 10793
rect 14742 10705 14770 10710
rect 15134 10738 15162 10743
rect 15134 10682 15162 10710
rect 15134 10654 15274 10682
rect 14238 10481 14266 10486
rect 14574 10514 14602 10519
rect 14574 10467 14602 10486
rect 13454 10425 13482 10430
rect 14742 10458 14770 10463
rect 15022 10458 15050 10463
rect 14742 10457 15050 10458
rect 14742 10431 14743 10457
rect 14769 10431 15023 10457
rect 15049 10431 15050 10457
rect 14742 10430 15050 10431
rect 14742 10425 14770 10430
rect 15022 10425 15050 10430
rect 15190 10401 15218 10407
rect 15190 10375 15191 10401
rect 15217 10375 15218 10401
rect 14854 10346 14882 10351
rect 14854 10299 14882 10318
rect 14518 10122 14546 10127
rect 13398 10066 13594 10094
rect 13342 9983 13343 10009
rect 13369 9983 13370 10009
rect 13342 9977 13370 9983
rect 13510 9617 13538 9623
rect 13510 9591 13511 9617
rect 13537 9591 13538 9617
rect 13230 9562 13258 9567
rect 13230 9515 13258 9534
rect 13286 9505 13314 9511
rect 13286 9479 13287 9505
rect 13313 9479 13314 9505
rect 13286 9282 13314 9479
rect 13286 9249 13314 9254
rect 13398 9505 13426 9511
rect 13398 9479 13399 9505
rect 13425 9479 13426 9505
rect 12894 9199 12895 9225
rect 12921 9199 12922 9225
rect 11326 9081 11354 9086
rect 11270 8023 11271 8049
rect 11297 8023 11298 8049
rect 11270 8017 11298 8023
rect 11662 8722 11690 8727
rect 11662 8049 11690 8694
rect 11662 8023 11663 8049
rect 11689 8023 11690 8049
rect 11438 7993 11466 7999
rect 11438 7967 11439 7993
rect 11465 7967 11466 7993
rect 11326 7937 11354 7943
rect 11326 7911 11327 7937
rect 11353 7911 11354 7937
rect 11270 7714 11298 7719
rect 11326 7714 11354 7911
rect 11438 7770 11466 7967
rect 11550 7994 11578 7999
rect 11550 7947 11578 7966
rect 11438 7737 11466 7742
rect 11270 7713 11354 7714
rect 11270 7687 11271 7713
rect 11297 7687 11354 7713
rect 11270 7686 11354 7687
rect 11270 7681 11298 7686
rect 10962 7630 11018 7658
rect 10934 7611 10962 7630
rect 11046 7322 11074 7327
rect 11046 7275 11074 7294
rect 10990 7266 11018 7271
rect 10990 7219 11018 7238
rect 11214 7210 11242 7215
rect 11214 7163 11242 7182
rect 11662 7210 11690 8023
rect 11942 7994 11970 7999
rect 11942 7947 11970 7966
rect 11886 7937 11914 7943
rect 11886 7911 11887 7937
rect 11913 7911 11914 7937
rect 11886 7658 11914 7911
rect 11998 7938 12026 7943
rect 11998 7891 12026 7910
rect 11886 7630 12250 7658
rect 12222 7574 12250 7630
rect 12670 7657 12698 7663
rect 12670 7631 12671 7657
rect 12697 7631 12698 7657
rect 12334 7601 12362 7607
rect 12334 7575 12335 7601
rect 12361 7575 12362 7601
rect 12334 7574 12362 7575
rect 11662 7177 11690 7182
rect 12110 7546 12138 7551
rect 12222 7546 12362 7574
rect 12670 7546 12698 7631
rect 10822 6903 10823 6929
rect 10849 6903 10850 6929
rect 10822 6897 10850 6903
rect 11102 7153 11130 7159
rect 11102 7127 11103 7153
rect 11129 7127 11130 7153
rect 10486 6847 10487 6873
rect 10513 6847 10514 6873
rect 10486 6841 10514 6847
rect 9534 6818 9562 6823
rect 9422 6817 9562 6818
rect 9422 6791 9535 6817
rect 9561 6791 9562 6817
rect 9422 6790 9562 6791
rect 9086 6537 9170 6538
rect 9086 6511 9087 6537
rect 9113 6511 9170 6537
rect 9086 6510 9170 6511
rect 9534 6538 9562 6790
rect 9086 6505 9114 6510
rect 9534 6505 9562 6510
rect 9758 6817 9786 6823
rect 9758 6791 9759 6817
rect 9785 6791 9786 6817
rect 9758 6482 9786 6791
rect 11102 6818 11130 7127
rect 12110 6985 12138 7518
rect 12110 6959 12111 6985
rect 12137 6959 12138 6985
rect 12110 6953 12138 6959
rect 11102 6785 11130 6790
rect 11886 6818 11914 6823
rect 10150 6538 10178 6543
rect 9982 6537 10178 6538
rect 9982 6511 10151 6537
rect 10177 6511 10178 6537
rect 9982 6510 10178 6511
rect 9982 6482 10010 6510
rect 10150 6505 10178 6510
rect 10374 6538 10402 6543
rect 10374 6491 10402 6510
rect 9758 6454 10010 6482
rect 9814 2170 9842 6454
rect 9918 6286 10050 6291
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 9918 6253 10050 6258
rect 9918 5502 10050 5507
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 9918 5469 10050 5474
rect 9918 4718 10050 4723
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 9918 4685 10050 4690
rect 11886 4214 11914 6790
rect 11774 4186 11914 4214
rect 9918 3934 10050 3939
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 9918 3901 10050 3906
rect 9918 3150 10050 3155
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 9918 3117 10050 3122
rect 9918 2366 10050 2371
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 9918 2333 10050 2338
rect 9870 2170 9898 2175
rect 9814 2169 9898 2170
rect 9814 2143 9871 2169
rect 9897 2143 9898 2169
rect 9814 2142 9898 2143
rect 9870 2137 9898 2142
rect 9758 2058 9786 2063
rect 9310 1834 9338 1839
rect 8806 1751 8807 1777
rect 8833 1751 8834 1777
rect 8806 1745 8834 1751
rect 9086 1833 9338 1834
rect 9086 1807 9311 1833
rect 9337 1807 9338 1833
rect 9086 1806 9338 1807
rect 9086 400 9114 1806
rect 9310 1801 9338 1806
rect 9758 400 9786 2030
rect 10374 2058 10402 2063
rect 10374 2011 10402 2030
rect 11774 1777 11802 4186
rect 11774 1751 11775 1777
rect 11801 1751 11802 1777
rect 11774 1745 11802 1751
rect 11886 1834 11914 1839
rect 11102 1721 11130 1727
rect 11102 1695 11103 1721
rect 11129 1695 11130 1721
rect 9918 1582 10050 1587
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 9918 1549 10050 1554
rect 11102 400 11130 1695
rect 11886 490 11914 1806
rect 12278 1777 12306 7546
rect 12670 7513 12698 7518
rect 12894 7546 12922 9199
rect 13286 9169 13314 9175
rect 13286 9143 13287 9169
rect 13313 9143 13314 9169
rect 13286 8722 13314 9143
rect 13342 8834 13370 8839
rect 13398 8834 13426 9479
rect 13510 9226 13538 9591
rect 13510 9193 13538 9198
rect 13566 9506 13594 10066
rect 14518 10066 14546 10094
rect 15022 10066 15050 10071
rect 14518 10065 15050 10066
rect 14518 10039 15023 10065
rect 15049 10039 15050 10065
rect 14518 10038 15050 10039
rect 13734 9954 13762 9959
rect 13622 9953 13762 9954
rect 13622 9927 13735 9953
rect 13761 9927 13762 9953
rect 13622 9926 13762 9927
rect 13622 9673 13650 9926
rect 13734 9921 13762 9926
rect 14182 9954 14210 9959
rect 13622 9647 13623 9673
rect 13649 9647 13650 9673
rect 13622 9641 13650 9647
rect 13734 9646 13930 9674
rect 13734 9617 13762 9646
rect 13734 9591 13735 9617
rect 13761 9591 13762 9617
rect 13734 9585 13762 9591
rect 13902 9618 13930 9646
rect 14070 9618 14098 9623
rect 13902 9617 14098 9618
rect 13902 9591 14071 9617
rect 14097 9591 14098 9617
rect 13902 9590 14098 9591
rect 14070 9585 14098 9590
rect 13846 9561 13874 9567
rect 13846 9535 13847 9561
rect 13873 9535 13874 9561
rect 13846 9506 13874 9535
rect 14182 9561 14210 9926
rect 14238 9786 14266 9791
rect 14238 9617 14266 9758
rect 14238 9591 14239 9617
rect 14265 9591 14266 9617
rect 14238 9585 14266 9591
rect 14182 9535 14183 9561
rect 14209 9535 14210 9561
rect 14182 9529 14210 9535
rect 13566 9478 13874 9506
rect 13342 8833 13426 8834
rect 13342 8807 13343 8833
rect 13369 8807 13426 8833
rect 13342 8806 13426 8807
rect 13454 9058 13482 9063
rect 13454 8833 13482 9030
rect 13454 8807 13455 8833
rect 13481 8807 13482 8833
rect 13342 8801 13370 8806
rect 13398 8722 13426 8727
rect 13286 8721 13426 8722
rect 13286 8695 13399 8721
rect 13425 8695 13426 8721
rect 13286 8694 13426 8695
rect 13398 8689 13426 8694
rect 13118 8050 13146 8055
rect 13118 8003 13146 8022
rect 13454 8049 13482 8807
rect 13454 8023 13455 8049
rect 13481 8023 13482 8049
rect 13454 8017 13482 8023
rect 13566 8833 13594 9478
rect 14350 9170 14378 9175
rect 14518 9170 14546 10038
rect 15022 10033 15050 10038
rect 14798 9954 14826 9959
rect 14798 9907 14826 9926
rect 15190 9786 15218 10375
rect 15246 10402 15274 10654
rect 17598 10598 17730 10603
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17598 10565 17730 10570
rect 15302 10402 15330 10407
rect 15246 10374 15302 10402
rect 15302 10355 15330 10374
rect 18830 10402 18858 10767
rect 20006 10794 20034 10799
rect 20006 10737 20034 10766
rect 20006 10711 20007 10737
rect 20033 10711 20034 10737
rect 20006 10705 20034 10711
rect 18830 10369 18858 10374
rect 18830 10010 18858 10015
rect 18830 9963 18858 9982
rect 18830 9898 18858 9903
rect 17598 9814 17730 9819
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17598 9781 17730 9786
rect 15190 9753 15218 9758
rect 18830 9617 18858 9870
rect 20006 9897 20034 9903
rect 20006 9871 20007 9897
rect 20033 9871 20034 9897
rect 20006 9786 20034 9871
rect 20006 9753 20034 9758
rect 18830 9591 18831 9617
rect 18857 9591 18858 9617
rect 18830 9585 18858 9591
rect 20006 9673 20034 9679
rect 20006 9647 20007 9673
rect 20033 9647 20034 9673
rect 20006 9450 20034 9647
rect 20006 9417 20034 9422
rect 18830 9226 18858 9231
rect 18830 9179 18858 9198
rect 14574 9170 14602 9175
rect 14518 9169 14602 9170
rect 14518 9143 14575 9169
rect 14601 9143 14602 9169
rect 14518 9142 14602 9143
rect 14350 9123 14378 9142
rect 13566 8807 13567 8833
rect 13593 8807 13594 8833
rect 13566 8050 13594 8807
rect 13566 8017 13594 8022
rect 13678 8050 13706 8055
rect 13902 8050 13930 8055
rect 13678 8049 13930 8050
rect 13678 8023 13679 8049
rect 13705 8023 13903 8049
rect 13929 8023 13930 8049
rect 13678 8022 13930 8023
rect 13678 8017 13706 8022
rect 13902 8017 13930 8022
rect 14014 8050 14042 8055
rect 13286 7994 13314 7999
rect 13286 7947 13314 7966
rect 14014 7993 14042 8022
rect 14014 7967 14015 7993
rect 14041 7967 14042 7993
rect 14014 7961 14042 7967
rect 13230 7937 13258 7943
rect 13230 7911 13231 7937
rect 13257 7911 13258 7937
rect 13006 7657 13034 7663
rect 13006 7631 13007 7657
rect 13033 7631 13034 7657
rect 13006 7546 13034 7631
rect 12922 7518 13034 7546
rect 12894 7265 12922 7518
rect 13230 7321 13258 7911
rect 13398 7938 13426 7943
rect 13398 7713 13426 7910
rect 13398 7687 13399 7713
rect 13425 7687 13426 7713
rect 13398 7681 13426 7687
rect 13622 7937 13650 7943
rect 13622 7911 13623 7937
rect 13649 7911 13650 7937
rect 13622 7602 13650 7911
rect 13734 7937 13762 7943
rect 13734 7911 13735 7937
rect 13761 7911 13762 7937
rect 13734 7770 13762 7911
rect 13958 7938 13986 7943
rect 13958 7891 13986 7910
rect 13734 7737 13762 7742
rect 13622 7569 13650 7574
rect 14294 7714 14322 7719
rect 13230 7295 13231 7321
rect 13257 7295 13258 7321
rect 13230 7289 13258 7295
rect 14294 7321 14322 7686
rect 14462 7602 14490 7607
rect 14462 7555 14490 7574
rect 14294 7295 14295 7321
rect 14321 7295 14322 7321
rect 14294 7289 14322 7295
rect 14574 7322 14602 9142
rect 20006 9114 20034 9119
rect 20006 9067 20034 9086
rect 17598 9030 17730 9035
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17598 8997 17730 9002
rect 17598 8246 17730 8251
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17598 8213 17730 8218
rect 20006 8105 20034 8111
rect 20006 8079 20007 8105
rect 20033 8079 20034 8105
rect 18942 8049 18970 8055
rect 18942 8023 18943 8049
rect 18969 8023 18970 8049
rect 14686 7994 14714 7999
rect 14630 7770 14658 7775
rect 14630 7713 14658 7742
rect 14686 7769 14714 7966
rect 14686 7743 14687 7769
rect 14713 7743 14714 7769
rect 14686 7737 14714 7743
rect 14630 7687 14631 7713
rect 14657 7687 14658 7713
rect 14630 7681 14658 7687
rect 14798 7714 14826 7719
rect 14798 7657 14826 7686
rect 14798 7631 14799 7657
rect 14825 7631 14826 7657
rect 14798 7625 14826 7631
rect 18830 7658 18858 7663
rect 18830 7611 18858 7630
rect 15022 7601 15050 7607
rect 15022 7575 15023 7601
rect 15049 7575 15050 7601
rect 14630 7322 14658 7327
rect 15022 7322 15050 7575
rect 18942 7602 18970 8023
rect 20006 7770 20034 8079
rect 20006 7737 20034 7742
rect 18942 7569 18970 7574
rect 20006 7601 20034 7607
rect 20006 7575 20007 7601
rect 20033 7575 20034 7601
rect 17598 7462 17730 7467
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17598 7429 17730 7434
rect 20006 7434 20034 7575
rect 20006 7401 20034 7406
rect 14574 7321 15050 7322
rect 14574 7295 14631 7321
rect 14657 7295 15050 7321
rect 14574 7294 15050 7295
rect 14630 7289 14658 7294
rect 12894 7239 12895 7265
rect 12921 7239 12922 7265
rect 12894 7233 12922 7239
rect 20118 7153 20146 7159
rect 20118 7127 20119 7153
rect 20145 7127 20146 7153
rect 20118 7098 20146 7127
rect 20118 7065 20146 7070
rect 17598 6678 17730 6683
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17598 6645 17730 6650
rect 17598 5894 17730 5899
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17598 5861 17730 5866
rect 17598 5110 17730 5115
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17598 5077 17730 5082
rect 17598 4326 17730 4331
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17598 4293 17730 4298
rect 17598 3542 17730 3547
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17598 3509 17730 3514
rect 17598 2758 17730 2763
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17598 2725 17730 2730
rect 17598 1974 17730 1979
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17598 1941 17730 1946
rect 12782 1834 12810 1839
rect 12782 1787 12810 1806
rect 12278 1751 12279 1777
rect 12305 1751 12306 1777
rect 12278 1745 12306 1751
rect 11774 462 11914 490
rect 11774 400 11802 462
rect 8064 0 8120 400
rect 9072 0 9128 400
rect 9744 0 9800 400
rect 11088 0 11144 400
rect 11760 0 11816 400
<< via2 >>
rect 2238 19221 2266 19222
rect 2238 19195 2239 19221
rect 2239 19195 2265 19221
rect 2265 19195 2266 19221
rect 2238 19194 2266 19195
rect 2290 19221 2318 19222
rect 2290 19195 2291 19221
rect 2291 19195 2317 19221
rect 2317 19195 2318 19221
rect 2290 19194 2318 19195
rect 2342 19221 2370 19222
rect 2342 19195 2343 19221
rect 2343 19195 2369 19221
rect 2369 19195 2370 19221
rect 2342 19194 2370 19195
rect 2238 18437 2266 18438
rect 2238 18411 2239 18437
rect 2239 18411 2265 18437
rect 2265 18411 2266 18437
rect 2238 18410 2266 18411
rect 2290 18437 2318 18438
rect 2290 18411 2291 18437
rect 2291 18411 2317 18437
rect 2317 18411 2318 18437
rect 2290 18410 2318 18411
rect 2342 18437 2370 18438
rect 2342 18411 2343 18437
rect 2343 18411 2369 18437
rect 2369 18411 2370 18437
rect 2342 18410 2370 18411
rect 8414 18326 8442 18354
rect 2238 17653 2266 17654
rect 2238 17627 2239 17653
rect 2239 17627 2265 17653
rect 2265 17627 2266 17653
rect 2238 17626 2266 17627
rect 2290 17653 2318 17654
rect 2290 17627 2291 17653
rect 2291 17627 2317 17653
rect 2317 17627 2318 17653
rect 2290 17626 2318 17627
rect 2342 17653 2370 17654
rect 2342 17627 2343 17653
rect 2343 17627 2369 17653
rect 2369 17627 2370 17653
rect 2342 17626 2370 17627
rect 2238 16869 2266 16870
rect 2238 16843 2239 16869
rect 2239 16843 2265 16869
rect 2265 16843 2266 16869
rect 2238 16842 2266 16843
rect 2290 16869 2318 16870
rect 2290 16843 2291 16869
rect 2291 16843 2317 16869
rect 2317 16843 2318 16869
rect 2290 16842 2318 16843
rect 2342 16869 2370 16870
rect 2342 16843 2343 16869
rect 2343 16843 2369 16869
rect 2369 16843 2370 16869
rect 2342 16842 2370 16843
rect 2238 16085 2266 16086
rect 2238 16059 2239 16085
rect 2239 16059 2265 16085
rect 2265 16059 2266 16085
rect 2238 16058 2266 16059
rect 2290 16085 2318 16086
rect 2290 16059 2291 16085
rect 2291 16059 2317 16085
rect 2317 16059 2318 16085
rect 2290 16058 2318 16059
rect 2342 16085 2370 16086
rect 2342 16059 2343 16085
rect 2343 16059 2369 16085
rect 2369 16059 2370 16085
rect 2342 16058 2370 16059
rect 2238 15301 2266 15302
rect 2238 15275 2239 15301
rect 2239 15275 2265 15301
rect 2265 15275 2266 15301
rect 2238 15274 2266 15275
rect 2290 15301 2318 15302
rect 2290 15275 2291 15301
rect 2291 15275 2317 15301
rect 2317 15275 2318 15301
rect 2290 15274 2318 15275
rect 2342 15301 2370 15302
rect 2342 15275 2343 15301
rect 2343 15275 2369 15301
rect 2369 15275 2370 15301
rect 2342 15274 2370 15275
rect 2238 14517 2266 14518
rect 2238 14491 2239 14517
rect 2239 14491 2265 14517
rect 2265 14491 2266 14517
rect 2238 14490 2266 14491
rect 2290 14517 2318 14518
rect 2290 14491 2291 14517
rect 2291 14491 2317 14517
rect 2317 14491 2318 14517
rect 2290 14490 2318 14491
rect 2342 14517 2370 14518
rect 2342 14491 2343 14517
rect 2343 14491 2369 14517
rect 2369 14491 2370 14517
rect 2342 14490 2370 14491
rect 9918 18829 9946 18830
rect 9918 18803 9919 18829
rect 9919 18803 9945 18829
rect 9945 18803 9946 18829
rect 9918 18802 9946 18803
rect 9970 18829 9998 18830
rect 9970 18803 9971 18829
rect 9971 18803 9997 18829
rect 9997 18803 9998 18829
rect 9970 18802 9998 18803
rect 10022 18829 10050 18830
rect 10022 18803 10023 18829
rect 10023 18803 10049 18829
rect 10049 18803 10050 18829
rect 10022 18802 10050 18803
rect 9422 18718 9450 18746
rect 9926 18745 9954 18746
rect 9926 18719 9927 18745
rect 9927 18719 9953 18745
rect 9953 18719 9954 18745
rect 9926 18718 9954 18719
rect 12446 19110 12474 19138
rect 10766 18718 10794 18746
rect 9030 18353 9058 18354
rect 9030 18327 9031 18353
rect 9031 18327 9057 18353
rect 9057 18327 9058 18353
rect 9030 18326 9058 18327
rect 2238 13733 2266 13734
rect 2238 13707 2239 13733
rect 2239 13707 2265 13733
rect 2265 13707 2266 13733
rect 2238 13706 2266 13707
rect 2290 13733 2318 13734
rect 2290 13707 2291 13733
rect 2291 13707 2317 13733
rect 2317 13707 2318 13733
rect 2290 13706 2318 13707
rect 2342 13733 2370 13734
rect 2342 13707 2343 13733
rect 2343 13707 2369 13733
rect 2369 13707 2370 13733
rect 2342 13706 2370 13707
rect 2086 13454 2114 13482
rect 966 11774 994 11802
rect 2238 12949 2266 12950
rect 2238 12923 2239 12949
rect 2239 12923 2265 12949
rect 2265 12923 2266 12949
rect 2238 12922 2266 12923
rect 2290 12949 2318 12950
rect 2290 12923 2291 12949
rect 2291 12923 2317 12949
rect 2317 12923 2318 12949
rect 2290 12922 2318 12923
rect 2342 12949 2370 12950
rect 2342 12923 2343 12949
rect 2343 12923 2369 12949
rect 2369 12923 2370 12949
rect 2342 12922 2370 12923
rect 2238 12165 2266 12166
rect 2238 12139 2239 12165
rect 2239 12139 2265 12165
rect 2265 12139 2266 12165
rect 2238 12138 2266 12139
rect 2290 12165 2318 12166
rect 2290 12139 2291 12165
rect 2291 12139 2317 12165
rect 2317 12139 2318 12165
rect 2290 12138 2318 12139
rect 2342 12165 2370 12166
rect 2342 12139 2343 12165
rect 2343 12139 2369 12165
rect 2369 12139 2370 12165
rect 2342 12138 2370 12139
rect 2142 11969 2170 11970
rect 2142 11943 2143 11969
rect 2143 11943 2169 11969
rect 2169 11943 2170 11969
rect 2142 11942 2170 11943
rect 6006 11942 6034 11970
rect 6006 11662 6034 11690
rect 7238 13089 7266 13090
rect 7238 13063 7239 13089
rect 7239 13063 7265 13089
rect 7265 13063 7266 13089
rect 7238 13062 7266 13063
rect 7630 13062 7658 13090
rect 7686 12782 7714 12810
rect 9918 18045 9946 18046
rect 9918 18019 9919 18045
rect 9919 18019 9945 18045
rect 9945 18019 9946 18045
rect 9918 18018 9946 18019
rect 9970 18045 9998 18046
rect 9970 18019 9971 18045
rect 9971 18019 9997 18045
rect 9997 18019 9998 18045
rect 9970 18018 9998 18019
rect 10022 18045 10050 18046
rect 10022 18019 10023 18045
rect 10023 18019 10049 18045
rect 10049 18019 10050 18045
rect 10022 18018 10050 18019
rect 9918 17261 9946 17262
rect 9918 17235 9919 17261
rect 9919 17235 9945 17261
rect 9945 17235 9946 17261
rect 9918 17234 9946 17235
rect 9970 17261 9998 17262
rect 9970 17235 9971 17261
rect 9971 17235 9997 17261
rect 9997 17235 9998 17261
rect 9970 17234 9998 17235
rect 10022 17261 10050 17262
rect 10022 17235 10023 17261
rect 10023 17235 10049 17261
rect 10049 17235 10050 17261
rect 10022 17234 10050 17235
rect 9918 16477 9946 16478
rect 9918 16451 9919 16477
rect 9919 16451 9945 16477
rect 9945 16451 9946 16477
rect 9918 16450 9946 16451
rect 9970 16477 9998 16478
rect 9970 16451 9971 16477
rect 9971 16451 9997 16477
rect 9997 16451 9998 16477
rect 9970 16450 9998 16451
rect 10022 16477 10050 16478
rect 10022 16451 10023 16477
rect 10023 16451 10049 16477
rect 10049 16451 10050 16477
rect 10022 16450 10050 16451
rect 8750 13398 8778 13426
rect 9310 13481 9338 13482
rect 9310 13455 9311 13481
rect 9311 13455 9337 13481
rect 9337 13455 9338 13481
rect 9310 13454 9338 13455
rect 8302 13230 8330 13258
rect 9086 13398 9114 13426
rect 9142 13230 9170 13258
rect 8806 12809 8834 12810
rect 8806 12783 8807 12809
rect 8807 12783 8833 12809
rect 8833 12783 8834 12809
rect 8806 12782 8834 12783
rect 6902 11942 6930 11970
rect 7574 11942 7602 11970
rect 7406 11577 7434 11578
rect 7406 11551 7407 11577
rect 7407 11551 7433 11577
rect 7433 11551 7434 11577
rect 7406 11550 7434 11551
rect 7238 11494 7266 11522
rect 2238 11381 2266 11382
rect 2238 11355 2239 11381
rect 2239 11355 2265 11381
rect 2265 11355 2266 11381
rect 2238 11354 2266 11355
rect 2290 11381 2318 11382
rect 2290 11355 2291 11381
rect 2291 11355 2317 11381
rect 2317 11355 2318 11381
rect 2290 11354 2318 11355
rect 2342 11381 2370 11382
rect 2342 11355 2343 11381
rect 2343 11355 2369 11381
rect 2369 11355 2370 11381
rect 2342 11354 2370 11355
rect 7350 11438 7378 11466
rect 5614 11046 5642 11074
rect 6902 11073 6930 11074
rect 6902 11047 6903 11073
rect 6903 11047 6929 11073
rect 6929 11047 6930 11073
rect 6902 11046 6930 11047
rect 7574 11550 7602 11578
rect 7686 11521 7714 11522
rect 7686 11495 7687 11521
rect 7687 11495 7713 11521
rect 7713 11495 7714 11521
rect 7686 11494 7714 11495
rect 7630 11158 7658 11186
rect 7406 11046 7434 11074
rect 7574 11073 7602 11074
rect 7574 11047 7575 11073
rect 7575 11047 7601 11073
rect 7601 11047 7602 11073
rect 7574 11046 7602 11047
rect 7014 10766 7042 10794
rect 2238 10597 2266 10598
rect 2238 10571 2239 10597
rect 2239 10571 2265 10597
rect 2265 10571 2266 10597
rect 2238 10570 2266 10571
rect 2290 10597 2318 10598
rect 2290 10571 2291 10597
rect 2291 10571 2317 10597
rect 2317 10571 2318 10597
rect 2290 10570 2318 10571
rect 2342 10597 2370 10598
rect 2342 10571 2343 10597
rect 2343 10571 2369 10597
rect 2369 10571 2370 10597
rect 2342 10570 2370 10571
rect 6398 10710 6426 10738
rect 7182 10737 7210 10738
rect 7182 10711 7183 10737
rect 7183 10711 7209 10737
rect 7209 10711 7210 10737
rect 7182 10710 7210 10711
rect 2238 9813 2266 9814
rect 2238 9787 2239 9813
rect 2239 9787 2265 9813
rect 2265 9787 2266 9813
rect 2238 9786 2266 9787
rect 2290 9813 2318 9814
rect 2290 9787 2291 9813
rect 2291 9787 2317 9813
rect 2317 9787 2318 9813
rect 2290 9786 2318 9787
rect 2342 9813 2370 9814
rect 2342 9787 2343 9813
rect 2343 9787 2369 9813
rect 2369 9787 2370 9813
rect 2342 9786 2370 9787
rect 7350 9534 7378 9562
rect 2086 9478 2114 9506
rect 6566 9225 6594 9226
rect 6566 9199 6567 9225
rect 6567 9199 6593 9225
rect 6593 9199 6594 9225
rect 6566 9198 6594 9199
rect 6230 9142 6258 9170
rect 2238 9029 2266 9030
rect 2238 9003 2239 9029
rect 2239 9003 2265 9029
rect 2265 9003 2266 9029
rect 2238 9002 2266 9003
rect 2290 9029 2318 9030
rect 2290 9003 2291 9029
rect 2291 9003 2317 9029
rect 2317 9003 2318 9029
rect 2290 9002 2318 9003
rect 2342 9029 2370 9030
rect 2342 9003 2343 9029
rect 2343 9003 2369 9029
rect 2369 9003 2370 9029
rect 2342 9002 2370 9003
rect 7462 10710 7490 10738
rect 7798 11158 7826 11186
rect 7966 11969 7994 11970
rect 7966 11943 7967 11969
rect 7967 11943 7993 11969
rect 7993 11943 7994 11969
rect 7966 11942 7994 11943
rect 8750 12054 8778 12082
rect 8414 11942 8442 11970
rect 8134 11689 8162 11690
rect 8134 11663 8135 11689
rect 8135 11663 8161 11689
rect 8161 11663 8162 11689
rect 8134 11662 8162 11663
rect 8302 11606 8330 11634
rect 7854 10990 7882 11018
rect 7910 11046 7938 11074
rect 7854 10793 7882 10794
rect 7854 10767 7855 10793
rect 7855 10767 7881 10793
rect 7881 10767 7882 10793
rect 7854 10766 7882 10767
rect 7742 10710 7770 10738
rect 8078 11129 8106 11130
rect 8078 11103 8079 11129
rect 8079 11103 8105 11129
rect 8105 11103 8106 11129
rect 8078 11102 8106 11103
rect 9918 15693 9946 15694
rect 9918 15667 9919 15693
rect 9919 15667 9945 15693
rect 9945 15667 9946 15693
rect 9918 15666 9946 15667
rect 9970 15693 9998 15694
rect 9970 15667 9971 15693
rect 9971 15667 9997 15693
rect 9997 15667 9998 15693
rect 9970 15666 9998 15667
rect 10022 15693 10050 15694
rect 10022 15667 10023 15693
rect 10023 15667 10049 15693
rect 10049 15667 10050 15693
rect 10022 15666 10050 15667
rect 9918 14909 9946 14910
rect 9918 14883 9919 14909
rect 9919 14883 9945 14909
rect 9945 14883 9946 14909
rect 9918 14882 9946 14883
rect 9970 14909 9998 14910
rect 9970 14883 9971 14909
rect 9971 14883 9997 14909
rect 9997 14883 9998 14909
rect 9970 14882 9998 14883
rect 10022 14909 10050 14910
rect 10022 14883 10023 14909
rect 10023 14883 10049 14909
rect 10049 14883 10050 14909
rect 10022 14882 10050 14883
rect 9918 14125 9946 14126
rect 9918 14099 9919 14125
rect 9919 14099 9945 14125
rect 9945 14099 9946 14125
rect 9918 14098 9946 14099
rect 9970 14125 9998 14126
rect 9970 14099 9971 14125
rect 9971 14099 9997 14125
rect 9997 14099 9998 14125
rect 9970 14098 9998 14099
rect 10022 14125 10050 14126
rect 10022 14099 10023 14125
rect 10023 14099 10049 14125
rect 10049 14099 10050 14125
rect 10022 14098 10050 14099
rect 10710 13873 10738 13874
rect 10710 13847 10711 13873
rect 10711 13847 10737 13873
rect 10737 13847 10738 13873
rect 10710 13846 10738 13847
rect 9646 13566 9674 13594
rect 9534 13454 9562 13482
rect 9478 12081 9506 12082
rect 9478 12055 9479 12081
rect 9479 12055 9505 12081
rect 9505 12055 9506 12081
rect 9478 12054 9506 12055
rect 8862 11942 8890 11970
rect 9086 11830 9114 11858
rect 8862 11438 8890 11466
rect 8974 11382 9002 11410
rect 9030 11297 9058 11298
rect 9030 11271 9031 11297
rect 9031 11271 9057 11297
rect 9057 11271 9058 11297
rect 9030 11270 9058 11271
rect 9142 11633 9170 11634
rect 9142 11607 9143 11633
rect 9143 11607 9169 11633
rect 9169 11607 9170 11633
rect 9142 11606 9170 11607
rect 9254 11465 9282 11466
rect 9254 11439 9255 11465
rect 9255 11439 9281 11465
rect 9281 11439 9282 11465
rect 9254 11438 9282 11439
rect 9142 11382 9170 11410
rect 8974 11129 9002 11130
rect 8974 11103 8975 11129
rect 8975 11103 9001 11129
rect 9001 11103 9002 11129
rect 8974 11102 9002 11103
rect 7518 9982 7546 10010
rect 7910 9366 7938 9394
rect 7630 9310 7658 9338
rect 7742 9225 7770 9226
rect 7742 9199 7743 9225
rect 7743 9199 7769 9225
rect 7769 9199 7770 9225
rect 7742 9198 7770 9199
rect 7798 9142 7826 9170
rect 7406 8750 7434 8778
rect 7630 8862 7658 8890
rect 7742 8833 7770 8834
rect 7742 8807 7743 8833
rect 7743 8807 7769 8833
rect 7769 8807 7770 8833
rect 7742 8806 7770 8807
rect 8022 9310 8050 9338
rect 8078 9198 8106 9226
rect 8190 10038 8218 10066
rect 8246 10654 8274 10682
rect 8190 9590 8218 9618
rect 8134 9142 8162 9170
rect 8358 10318 8386 10346
rect 8694 10065 8722 10066
rect 8694 10039 8695 10065
rect 8695 10039 8721 10065
rect 8721 10039 8722 10065
rect 8694 10038 8722 10039
rect 8470 9617 8498 9618
rect 8470 9591 8471 9617
rect 8471 9591 8497 9617
rect 8497 9591 8498 9617
rect 8470 9590 8498 9591
rect 8806 9590 8834 9618
rect 8078 8862 8106 8890
rect 8806 9225 8834 9226
rect 8806 9199 8807 9225
rect 8807 9199 8833 9225
rect 8833 9199 8834 9225
rect 8806 9198 8834 9199
rect 8974 9617 9002 9618
rect 8974 9591 8975 9617
rect 8975 9591 9001 9617
rect 9001 9591 9002 9617
rect 8974 9590 9002 9591
rect 9918 13341 9946 13342
rect 9918 13315 9919 13341
rect 9919 13315 9945 13341
rect 9945 13315 9946 13341
rect 9918 13314 9946 13315
rect 9970 13341 9998 13342
rect 9970 13315 9971 13341
rect 9971 13315 9997 13341
rect 9997 13315 9998 13341
rect 9970 13314 9998 13315
rect 10022 13341 10050 13342
rect 10022 13315 10023 13341
rect 10023 13315 10049 13341
rect 10049 13315 10050 13341
rect 10022 13314 10050 13315
rect 9646 13257 9674 13258
rect 9646 13231 9647 13257
rect 9647 13231 9673 13257
rect 9673 13231 9674 13257
rect 9646 13230 9674 13231
rect 9758 13145 9786 13146
rect 9758 13119 9759 13145
rect 9759 13119 9785 13145
rect 9785 13119 9786 13145
rect 9758 13118 9786 13119
rect 10094 13118 10122 13146
rect 9918 12557 9946 12558
rect 9918 12531 9919 12557
rect 9919 12531 9945 12557
rect 9945 12531 9946 12557
rect 9918 12530 9946 12531
rect 9970 12557 9998 12558
rect 9970 12531 9971 12557
rect 9971 12531 9997 12557
rect 9997 12531 9998 12557
rect 9970 12530 9998 12531
rect 10022 12557 10050 12558
rect 10022 12531 10023 12557
rect 10023 12531 10049 12557
rect 10049 12531 10050 12557
rect 10022 12530 10050 12531
rect 9814 12054 9842 12082
rect 9366 11774 9394 11802
rect 9982 11969 10010 11970
rect 9982 11943 9983 11969
rect 9983 11943 10009 11969
rect 10009 11943 10010 11969
rect 9982 11942 10010 11943
rect 10094 11830 10122 11858
rect 9646 11550 9674 11578
rect 9198 11102 9226 11130
rect 9142 10430 9170 10458
rect 9478 10934 9506 10962
rect 9422 10822 9450 10850
rect 9030 9198 9058 9226
rect 8582 8862 8610 8890
rect 8974 8862 9002 8890
rect 8134 8833 8162 8834
rect 8134 8807 8135 8833
rect 8135 8807 8161 8833
rect 8161 8807 8162 8833
rect 8134 8806 8162 8807
rect 8862 8777 8890 8778
rect 8862 8751 8863 8777
rect 8863 8751 8889 8777
rect 8889 8751 8890 8777
rect 8862 8750 8890 8751
rect 7686 8302 7714 8330
rect 2238 8245 2266 8246
rect 2238 8219 2239 8245
rect 2239 8219 2265 8245
rect 2265 8219 2266 8245
rect 2238 8218 2266 8219
rect 2290 8245 2318 8246
rect 2290 8219 2291 8245
rect 2291 8219 2317 8245
rect 2317 8219 2318 8245
rect 2290 8218 2318 8219
rect 2342 8245 2370 8246
rect 2342 8219 2343 8245
rect 2343 8219 2369 8245
rect 2369 8219 2370 8245
rect 2342 8218 2370 8219
rect 7630 8078 7658 8106
rect 2142 8049 2170 8050
rect 2142 8023 2143 8049
rect 2143 8023 2169 8049
rect 2169 8023 2170 8049
rect 2142 8022 2170 8023
rect 6062 8022 6090 8050
rect 966 7742 994 7770
rect 7126 7910 7154 7938
rect 7686 8022 7714 8050
rect 8078 8078 8106 8106
rect 8134 8694 8162 8722
rect 9814 11774 9842 11802
rect 9918 11773 9946 11774
rect 9918 11747 9919 11773
rect 9919 11747 9945 11773
rect 9945 11747 9946 11773
rect 9918 11746 9946 11747
rect 9970 11773 9998 11774
rect 9970 11747 9971 11773
rect 9971 11747 9997 11773
rect 9997 11747 9998 11773
rect 9970 11746 9998 11747
rect 10022 11773 10050 11774
rect 10022 11747 10023 11773
rect 10023 11747 10049 11773
rect 10049 11747 10050 11773
rect 10022 11746 10050 11747
rect 9758 11662 9786 11690
rect 9870 11129 9898 11130
rect 9870 11103 9871 11129
rect 9871 11103 9897 11129
rect 9897 11103 9898 11129
rect 9870 11102 9898 11103
rect 9646 10934 9674 10962
rect 9534 10430 9562 10458
rect 9646 10737 9674 10738
rect 9646 10711 9647 10737
rect 9647 10711 9673 10737
rect 9673 10711 9674 10737
rect 9646 10710 9674 10711
rect 9646 10262 9674 10290
rect 9534 10065 9562 10066
rect 9534 10039 9535 10065
rect 9535 10039 9561 10065
rect 9561 10039 9562 10065
rect 9534 10038 9562 10039
rect 9918 10989 9946 10990
rect 9814 10934 9842 10962
rect 9918 10963 9919 10989
rect 9919 10963 9945 10989
rect 9945 10963 9946 10989
rect 9918 10962 9946 10963
rect 9970 10989 9998 10990
rect 9970 10963 9971 10989
rect 9971 10963 9997 10989
rect 9997 10963 9998 10989
rect 9970 10962 9998 10963
rect 10022 10989 10050 10990
rect 10022 10963 10023 10989
rect 10023 10963 10049 10989
rect 10049 10963 10050 10989
rect 10022 10962 10050 10963
rect 10710 13593 10738 13594
rect 10710 13567 10711 13593
rect 10711 13567 10737 13593
rect 10737 13567 10738 13593
rect 10710 13566 10738 13567
rect 10766 13481 10794 13482
rect 10766 13455 10767 13481
rect 10767 13455 10793 13481
rect 10793 13455 10794 13481
rect 10766 13454 10794 13455
rect 10654 13398 10682 13426
rect 11382 18745 11410 18746
rect 11382 18719 11383 18745
rect 11383 18719 11409 18745
rect 11409 18719 11410 18745
rect 11382 18718 11410 18719
rect 10934 13929 10962 13930
rect 10934 13903 10935 13929
rect 10935 13903 10961 13929
rect 10961 13903 10962 13929
rect 10934 13902 10962 13903
rect 13062 19137 13090 19138
rect 13062 19111 13063 19137
rect 13063 19111 13089 19137
rect 13089 19111 13090 19137
rect 13062 19110 13090 19111
rect 17598 19221 17626 19222
rect 17598 19195 17599 19221
rect 17599 19195 17625 19221
rect 17625 19195 17626 19221
rect 17598 19194 17626 19195
rect 17650 19221 17678 19222
rect 17650 19195 17651 19221
rect 17651 19195 17677 19221
rect 17677 19195 17678 19221
rect 17650 19194 17678 19195
rect 17702 19221 17730 19222
rect 17702 19195 17703 19221
rect 17703 19195 17729 19221
rect 17729 19195 17730 19221
rect 17702 19194 17730 19195
rect 12782 18718 12810 18746
rect 13398 18745 13426 18746
rect 13398 18719 13399 18745
rect 13399 18719 13425 18745
rect 13425 18719 13426 18745
rect 13398 18718 13426 18719
rect 11494 13902 11522 13930
rect 11102 13846 11130 13874
rect 10878 13201 10906 13202
rect 10878 13175 10879 13201
rect 10879 13175 10905 13201
rect 10905 13175 10906 13201
rect 10878 13174 10906 13175
rect 11270 13230 11298 13258
rect 11214 13118 11242 13146
rect 11998 13790 12026 13818
rect 11662 13398 11690 13426
rect 11886 13286 11914 13314
rect 11718 13257 11746 13258
rect 11718 13231 11719 13257
rect 11719 13231 11745 13257
rect 11745 13231 11746 13257
rect 11718 13230 11746 13231
rect 10878 11857 10906 11858
rect 10878 11831 10879 11857
rect 10879 11831 10905 11857
rect 10905 11831 10906 11857
rect 10878 11830 10906 11831
rect 10822 11662 10850 11690
rect 10878 11606 10906 11634
rect 10822 11521 10850 11522
rect 10822 11495 10823 11521
rect 10823 11495 10849 11521
rect 10849 11495 10850 11521
rect 10822 11494 10850 11495
rect 10654 11102 10682 11130
rect 9926 10849 9954 10850
rect 9926 10823 9927 10849
rect 9927 10823 9953 10849
rect 9953 10823 9954 10849
rect 9926 10822 9954 10823
rect 10598 10849 10626 10850
rect 10598 10823 10599 10849
rect 10599 10823 10625 10849
rect 10625 10823 10626 10849
rect 10598 10822 10626 10823
rect 10038 10401 10066 10402
rect 10038 10375 10039 10401
rect 10039 10375 10065 10401
rect 10065 10375 10066 10401
rect 10038 10374 10066 10375
rect 10150 10262 10178 10290
rect 9918 10205 9946 10206
rect 9918 10179 9919 10205
rect 9919 10179 9945 10205
rect 9945 10179 9946 10205
rect 9918 10178 9946 10179
rect 9970 10205 9998 10206
rect 9970 10179 9971 10205
rect 9971 10179 9997 10205
rect 9997 10179 9998 10205
rect 9970 10178 9998 10179
rect 10022 10205 10050 10206
rect 10022 10179 10023 10205
rect 10023 10179 10049 10205
rect 10049 10179 10050 10205
rect 10022 10178 10050 10179
rect 9814 9926 9842 9954
rect 9422 9478 9450 9506
rect 9478 9422 9506 9450
rect 9310 9198 9338 9226
rect 9366 9142 9394 9170
rect 9254 8974 9282 9002
rect 9310 9030 9338 9058
rect 9198 8889 9226 8890
rect 9198 8863 9199 8889
rect 9199 8863 9225 8889
rect 9225 8863 9226 8889
rect 9198 8862 9226 8863
rect 8190 8302 8218 8330
rect 8974 8329 9002 8330
rect 8974 8303 8975 8329
rect 8975 8303 9001 8329
rect 9001 8303 9002 8329
rect 8974 8302 9002 8303
rect 7686 7686 7714 7714
rect 6734 7574 6762 7602
rect 2238 7461 2266 7462
rect 2238 7435 2239 7461
rect 2239 7435 2265 7461
rect 2265 7435 2266 7461
rect 2238 7434 2266 7435
rect 2290 7461 2318 7462
rect 2290 7435 2291 7461
rect 2291 7435 2317 7461
rect 2317 7435 2318 7461
rect 2290 7434 2318 7435
rect 2342 7461 2370 7462
rect 2342 7435 2343 7461
rect 2343 7435 2369 7461
rect 2369 7435 2370 7461
rect 2342 7434 2370 7435
rect 7518 7574 7546 7602
rect 7686 7462 7714 7490
rect 6958 6734 6986 6762
rect 2238 6677 2266 6678
rect 2238 6651 2239 6677
rect 2239 6651 2265 6677
rect 2265 6651 2266 6677
rect 2238 6650 2266 6651
rect 2290 6677 2318 6678
rect 2290 6651 2291 6677
rect 2291 6651 2317 6677
rect 2317 6651 2318 6677
rect 2290 6650 2318 6651
rect 2342 6677 2370 6678
rect 2342 6651 2343 6677
rect 2343 6651 2369 6677
rect 2369 6651 2370 6677
rect 2342 6650 2370 6651
rect 8078 7937 8106 7938
rect 8078 7911 8079 7937
rect 8079 7911 8105 7937
rect 8105 7911 8106 7937
rect 8078 7910 8106 7911
rect 8246 7630 8274 7658
rect 7966 7321 7994 7322
rect 7966 7295 7967 7321
rect 7967 7295 7993 7321
rect 7993 7295 7994 7321
rect 7966 7294 7994 7295
rect 9534 9086 9562 9114
rect 9478 8974 9506 9002
rect 9478 8694 9506 8722
rect 9814 9478 9842 9506
rect 10374 10681 10402 10682
rect 10374 10655 10375 10681
rect 10375 10655 10401 10681
rect 10401 10655 10402 10681
rect 10374 10654 10402 10655
rect 10206 9590 10234 9618
rect 9918 9421 9946 9422
rect 9918 9395 9919 9421
rect 9919 9395 9945 9421
rect 9945 9395 9946 9421
rect 9918 9394 9946 9395
rect 9970 9421 9998 9422
rect 9970 9395 9971 9421
rect 9971 9395 9997 9421
rect 9997 9395 9998 9421
rect 9970 9394 9998 9395
rect 10022 9421 10050 9422
rect 10022 9395 10023 9421
rect 10023 9395 10049 9421
rect 10049 9395 10050 9421
rect 10022 9394 10050 9395
rect 10038 9281 10066 9282
rect 10038 9255 10039 9281
rect 10039 9255 10065 9281
rect 10065 9255 10066 9281
rect 10038 9254 10066 9255
rect 9702 9198 9730 9226
rect 9646 9030 9674 9058
rect 10766 10934 10794 10962
rect 10654 10430 10682 10458
rect 10262 9310 10290 9338
rect 10262 9113 10290 9114
rect 10262 9087 10263 9113
rect 10263 9087 10289 9113
rect 10289 9087 10290 9113
rect 10262 9086 10290 9087
rect 9702 8329 9730 8330
rect 9702 8303 9703 8329
rect 9703 8303 9729 8329
rect 9729 8303 9730 8329
rect 9702 8302 9730 8303
rect 8862 7574 8890 7602
rect 8806 7294 8834 7322
rect 8806 6958 8834 6986
rect 7798 6510 7826 6538
rect 8246 6761 8274 6762
rect 8246 6735 8247 6761
rect 8247 6735 8273 6761
rect 8273 6735 8274 6761
rect 8246 6734 8274 6735
rect 8190 6537 8218 6538
rect 8190 6511 8191 6537
rect 8191 6511 8217 6537
rect 8217 6511 8218 6537
rect 8190 6510 8218 6511
rect 8750 6510 8778 6538
rect 2238 5893 2266 5894
rect 2238 5867 2239 5893
rect 2239 5867 2265 5893
rect 2265 5867 2266 5893
rect 2238 5866 2266 5867
rect 2290 5893 2318 5894
rect 2290 5867 2291 5893
rect 2291 5867 2317 5893
rect 2317 5867 2318 5893
rect 2290 5866 2318 5867
rect 2342 5893 2370 5894
rect 2342 5867 2343 5893
rect 2343 5867 2369 5893
rect 2369 5867 2370 5893
rect 2342 5866 2370 5867
rect 2238 5109 2266 5110
rect 2238 5083 2239 5109
rect 2239 5083 2265 5109
rect 2265 5083 2266 5109
rect 2238 5082 2266 5083
rect 2290 5109 2318 5110
rect 2290 5083 2291 5109
rect 2291 5083 2317 5109
rect 2317 5083 2318 5109
rect 2290 5082 2318 5083
rect 2342 5109 2370 5110
rect 2342 5083 2343 5109
rect 2343 5083 2369 5109
rect 2369 5083 2370 5109
rect 2342 5082 2370 5083
rect 2238 4325 2266 4326
rect 2238 4299 2239 4325
rect 2239 4299 2265 4325
rect 2265 4299 2266 4325
rect 2238 4298 2266 4299
rect 2290 4325 2318 4326
rect 2290 4299 2291 4325
rect 2291 4299 2317 4325
rect 2317 4299 2318 4325
rect 2290 4298 2318 4299
rect 2342 4325 2370 4326
rect 2342 4299 2343 4325
rect 2343 4299 2369 4325
rect 2369 4299 2370 4325
rect 2342 4298 2370 4299
rect 2238 3541 2266 3542
rect 2238 3515 2239 3541
rect 2239 3515 2265 3541
rect 2265 3515 2266 3541
rect 2238 3514 2266 3515
rect 2290 3541 2318 3542
rect 2290 3515 2291 3541
rect 2291 3515 2317 3541
rect 2317 3515 2318 3541
rect 2290 3514 2318 3515
rect 2342 3541 2370 3542
rect 2342 3515 2343 3541
rect 2343 3515 2369 3541
rect 2369 3515 2370 3541
rect 2342 3514 2370 3515
rect 2238 2757 2266 2758
rect 2238 2731 2239 2757
rect 2239 2731 2265 2757
rect 2265 2731 2266 2757
rect 2238 2730 2266 2731
rect 2290 2757 2318 2758
rect 2290 2731 2291 2757
rect 2291 2731 2317 2757
rect 2317 2731 2318 2757
rect 2290 2730 2318 2731
rect 2342 2757 2370 2758
rect 2342 2731 2343 2757
rect 2343 2731 2369 2757
rect 2369 2731 2370 2757
rect 2342 2730 2370 2731
rect 8078 2590 8106 2618
rect 2238 1973 2266 1974
rect 2238 1947 2239 1973
rect 2239 1947 2265 1973
rect 2265 1947 2266 1973
rect 2238 1946 2266 1947
rect 2290 1973 2318 1974
rect 2290 1947 2291 1973
rect 2291 1947 2317 1973
rect 2317 1947 2318 1973
rect 2290 1946 2318 1947
rect 2342 1973 2370 1974
rect 2342 1947 2343 1973
rect 2343 1947 2369 1973
rect 2369 1947 2370 1973
rect 2342 1946 2370 1947
rect 8694 2617 8722 2618
rect 8694 2591 8695 2617
rect 8695 2591 8721 2617
rect 8721 2591 8722 2617
rect 8694 2590 8722 2591
rect 8974 7657 9002 7658
rect 8974 7631 8975 7657
rect 8975 7631 9001 7657
rect 9001 7631 9002 7657
rect 8974 7630 9002 7631
rect 9366 7657 9394 7658
rect 9366 7631 9367 7657
rect 9367 7631 9393 7657
rect 9393 7631 9394 7657
rect 9366 7630 9394 7631
rect 9590 7630 9618 7658
rect 9086 7574 9114 7602
rect 9142 7126 9170 7154
rect 9030 6985 9058 6986
rect 9030 6959 9031 6985
rect 9031 6959 9057 6985
rect 9057 6959 9058 6985
rect 9030 6958 9058 6959
rect 9926 8833 9954 8834
rect 9926 8807 9927 8833
rect 9927 8807 9953 8833
rect 9953 8807 9954 8833
rect 9926 8806 9954 8807
rect 10094 8721 10122 8722
rect 10094 8695 10095 8721
rect 10095 8695 10121 8721
rect 10121 8695 10122 8721
rect 10094 8694 10122 8695
rect 9918 8637 9946 8638
rect 9918 8611 9919 8637
rect 9919 8611 9945 8637
rect 9945 8611 9946 8637
rect 9918 8610 9946 8611
rect 9970 8637 9998 8638
rect 9970 8611 9971 8637
rect 9971 8611 9997 8637
rect 9997 8611 9998 8637
rect 9970 8610 9998 8611
rect 10022 8637 10050 8638
rect 10022 8611 10023 8637
rect 10023 8611 10049 8637
rect 10049 8611 10050 8637
rect 10022 8610 10050 8611
rect 10262 8833 10290 8834
rect 10262 8807 10263 8833
rect 10263 8807 10289 8833
rect 10289 8807 10290 8833
rect 10262 8806 10290 8807
rect 10150 8358 10178 8386
rect 10094 8302 10122 8330
rect 10598 9254 10626 9282
rect 10654 9225 10682 9226
rect 10654 9199 10655 9225
rect 10655 9199 10681 9225
rect 10681 9199 10682 9225
rect 10654 9198 10682 9199
rect 10598 9169 10626 9170
rect 10598 9143 10599 9169
rect 10599 9143 10625 9169
rect 10625 9143 10626 9169
rect 10598 9142 10626 9143
rect 10374 8862 10402 8890
rect 10654 8862 10682 8890
rect 10710 8806 10738 8834
rect 10430 8358 10458 8386
rect 10094 7910 10122 7938
rect 9918 7853 9946 7854
rect 9918 7827 9919 7853
rect 9919 7827 9945 7853
rect 9945 7827 9946 7853
rect 9918 7826 9946 7827
rect 9970 7853 9998 7854
rect 9970 7827 9971 7853
rect 9971 7827 9997 7853
rect 9997 7827 9998 7853
rect 9970 7826 9998 7827
rect 10022 7853 10050 7854
rect 10022 7827 10023 7853
rect 10023 7827 10049 7853
rect 10049 7827 10050 7853
rect 10022 7826 10050 7827
rect 9814 7574 9842 7602
rect 9870 7686 9898 7714
rect 10318 7742 10346 7770
rect 10654 7937 10682 7938
rect 10654 7911 10655 7937
rect 10655 7911 10681 7937
rect 10681 7911 10682 7937
rect 10654 7910 10682 7911
rect 11326 12025 11354 12026
rect 11326 11999 11327 12025
rect 11327 11999 11353 12025
rect 11353 11999 11354 12025
rect 11326 11998 11354 11999
rect 11550 12054 11578 12082
rect 11774 13201 11802 13202
rect 11774 13175 11775 13201
rect 11775 13175 11801 13201
rect 11801 13175 11802 13201
rect 11774 13174 11802 13175
rect 11886 13118 11914 13146
rect 12166 13342 12194 13370
rect 12670 13817 12698 13818
rect 12670 13791 12671 13817
rect 12671 13791 12697 13817
rect 12697 13791 12698 13817
rect 12670 13790 12698 13791
rect 12614 13342 12642 13370
rect 17598 18437 17626 18438
rect 17598 18411 17599 18437
rect 17599 18411 17625 18437
rect 17625 18411 17626 18437
rect 17598 18410 17626 18411
rect 17650 18437 17678 18438
rect 17650 18411 17651 18437
rect 17651 18411 17677 18437
rect 17677 18411 17678 18437
rect 17650 18410 17678 18411
rect 17702 18437 17730 18438
rect 17702 18411 17703 18437
rect 17703 18411 17729 18437
rect 17729 18411 17730 18437
rect 17702 18410 17730 18411
rect 17598 17653 17626 17654
rect 17598 17627 17599 17653
rect 17599 17627 17625 17653
rect 17625 17627 17626 17653
rect 17598 17626 17626 17627
rect 17650 17653 17678 17654
rect 17650 17627 17651 17653
rect 17651 17627 17677 17653
rect 17677 17627 17678 17653
rect 17650 17626 17678 17627
rect 17702 17653 17730 17654
rect 17702 17627 17703 17653
rect 17703 17627 17729 17653
rect 17729 17627 17730 17653
rect 17702 17626 17730 17627
rect 17598 16869 17626 16870
rect 17598 16843 17599 16869
rect 17599 16843 17625 16869
rect 17625 16843 17626 16869
rect 17598 16842 17626 16843
rect 17650 16869 17678 16870
rect 17650 16843 17651 16869
rect 17651 16843 17677 16869
rect 17677 16843 17678 16869
rect 17650 16842 17678 16843
rect 17702 16869 17730 16870
rect 17702 16843 17703 16869
rect 17703 16843 17729 16869
rect 17729 16843 17730 16869
rect 17702 16842 17730 16843
rect 17598 16085 17626 16086
rect 17598 16059 17599 16085
rect 17599 16059 17625 16085
rect 17625 16059 17626 16085
rect 17598 16058 17626 16059
rect 17650 16085 17678 16086
rect 17650 16059 17651 16085
rect 17651 16059 17677 16085
rect 17677 16059 17678 16085
rect 17650 16058 17678 16059
rect 17702 16085 17730 16086
rect 17702 16059 17703 16085
rect 17703 16059 17729 16085
rect 17729 16059 17730 16085
rect 17702 16058 17730 16059
rect 17598 15301 17626 15302
rect 17598 15275 17599 15301
rect 17599 15275 17625 15301
rect 17625 15275 17626 15301
rect 17598 15274 17626 15275
rect 17650 15301 17678 15302
rect 17650 15275 17651 15301
rect 17651 15275 17677 15301
rect 17677 15275 17678 15301
rect 17650 15274 17678 15275
rect 17702 15301 17730 15302
rect 17702 15275 17703 15301
rect 17703 15275 17729 15301
rect 17729 15275 17730 15301
rect 17702 15274 17730 15275
rect 17598 14517 17626 14518
rect 17598 14491 17599 14517
rect 17599 14491 17625 14517
rect 17625 14491 17626 14517
rect 17598 14490 17626 14491
rect 17650 14517 17678 14518
rect 17650 14491 17651 14517
rect 17651 14491 17677 14517
rect 17677 14491 17678 14517
rect 17650 14490 17678 14491
rect 17702 14517 17730 14518
rect 17702 14491 17703 14517
rect 17703 14491 17729 14517
rect 17729 14491 17730 14517
rect 17702 14490 17730 14491
rect 13006 13929 13034 13930
rect 13006 13903 13007 13929
rect 13007 13903 13033 13929
rect 13033 13903 13034 13929
rect 13006 13902 13034 13903
rect 12558 13286 12586 13314
rect 12222 13257 12250 13258
rect 12222 13231 12223 13257
rect 12223 13231 12249 13257
rect 12249 13231 12250 13257
rect 12222 13230 12250 13231
rect 17598 13733 17626 13734
rect 17598 13707 17599 13733
rect 17599 13707 17625 13733
rect 17625 13707 17626 13733
rect 17598 13706 17626 13707
rect 17650 13733 17678 13734
rect 17650 13707 17651 13733
rect 17651 13707 17677 13733
rect 17677 13707 17678 13733
rect 17650 13706 17678 13707
rect 17702 13733 17730 13734
rect 17702 13707 17703 13733
rect 17703 13707 17729 13733
rect 17729 13707 17730 13733
rect 17702 13706 17730 13707
rect 12950 13230 12978 13258
rect 12334 13201 12362 13202
rect 12334 13175 12335 13201
rect 12335 13175 12361 13201
rect 12361 13175 12362 13201
rect 12334 13174 12362 13175
rect 12670 13201 12698 13202
rect 12670 13175 12671 13201
rect 12671 13175 12697 13201
rect 12697 13175 12698 13201
rect 12670 13174 12698 13175
rect 12726 13145 12754 13146
rect 12726 13119 12727 13145
rect 12727 13119 12753 13145
rect 12753 13119 12754 13145
rect 12726 13118 12754 13119
rect 17598 12949 17626 12950
rect 17598 12923 17599 12949
rect 17599 12923 17625 12949
rect 17625 12923 17626 12949
rect 17598 12922 17626 12923
rect 17650 12949 17678 12950
rect 17650 12923 17651 12949
rect 17651 12923 17677 12949
rect 17677 12923 17678 12949
rect 17650 12922 17678 12923
rect 17702 12949 17730 12950
rect 17702 12923 17703 12949
rect 17703 12923 17729 12949
rect 17729 12923 17730 12949
rect 17702 12922 17730 12923
rect 12110 12334 12138 12362
rect 11550 11577 11578 11578
rect 11550 11551 11551 11577
rect 11551 11551 11577 11577
rect 11577 11551 11578 11577
rect 11550 11550 11578 11551
rect 11606 11521 11634 11522
rect 11606 11495 11607 11521
rect 11607 11495 11633 11521
rect 11633 11495 11634 11521
rect 11606 11494 11634 11495
rect 11214 11102 11242 11130
rect 11102 10934 11130 10962
rect 10878 10486 10906 10514
rect 11046 10345 11074 10346
rect 11046 10319 11047 10345
rect 11047 10319 11073 10345
rect 11073 10319 11074 10345
rect 11046 10318 11074 10319
rect 10878 10289 10906 10290
rect 10878 10263 10879 10289
rect 10879 10263 10905 10289
rect 10905 10263 10906 10289
rect 10878 10262 10906 10263
rect 11158 10038 11186 10066
rect 11662 11270 11690 11298
rect 11774 11606 11802 11634
rect 11774 11046 11802 11074
rect 11718 10793 11746 10794
rect 11718 10767 11719 10793
rect 11719 10767 11745 10793
rect 11745 10767 11746 10793
rect 11718 10766 11746 10767
rect 11326 10654 11354 10682
rect 11270 10457 11298 10458
rect 11270 10431 11271 10457
rect 11271 10431 11297 10457
rect 11297 10431 11298 10457
rect 11270 10430 11298 10431
rect 11214 9758 11242 9786
rect 10822 9478 10850 9506
rect 10934 9337 10962 9338
rect 10934 9311 10935 9337
rect 10935 9311 10961 9337
rect 10961 9311 10962 9337
rect 10934 9310 10962 9311
rect 10822 8721 10850 8722
rect 10822 8695 10823 8721
rect 10823 8695 10849 8721
rect 10849 8695 10850 8721
rect 10822 8694 10850 8695
rect 10822 7937 10850 7938
rect 10822 7911 10823 7937
rect 10823 7911 10849 7937
rect 10849 7911 10850 7937
rect 10822 7910 10850 7911
rect 10430 7713 10458 7714
rect 10430 7687 10431 7713
rect 10431 7687 10457 7713
rect 10457 7687 10458 7713
rect 10430 7686 10458 7687
rect 10486 7630 10514 7658
rect 10262 7238 10290 7266
rect 10374 7209 10402 7210
rect 10374 7183 10375 7209
rect 10375 7183 10401 7209
rect 10401 7183 10402 7209
rect 10374 7182 10402 7183
rect 9758 7153 9786 7154
rect 9758 7127 9759 7153
rect 9759 7127 9785 7153
rect 9785 7127 9786 7153
rect 9758 7126 9786 7127
rect 9918 7069 9946 7070
rect 9918 7043 9919 7069
rect 9919 7043 9945 7069
rect 9945 7043 9946 7069
rect 9918 7042 9946 7043
rect 9970 7069 9998 7070
rect 9970 7043 9971 7069
rect 9971 7043 9997 7069
rect 9997 7043 9998 7069
rect 9970 7042 9998 7043
rect 10022 7069 10050 7070
rect 10022 7043 10023 7069
rect 10023 7043 10049 7069
rect 10049 7043 10050 7069
rect 10022 7042 10050 7043
rect 10542 7601 10570 7602
rect 10542 7575 10543 7601
rect 10543 7575 10569 7601
rect 10569 7575 10570 7601
rect 10542 7574 10570 7575
rect 10710 7294 10738 7322
rect 11270 10094 11298 10122
rect 12614 12054 12642 12082
rect 12222 11998 12250 12026
rect 12558 11998 12586 12026
rect 12166 11886 12194 11914
rect 12614 11913 12642 11914
rect 12614 11887 12615 11913
rect 12615 11887 12641 11913
rect 12641 11887 12642 11913
rect 12614 11886 12642 11887
rect 12278 11633 12306 11634
rect 12278 11607 12279 11633
rect 12279 11607 12305 11633
rect 12305 11607 12306 11633
rect 12278 11606 12306 11607
rect 12558 11606 12586 11634
rect 11942 11270 11970 11298
rect 12278 11185 12306 11186
rect 12278 11159 12279 11185
rect 12279 11159 12305 11185
rect 12305 11159 12306 11185
rect 12278 11158 12306 11159
rect 12614 11577 12642 11578
rect 12614 11551 12615 11577
rect 12615 11551 12641 11577
rect 12641 11551 12642 11577
rect 12614 11550 12642 11551
rect 12894 12361 12922 12362
rect 12894 12335 12895 12361
rect 12895 12335 12921 12361
rect 12921 12335 12922 12361
rect 12894 12334 12922 12335
rect 17598 12165 17626 12166
rect 17598 12139 17599 12165
rect 17599 12139 17625 12165
rect 17625 12139 17626 12165
rect 17598 12138 17626 12139
rect 17650 12165 17678 12166
rect 17650 12139 17651 12165
rect 17651 12139 17677 12165
rect 17677 12139 17678 12165
rect 17650 12138 17678 12139
rect 17702 12165 17730 12166
rect 17702 12139 17703 12165
rect 17703 12139 17729 12165
rect 17729 12139 17730 12165
rect 17702 12138 17730 12139
rect 13678 12025 13706 12026
rect 13678 11999 13679 12025
rect 13679 11999 13705 12025
rect 13705 11999 13706 12025
rect 13678 11998 13706 11999
rect 13902 11998 13930 12026
rect 18830 11969 18858 11970
rect 18830 11943 18831 11969
rect 18831 11943 18857 11969
rect 18857 11943 18858 11969
rect 18830 11942 18858 11943
rect 14014 11857 14042 11858
rect 14014 11831 14015 11857
rect 14015 11831 14041 11857
rect 14041 11831 14042 11857
rect 14014 11830 14042 11831
rect 20006 12110 20034 12138
rect 18942 11830 18970 11858
rect 13678 11606 13706 11634
rect 13174 11550 13202 11578
rect 12446 11073 12474 11074
rect 12446 11047 12447 11073
rect 12447 11047 12473 11073
rect 12473 11047 12474 11073
rect 12446 11046 12474 11047
rect 11830 10934 11858 10962
rect 20006 11774 20034 11802
rect 14294 11577 14322 11578
rect 14294 11551 14295 11577
rect 14295 11551 14321 11577
rect 14321 11551 14322 11577
rect 14294 11550 14322 11551
rect 18830 11577 18858 11578
rect 18830 11551 18831 11577
rect 18831 11551 18857 11577
rect 18857 11551 18858 11577
rect 18830 11550 18858 11551
rect 13230 11494 13258 11522
rect 14070 11521 14098 11522
rect 14070 11495 14071 11521
rect 14071 11495 14097 11521
rect 14097 11495 14098 11521
rect 14070 11494 14098 11495
rect 20006 11465 20034 11466
rect 20006 11439 20007 11465
rect 20007 11439 20033 11465
rect 20033 11439 20034 11465
rect 20006 11438 20034 11439
rect 17598 11381 17626 11382
rect 17598 11355 17599 11381
rect 17599 11355 17625 11381
rect 17625 11355 17626 11381
rect 17598 11354 17626 11355
rect 17650 11381 17678 11382
rect 17650 11355 17651 11381
rect 17651 11355 17677 11381
rect 17677 11355 17678 11381
rect 17650 11354 17678 11355
rect 17702 11381 17730 11382
rect 17702 11355 17703 11381
rect 17703 11355 17729 11381
rect 17729 11355 17730 11381
rect 17702 11354 17730 11355
rect 18830 11185 18858 11186
rect 18830 11159 18831 11185
rect 18831 11159 18857 11185
rect 18857 11159 18858 11185
rect 18830 11158 18858 11159
rect 13286 11129 13314 11130
rect 13286 11103 13287 11129
rect 13287 11103 13313 11129
rect 13313 11103 13314 11129
rect 13286 11102 13314 11103
rect 11438 10318 11466 10346
rect 11662 10401 11690 10402
rect 11662 10375 11663 10401
rect 11663 10375 11689 10401
rect 11689 10375 11690 10401
rect 11662 10374 11690 10375
rect 11886 10486 11914 10514
rect 11998 10094 12026 10122
rect 12166 10793 12194 10794
rect 12166 10767 12167 10793
rect 12167 10767 12193 10793
rect 12193 10767 12194 10793
rect 12166 10766 12194 10767
rect 13174 10766 13202 10794
rect 12110 10038 12138 10066
rect 12558 10038 12586 10066
rect 12614 10094 12642 10122
rect 12334 9982 12362 10010
rect 12894 10094 12922 10122
rect 12670 10065 12698 10066
rect 12670 10039 12671 10065
rect 12671 10039 12697 10065
rect 12697 10039 12698 10065
rect 12670 10038 12698 10039
rect 11718 9534 11746 9562
rect 11046 8694 11074 8722
rect 12726 9142 12754 9170
rect 13174 10094 13202 10122
rect 13342 10094 13370 10122
rect 13678 10793 13706 10794
rect 13678 10767 13679 10793
rect 13679 10767 13705 10793
rect 13705 10767 13706 10793
rect 13678 10766 13706 10767
rect 20006 11102 20034 11130
rect 14910 11073 14938 11074
rect 14910 11047 14911 11073
rect 14911 11047 14937 11073
rect 14937 11047 14938 11073
rect 14910 11046 14938 11047
rect 14742 10710 14770 10738
rect 15134 10737 15162 10738
rect 15134 10711 15135 10737
rect 15135 10711 15161 10737
rect 15161 10711 15162 10737
rect 15134 10710 15162 10711
rect 14238 10486 14266 10514
rect 14574 10513 14602 10514
rect 14574 10487 14575 10513
rect 14575 10487 14601 10513
rect 14601 10487 14602 10513
rect 14574 10486 14602 10487
rect 13454 10430 13482 10458
rect 14854 10345 14882 10346
rect 14854 10319 14855 10345
rect 14855 10319 14881 10345
rect 14881 10319 14882 10345
rect 14854 10318 14882 10319
rect 14518 10094 14546 10122
rect 13230 9561 13258 9562
rect 13230 9535 13231 9561
rect 13231 9535 13257 9561
rect 13257 9535 13258 9561
rect 13230 9534 13258 9535
rect 13286 9254 13314 9282
rect 11326 9086 11354 9114
rect 11662 8694 11690 8722
rect 11550 7993 11578 7994
rect 11550 7967 11551 7993
rect 11551 7967 11577 7993
rect 11577 7967 11578 7993
rect 11550 7966 11578 7967
rect 11438 7742 11466 7770
rect 10934 7657 10962 7658
rect 10934 7631 10935 7657
rect 10935 7631 10961 7657
rect 10961 7631 10962 7657
rect 10934 7630 10962 7631
rect 11046 7321 11074 7322
rect 11046 7295 11047 7321
rect 11047 7295 11073 7321
rect 11073 7295 11074 7321
rect 11046 7294 11074 7295
rect 10990 7265 11018 7266
rect 10990 7239 10991 7265
rect 10991 7239 11017 7265
rect 11017 7239 11018 7265
rect 10990 7238 11018 7239
rect 11214 7209 11242 7210
rect 11214 7183 11215 7209
rect 11215 7183 11241 7209
rect 11241 7183 11242 7209
rect 11214 7182 11242 7183
rect 11942 7993 11970 7994
rect 11942 7967 11943 7993
rect 11943 7967 11969 7993
rect 11969 7967 11970 7993
rect 11942 7966 11970 7967
rect 11998 7937 12026 7938
rect 11998 7911 11999 7937
rect 11999 7911 12025 7937
rect 12025 7911 12026 7937
rect 11998 7910 12026 7911
rect 11662 7182 11690 7210
rect 12110 7518 12138 7546
rect 9534 6510 9562 6538
rect 11102 6790 11130 6818
rect 11886 6817 11914 6818
rect 11886 6791 11887 6817
rect 11887 6791 11913 6817
rect 11913 6791 11914 6817
rect 11886 6790 11914 6791
rect 10374 6537 10402 6538
rect 10374 6511 10375 6537
rect 10375 6511 10401 6537
rect 10401 6511 10402 6537
rect 10374 6510 10402 6511
rect 9918 6285 9946 6286
rect 9918 6259 9919 6285
rect 9919 6259 9945 6285
rect 9945 6259 9946 6285
rect 9918 6258 9946 6259
rect 9970 6285 9998 6286
rect 9970 6259 9971 6285
rect 9971 6259 9997 6285
rect 9997 6259 9998 6285
rect 9970 6258 9998 6259
rect 10022 6285 10050 6286
rect 10022 6259 10023 6285
rect 10023 6259 10049 6285
rect 10049 6259 10050 6285
rect 10022 6258 10050 6259
rect 9918 5501 9946 5502
rect 9918 5475 9919 5501
rect 9919 5475 9945 5501
rect 9945 5475 9946 5501
rect 9918 5474 9946 5475
rect 9970 5501 9998 5502
rect 9970 5475 9971 5501
rect 9971 5475 9997 5501
rect 9997 5475 9998 5501
rect 9970 5474 9998 5475
rect 10022 5501 10050 5502
rect 10022 5475 10023 5501
rect 10023 5475 10049 5501
rect 10049 5475 10050 5501
rect 10022 5474 10050 5475
rect 9918 4717 9946 4718
rect 9918 4691 9919 4717
rect 9919 4691 9945 4717
rect 9945 4691 9946 4717
rect 9918 4690 9946 4691
rect 9970 4717 9998 4718
rect 9970 4691 9971 4717
rect 9971 4691 9997 4717
rect 9997 4691 9998 4717
rect 9970 4690 9998 4691
rect 10022 4717 10050 4718
rect 10022 4691 10023 4717
rect 10023 4691 10049 4717
rect 10049 4691 10050 4717
rect 10022 4690 10050 4691
rect 9918 3933 9946 3934
rect 9918 3907 9919 3933
rect 9919 3907 9945 3933
rect 9945 3907 9946 3933
rect 9918 3906 9946 3907
rect 9970 3933 9998 3934
rect 9970 3907 9971 3933
rect 9971 3907 9997 3933
rect 9997 3907 9998 3933
rect 9970 3906 9998 3907
rect 10022 3933 10050 3934
rect 10022 3907 10023 3933
rect 10023 3907 10049 3933
rect 10049 3907 10050 3933
rect 10022 3906 10050 3907
rect 9918 3149 9946 3150
rect 9918 3123 9919 3149
rect 9919 3123 9945 3149
rect 9945 3123 9946 3149
rect 9918 3122 9946 3123
rect 9970 3149 9998 3150
rect 9970 3123 9971 3149
rect 9971 3123 9997 3149
rect 9997 3123 9998 3149
rect 9970 3122 9998 3123
rect 10022 3149 10050 3150
rect 10022 3123 10023 3149
rect 10023 3123 10049 3149
rect 10049 3123 10050 3149
rect 10022 3122 10050 3123
rect 9918 2365 9946 2366
rect 9918 2339 9919 2365
rect 9919 2339 9945 2365
rect 9945 2339 9946 2365
rect 9918 2338 9946 2339
rect 9970 2365 9998 2366
rect 9970 2339 9971 2365
rect 9971 2339 9997 2365
rect 9997 2339 9998 2365
rect 9970 2338 9998 2339
rect 10022 2365 10050 2366
rect 10022 2339 10023 2365
rect 10023 2339 10049 2365
rect 10049 2339 10050 2365
rect 10022 2338 10050 2339
rect 9758 2030 9786 2058
rect 10374 2057 10402 2058
rect 10374 2031 10375 2057
rect 10375 2031 10401 2057
rect 10401 2031 10402 2057
rect 10374 2030 10402 2031
rect 11886 1806 11914 1834
rect 9918 1581 9946 1582
rect 9918 1555 9919 1581
rect 9919 1555 9945 1581
rect 9945 1555 9946 1581
rect 9918 1554 9946 1555
rect 9970 1581 9998 1582
rect 9970 1555 9971 1581
rect 9971 1555 9997 1581
rect 9997 1555 9998 1581
rect 9970 1554 9998 1555
rect 10022 1581 10050 1582
rect 10022 1555 10023 1581
rect 10023 1555 10049 1581
rect 10049 1555 10050 1581
rect 10022 1554 10050 1555
rect 12670 7518 12698 7546
rect 13510 9198 13538 9226
rect 14182 9926 14210 9954
rect 14238 9758 14266 9786
rect 13454 9030 13482 9058
rect 13118 8049 13146 8050
rect 13118 8023 13119 8049
rect 13119 8023 13145 8049
rect 13145 8023 13146 8049
rect 13118 8022 13146 8023
rect 14350 9169 14378 9170
rect 14350 9143 14351 9169
rect 14351 9143 14377 9169
rect 14377 9143 14378 9169
rect 14350 9142 14378 9143
rect 14798 9953 14826 9954
rect 14798 9927 14799 9953
rect 14799 9927 14825 9953
rect 14825 9927 14826 9953
rect 14798 9926 14826 9927
rect 17598 10597 17626 10598
rect 17598 10571 17599 10597
rect 17599 10571 17625 10597
rect 17625 10571 17626 10597
rect 17598 10570 17626 10571
rect 17650 10597 17678 10598
rect 17650 10571 17651 10597
rect 17651 10571 17677 10597
rect 17677 10571 17678 10597
rect 17650 10570 17678 10571
rect 17702 10597 17730 10598
rect 17702 10571 17703 10597
rect 17703 10571 17729 10597
rect 17729 10571 17730 10597
rect 17702 10570 17730 10571
rect 15302 10401 15330 10402
rect 15302 10375 15303 10401
rect 15303 10375 15329 10401
rect 15329 10375 15330 10401
rect 15302 10374 15330 10375
rect 20006 10766 20034 10794
rect 18830 10374 18858 10402
rect 18830 10009 18858 10010
rect 18830 9983 18831 10009
rect 18831 9983 18857 10009
rect 18857 9983 18858 10009
rect 18830 9982 18858 9983
rect 18830 9870 18858 9898
rect 15190 9758 15218 9786
rect 17598 9813 17626 9814
rect 17598 9787 17599 9813
rect 17599 9787 17625 9813
rect 17625 9787 17626 9813
rect 17598 9786 17626 9787
rect 17650 9813 17678 9814
rect 17650 9787 17651 9813
rect 17651 9787 17677 9813
rect 17677 9787 17678 9813
rect 17650 9786 17678 9787
rect 17702 9813 17730 9814
rect 17702 9787 17703 9813
rect 17703 9787 17729 9813
rect 17729 9787 17730 9813
rect 17702 9786 17730 9787
rect 20006 9758 20034 9786
rect 20006 9422 20034 9450
rect 18830 9225 18858 9226
rect 18830 9199 18831 9225
rect 18831 9199 18857 9225
rect 18857 9199 18858 9225
rect 18830 9198 18858 9199
rect 13566 8022 13594 8050
rect 14014 8022 14042 8050
rect 13286 7993 13314 7994
rect 13286 7967 13287 7993
rect 13287 7967 13313 7993
rect 13313 7967 13314 7993
rect 13286 7966 13314 7967
rect 12894 7518 12922 7546
rect 13398 7910 13426 7938
rect 13958 7937 13986 7938
rect 13958 7911 13959 7937
rect 13959 7911 13985 7937
rect 13985 7911 13986 7937
rect 13958 7910 13986 7911
rect 13734 7742 13762 7770
rect 13622 7574 13650 7602
rect 14294 7686 14322 7714
rect 14462 7601 14490 7602
rect 14462 7575 14463 7601
rect 14463 7575 14489 7601
rect 14489 7575 14490 7601
rect 14462 7574 14490 7575
rect 20006 9113 20034 9114
rect 20006 9087 20007 9113
rect 20007 9087 20033 9113
rect 20033 9087 20034 9113
rect 20006 9086 20034 9087
rect 17598 9029 17626 9030
rect 17598 9003 17599 9029
rect 17599 9003 17625 9029
rect 17625 9003 17626 9029
rect 17598 9002 17626 9003
rect 17650 9029 17678 9030
rect 17650 9003 17651 9029
rect 17651 9003 17677 9029
rect 17677 9003 17678 9029
rect 17650 9002 17678 9003
rect 17702 9029 17730 9030
rect 17702 9003 17703 9029
rect 17703 9003 17729 9029
rect 17729 9003 17730 9029
rect 17702 9002 17730 9003
rect 17598 8245 17626 8246
rect 17598 8219 17599 8245
rect 17599 8219 17625 8245
rect 17625 8219 17626 8245
rect 17598 8218 17626 8219
rect 17650 8245 17678 8246
rect 17650 8219 17651 8245
rect 17651 8219 17677 8245
rect 17677 8219 17678 8245
rect 17650 8218 17678 8219
rect 17702 8245 17730 8246
rect 17702 8219 17703 8245
rect 17703 8219 17729 8245
rect 17729 8219 17730 8245
rect 17702 8218 17730 8219
rect 14686 7966 14714 7994
rect 14630 7742 14658 7770
rect 14798 7686 14826 7714
rect 18830 7657 18858 7658
rect 18830 7631 18831 7657
rect 18831 7631 18857 7657
rect 18857 7631 18858 7657
rect 18830 7630 18858 7631
rect 20006 7742 20034 7770
rect 18942 7574 18970 7602
rect 17598 7461 17626 7462
rect 17598 7435 17599 7461
rect 17599 7435 17625 7461
rect 17625 7435 17626 7461
rect 17598 7434 17626 7435
rect 17650 7461 17678 7462
rect 17650 7435 17651 7461
rect 17651 7435 17677 7461
rect 17677 7435 17678 7461
rect 17650 7434 17678 7435
rect 17702 7461 17730 7462
rect 17702 7435 17703 7461
rect 17703 7435 17729 7461
rect 17729 7435 17730 7461
rect 17702 7434 17730 7435
rect 20006 7406 20034 7434
rect 20118 7070 20146 7098
rect 17598 6677 17626 6678
rect 17598 6651 17599 6677
rect 17599 6651 17625 6677
rect 17625 6651 17626 6677
rect 17598 6650 17626 6651
rect 17650 6677 17678 6678
rect 17650 6651 17651 6677
rect 17651 6651 17677 6677
rect 17677 6651 17678 6677
rect 17650 6650 17678 6651
rect 17702 6677 17730 6678
rect 17702 6651 17703 6677
rect 17703 6651 17729 6677
rect 17729 6651 17730 6677
rect 17702 6650 17730 6651
rect 17598 5893 17626 5894
rect 17598 5867 17599 5893
rect 17599 5867 17625 5893
rect 17625 5867 17626 5893
rect 17598 5866 17626 5867
rect 17650 5893 17678 5894
rect 17650 5867 17651 5893
rect 17651 5867 17677 5893
rect 17677 5867 17678 5893
rect 17650 5866 17678 5867
rect 17702 5893 17730 5894
rect 17702 5867 17703 5893
rect 17703 5867 17729 5893
rect 17729 5867 17730 5893
rect 17702 5866 17730 5867
rect 17598 5109 17626 5110
rect 17598 5083 17599 5109
rect 17599 5083 17625 5109
rect 17625 5083 17626 5109
rect 17598 5082 17626 5083
rect 17650 5109 17678 5110
rect 17650 5083 17651 5109
rect 17651 5083 17677 5109
rect 17677 5083 17678 5109
rect 17650 5082 17678 5083
rect 17702 5109 17730 5110
rect 17702 5083 17703 5109
rect 17703 5083 17729 5109
rect 17729 5083 17730 5109
rect 17702 5082 17730 5083
rect 17598 4325 17626 4326
rect 17598 4299 17599 4325
rect 17599 4299 17625 4325
rect 17625 4299 17626 4325
rect 17598 4298 17626 4299
rect 17650 4325 17678 4326
rect 17650 4299 17651 4325
rect 17651 4299 17677 4325
rect 17677 4299 17678 4325
rect 17650 4298 17678 4299
rect 17702 4325 17730 4326
rect 17702 4299 17703 4325
rect 17703 4299 17729 4325
rect 17729 4299 17730 4325
rect 17702 4298 17730 4299
rect 17598 3541 17626 3542
rect 17598 3515 17599 3541
rect 17599 3515 17625 3541
rect 17625 3515 17626 3541
rect 17598 3514 17626 3515
rect 17650 3541 17678 3542
rect 17650 3515 17651 3541
rect 17651 3515 17677 3541
rect 17677 3515 17678 3541
rect 17650 3514 17678 3515
rect 17702 3541 17730 3542
rect 17702 3515 17703 3541
rect 17703 3515 17729 3541
rect 17729 3515 17730 3541
rect 17702 3514 17730 3515
rect 17598 2757 17626 2758
rect 17598 2731 17599 2757
rect 17599 2731 17625 2757
rect 17625 2731 17626 2757
rect 17598 2730 17626 2731
rect 17650 2757 17678 2758
rect 17650 2731 17651 2757
rect 17651 2731 17677 2757
rect 17677 2731 17678 2757
rect 17650 2730 17678 2731
rect 17702 2757 17730 2758
rect 17702 2731 17703 2757
rect 17703 2731 17729 2757
rect 17729 2731 17730 2757
rect 17702 2730 17730 2731
rect 17598 1973 17626 1974
rect 17598 1947 17599 1973
rect 17599 1947 17625 1973
rect 17625 1947 17626 1973
rect 17598 1946 17626 1947
rect 17650 1973 17678 1974
rect 17650 1947 17651 1973
rect 17651 1947 17677 1973
rect 17677 1947 17678 1973
rect 17650 1946 17678 1947
rect 17702 1973 17730 1974
rect 17702 1947 17703 1973
rect 17703 1947 17729 1973
rect 17729 1947 17730 1973
rect 17702 1946 17730 1947
rect 12782 1833 12810 1834
rect 12782 1807 12783 1833
rect 12783 1807 12809 1833
rect 12809 1807 12810 1833
rect 12782 1806 12810 1807
<< metal3 >>
rect 2233 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2375 19222
rect 17593 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17735 19222
rect 12441 19110 12446 19138
rect 12474 19110 13062 19138
rect 13090 19110 13095 19138
rect 9913 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10055 18830
rect 9417 18718 9422 18746
rect 9450 18718 9926 18746
rect 9954 18718 9959 18746
rect 10761 18718 10766 18746
rect 10794 18718 11382 18746
rect 11410 18718 11415 18746
rect 12777 18718 12782 18746
rect 12810 18718 13398 18746
rect 13426 18718 13431 18746
rect 2233 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2375 18438
rect 17593 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17735 18438
rect 8409 18326 8414 18354
rect 8442 18326 9030 18354
rect 9058 18326 9063 18354
rect 9913 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10055 18046
rect 2233 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2375 17654
rect 17593 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17735 17654
rect 9913 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10055 17262
rect 2233 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2375 16870
rect 17593 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17735 16870
rect 9913 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10055 16478
rect 2233 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2375 16086
rect 17593 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17735 16086
rect 9913 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10055 15694
rect 2233 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2375 15302
rect 17593 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17735 15302
rect 9913 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10055 14910
rect 2233 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2375 14518
rect 17593 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17735 14518
rect 9913 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10055 14126
rect 10929 13902 10934 13930
rect 10962 13902 11494 13930
rect 11522 13902 13006 13930
rect 13034 13902 13039 13930
rect 10705 13846 10710 13874
rect 10738 13846 11102 13874
rect 11130 13846 11135 13874
rect 11993 13790 11998 13818
rect 12026 13790 12670 13818
rect 12698 13790 12703 13818
rect 2233 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2375 13734
rect 17593 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17735 13734
rect 9641 13566 9646 13594
rect 9674 13566 10710 13594
rect 10738 13566 10743 13594
rect 0 13482 400 13496
rect 0 13454 2086 13482
rect 2114 13454 2119 13482
rect 9305 13454 9310 13482
rect 9338 13454 9534 13482
rect 9562 13454 10766 13482
rect 10794 13454 10799 13482
rect 0 13440 400 13454
rect 8745 13398 8750 13426
rect 8778 13398 9086 13426
rect 9114 13398 9119 13426
rect 10649 13398 10654 13426
rect 10682 13398 11662 13426
rect 11690 13398 11695 13426
rect 10374 13342 12166 13370
rect 12194 13342 12614 13370
rect 12642 13342 12647 13370
rect 9913 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10055 13342
rect 10374 13258 10402 13342
rect 11881 13286 11886 13314
rect 11914 13286 12558 13314
rect 12586 13286 12591 13314
rect 8297 13230 8302 13258
rect 8330 13230 9142 13258
rect 9170 13230 9646 13258
rect 9674 13230 10402 13258
rect 11265 13230 11270 13258
rect 11298 13230 11718 13258
rect 11746 13230 11751 13258
rect 12217 13230 12222 13258
rect 12250 13230 12950 13258
rect 12978 13230 12983 13258
rect 10873 13174 10878 13202
rect 10906 13174 11774 13202
rect 11802 13174 11807 13202
rect 12329 13174 12334 13202
rect 12362 13174 12670 13202
rect 12698 13174 12703 13202
rect 9753 13118 9758 13146
rect 9786 13118 10094 13146
rect 10122 13118 11214 13146
rect 11242 13118 11247 13146
rect 11881 13118 11886 13146
rect 11914 13118 12726 13146
rect 12754 13118 12759 13146
rect 7233 13062 7238 13090
rect 7266 13062 7630 13090
rect 7658 13062 7663 13090
rect 2233 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2375 12950
rect 17593 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17735 12950
rect 7681 12782 7686 12810
rect 7714 12782 8806 12810
rect 8834 12782 8839 12810
rect 9913 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10055 12558
rect 12105 12334 12110 12362
rect 12138 12334 12894 12362
rect 12922 12334 12927 12362
rect 2233 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2375 12166
rect 17593 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17735 12166
rect 20600 12138 21000 12152
rect 20001 12110 20006 12138
rect 20034 12110 21000 12138
rect 20600 12096 21000 12110
rect 8745 12054 8750 12082
rect 8778 12054 9478 12082
rect 9506 12054 9511 12082
rect 9809 12054 9814 12082
rect 9842 12054 11550 12082
rect 11578 12054 12614 12082
rect 12642 12054 12647 12082
rect 11321 11998 11326 12026
rect 11354 11998 12222 12026
rect 12250 11998 12558 12026
rect 12586 11998 12591 12026
rect 13673 11998 13678 12026
rect 13706 11998 13902 12026
rect 13930 11998 15974 12026
rect 15946 11970 15974 11998
rect 2137 11942 2142 11970
rect 2170 11942 6006 11970
rect 6034 11942 6039 11970
rect 6897 11942 6902 11970
rect 6930 11942 7574 11970
rect 7602 11942 7966 11970
rect 7994 11942 8414 11970
rect 8442 11942 8862 11970
rect 8890 11942 9982 11970
rect 10010 11942 10015 11970
rect 15946 11942 18830 11970
rect 18858 11942 18863 11970
rect 12161 11886 12166 11914
rect 12194 11886 12614 11914
rect 12642 11886 12647 11914
rect 9081 11830 9086 11858
rect 9114 11830 10094 11858
rect 10122 11830 10878 11858
rect 10906 11830 10911 11858
rect 14009 11830 14014 11858
rect 14042 11830 18942 11858
rect 18970 11830 18975 11858
rect 0 11802 400 11816
rect 20600 11802 21000 11816
rect 0 11774 966 11802
rect 994 11774 999 11802
rect 9361 11774 9366 11802
rect 9394 11774 9814 11802
rect 9842 11774 9847 11802
rect 20001 11774 20006 11802
rect 20034 11774 21000 11802
rect 0 11760 400 11774
rect 9913 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10055 11774
rect 20600 11760 21000 11774
rect 6001 11662 6006 11690
rect 6034 11662 8134 11690
rect 8162 11662 8167 11690
rect 9753 11662 9758 11690
rect 9786 11662 10822 11690
rect 10850 11662 10855 11690
rect 8297 11606 8302 11634
rect 8330 11606 9142 11634
rect 9170 11606 9175 11634
rect 10873 11606 10878 11634
rect 10906 11606 11774 11634
rect 11802 11606 12278 11634
rect 12306 11606 12311 11634
rect 12553 11606 12558 11634
rect 12586 11606 13678 11634
rect 13706 11606 13711 11634
rect 7401 11550 7406 11578
rect 7434 11550 7574 11578
rect 7602 11550 7607 11578
rect 9641 11550 9646 11578
rect 9674 11550 11550 11578
rect 11578 11550 11583 11578
rect 12609 11550 12614 11578
rect 12642 11550 13174 11578
rect 13202 11550 14294 11578
rect 14322 11550 14327 11578
rect 15946 11550 18830 11578
rect 18858 11550 18863 11578
rect 15946 11522 15974 11550
rect 7233 11494 7238 11522
rect 7266 11494 7686 11522
rect 7714 11494 7719 11522
rect 10817 11494 10822 11522
rect 10850 11494 11606 11522
rect 11634 11494 11639 11522
rect 13225 11494 13230 11522
rect 13258 11494 14070 11522
rect 14098 11494 15974 11522
rect 20600 11466 21000 11480
rect 7345 11438 7350 11466
rect 7378 11438 8862 11466
rect 8890 11438 9254 11466
rect 9282 11438 9287 11466
rect 20001 11438 20006 11466
rect 20034 11438 21000 11466
rect 20600 11424 21000 11438
rect 8969 11382 8974 11410
rect 9002 11382 9142 11410
rect 9170 11382 9175 11410
rect 2233 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2375 11382
rect 17593 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17735 11382
rect 9025 11270 9030 11298
rect 9058 11270 11662 11298
rect 11690 11270 11942 11298
rect 11970 11270 11975 11298
rect 7625 11158 7630 11186
rect 7658 11158 7798 11186
rect 7826 11158 12278 11186
rect 12306 11158 12311 11186
rect 15946 11158 18830 11186
rect 18858 11158 18863 11186
rect 8073 11102 8078 11130
rect 8106 11102 8974 11130
rect 9002 11102 9198 11130
rect 9226 11102 9231 11130
rect 9865 11102 9870 11130
rect 9898 11102 10654 11130
rect 10682 11102 10687 11130
rect 11209 11102 11214 11130
rect 11242 11102 13286 11130
rect 13314 11102 13319 11130
rect 15946 11074 15974 11158
rect 20600 11130 21000 11144
rect 20001 11102 20006 11130
rect 20034 11102 21000 11130
rect 20600 11088 21000 11102
rect 5609 11046 5614 11074
rect 5642 11046 6902 11074
rect 6930 11046 7406 11074
rect 7434 11046 7574 11074
rect 7602 11046 7910 11074
rect 7938 11046 7943 11074
rect 11769 11046 11774 11074
rect 11802 11046 12446 11074
rect 12474 11046 12479 11074
rect 14905 11046 14910 11074
rect 14938 11046 15974 11074
rect 7835 10990 7854 11018
rect 7882 10990 7887 11018
rect 9913 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10055 10990
rect 9473 10934 9478 10962
rect 9506 10934 9646 10962
rect 9674 10934 9814 10962
rect 9842 10934 9847 10962
rect 10761 10934 10766 10962
rect 10794 10934 11102 10962
rect 11130 10934 11830 10962
rect 11858 10934 11863 10962
rect 9417 10822 9422 10850
rect 9450 10822 9926 10850
rect 9954 10822 10598 10850
rect 10626 10822 10631 10850
rect 20600 10794 21000 10808
rect 7009 10766 7014 10794
rect 7042 10766 7854 10794
rect 7882 10766 7887 10794
rect 11713 10766 11718 10794
rect 11746 10766 12166 10794
rect 12194 10766 12199 10794
rect 13169 10766 13174 10794
rect 13202 10766 13678 10794
rect 13706 10766 13711 10794
rect 20001 10766 20006 10794
rect 20034 10766 21000 10794
rect 20600 10752 21000 10766
rect 6393 10710 6398 10738
rect 6426 10710 7182 10738
rect 7210 10710 7215 10738
rect 7457 10710 7462 10738
rect 7490 10710 7742 10738
rect 7770 10710 9646 10738
rect 9674 10710 9679 10738
rect 14737 10710 14742 10738
rect 14770 10710 15134 10738
rect 15162 10710 15167 10738
rect 8241 10654 8246 10682
rect 8274 10654 10374 10682
rect 10402 10654 11326 10682
rect 11354 10654 11359 10682
rect 2233 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2375 10598
rect 17593 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17735 10598
rect 10873 10486 10878 10514
rect 10906 10486 11886 10514
rect 11914 10486 11919 10514
rect 14233 10486 14238 10514
rect 14266 10486 14574 10514
rect 14602 10486 14607 10514
rect 9137 10430 9142 10458
rect 9170 10430 9534 10458
rect 9562 10430 10654 10458
rect 10682 10430 10687 10458
rect 11265 10430 11270 10458
rect 11298 10430 13454 10458
rect 13482 10430 14882 10458
rect 10033 10374 10038 10402
rect 10066 10374 11662 10402
rect 11690 10374 11695 10402
rect 14854 10346 14882 10430
rect 15297 10374 15302 10402
rect 15330 10374 18830 10402
rect 18858 10374 18863 10402
rect 8353 10318 8358 10346
rect 8386 10318 11046 10346
rect 11074 10318 11438 10346
rect 11466 10318 11471 10346
rect 14849 10318 14854 10346
rect 14882 10318 14887 10346
rect 9641 10262 9646 10290
rect 9674 10262 10150 10290
rect 10178 10262 10878 10290
rect 10906 10262 10911 10290
rect 9913 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10055 10206
rect 11265 10094 11270 10122
rect 11298 10094 11998 10122
rect 12026 10094 12031 10122
rect 12609 10094 12614 10122
rect 12642 10094 12894 10122
rect 12922 10094 13174 10122
rect 13202 10094 13342 10122
rect 13370 10094 14518 10122
rect 14546 10094 14551 10122
rect 8185 10038 8190 10066
rect 8218 10038 8694 10066
rect 8722 10038 9534 10066
rect 9562 10038 11158 10066
rect 11186 10038 11191 10066
rect 12105 10038 12110 10066
rect 12138 10038 12558 10066
rect 12586 10038 12591 10066
rect 12665 10038 12670 10066
rect 12698 10038 15974 10066
rect 12670 10010 12698 10038
rect 7513 9982 7518 10010
rect 7546 9982 7551 10010
rect 12329 9982 12334 10010
rect 12362 9982 12698 10010
rect 15946 10010 15974 10038
rect 15946 9982 18830 10010
rect 18858 9982 18863 10010
rect 7518 9954 7546 9982
rect 7518 9926 9814 9954
rect 9842 9926 9847 9954
rect 14177 9926 14182 9954
rect 14210 9926 14798 9954
rect 14826 9926 15974 9954
rect 15946 9898 15974 9926
rect 15946 9870 18830 9898
rect 18858 9870 18863 9898
rect 2233 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2375 9814
rect 17593 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17735 9814
rect 20600 9786 21000 9800
rect 11209 9758 11214 9786
rect 11242 9758 14238 9786
rect 14266 9758 15190 9786
rect 15218 9758 15223 9786
rect 20001 9758 20006 9786
rect 20034 9758 21000 9786
rect 20600 9744 21000 9758
rect 8185 9590 8190 9618
rect 8218 9590 8470 9618
rect 8498 9590 8806 9618
rect 8834 9590 8839 9618
rect 8969 9590 8974 9618
rect 9002 9590 10206 9618
rect 10234 9590 10239 9618
rect 8974 9562 9002 9590
rect 7345 9534 7350 9562
rect 7378 9534 9002 9562
rect 11713 9534 11718 9562
rect 11746 9534 13230 9562
rect 13258 9534 13263 9562
rect 2081 9478 2086 9506
rect 2114 9478 9422 9506
rect 9450 9478 9455 9506
rect 9809 9478 9814 9506
rect 9842 9478 10822 9506
rect 10850 9478 10855 9506
rect 20600 9450 21000 9464
rect 7849 9422 7854 9450
rect 7882 9422 9478 9450
rect 9506 9422 9511 9450
rect 20001 9422 20006 9450
rect 20034 9422 21000 9450
rect 7910 9394 7938 9422
rect 9913 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10055 9422
rect 20600 9408 21000 9422
rect 7905 9366 7910 9394
rect 7938 9366 7943 9394
rect 7625 9310 7630 9338
rect 7658 9310 8022 9338
rect 8050 9310 8055 9338
rect 10257 9310 10262 9338
rect 10290 9310 10934 9338
rect 10962 9310 10967 9338
rect 10033 9254 10038 9282
rect 10066 9254 10598 9282
rect 10626 9254 10631 9282
rect 13281 9254 13286 9282
rect 13314 9254 14378 9282
rect 6561 9198 6566 9226
rect 6594 9198 7742 9226
rect 7770 9198 7775 9226
rect 8073 9198 8078 9226
rect 8106 9198 8806 9226
rect 8834 9198 8839 9226
rect 9025 9198 9030 9226
rect 9058 9198 9310 9226
rect 9338 9198 9702 9226
rect 9730 9198 9735 9226
rect 10649 9198 10654 9226
rect 10682 9198 13510 9226
rect 13538 9198 13543 9226
rect 8806 9170 8834 9198
rect 14350 9170 14378 9254
rect 15946 9198 18830 9226
rect 18858 9198 18863 9226
rect 15946 9170 15974 9198
rect 6225 9142 6230 9170
rect 6258 9142 7798 9170
rect 7826 9142 8134 9170
rect 8162 9142 8167 9170
rect 8806 9142 9366 9170
rect 9394 9142 9399 9170
rect 10593 9142 10598 9170
rect 10626 9142 12726 9170
rect 12754 9142 13454 9170
rect 14345 9142 14350 9170
rect 14378 9142 15974 9170
rect 9529 9086 9534 9114
rect 9562 9086 10262 9114
rect 10290 9086 11326 9114
rect 11354 9086 11359 9114
rect 9305 9030 9310 9058
rect 9338 9030 9646 9058
rect 9674 9030 9679 9058
rect 13426 9030 13454 9142
rect 20600 9114 21000 9128
rect 20001 9086 20006 9114
rect 20034 9086 21000 9114
rect 20600 9072 21000 9086
rect 13482 9030 13487 9058
rect 2233 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2375 9030
rect 17593 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17735 9030
rect 9249 8974 9254 9002
rect 9282 8974 9478 9002
rect 9506 8974 9511 9002
rect 7625 8862 7630 8890
rect 7658 8862 8078 8890
rect 8106 8862 8111 8890
rect 8577 8862 8582 8890
rect 8610 8862 8974 8890
rect 9002 8862 9198 8890
rect 9226 8862 10374 8890
rect 10402 8862 10654 8890
rect 10682 8862 10687 8890
rect 7737 8806 7742 8834
rect 7770 8806 8134 8834
rect 8162 8806 8167 8834
rect 9921 8806 9926 8834
rect 9954 8806 10262 8834
rect 10290 8806 10710 8834
rect 10738 8806 10743 8834
rect 7401 8750 7406 8778
rect 7434 8750 8862 8778
rect 8890 8750 8895 8778
rect 8129 8694 8134 8722
rect 8162 8694 9478 8722
rect 9506 8694 10094 8722
rect 10122 8694 10127 8722
rect 10817 8694 10822 8722
rect 10850 8694 11046 8722
rect 11074 8694 11662 8722
rect 11690 8694 11695 8722
rect 9913 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10055 8638
rect 10145 8358 10150 8386
rect 10178 8358 10430 8386
rect 10458 8358 10463 8386
rect 7681 8302 7686 8330
rect 7714 8302 8190 8330
rect 8218 8302 8974 8330
rect 9002 8302 9007 8330
rect 9697 8302 9702 8330
rect 9730 8302 10094 8330
rect 10122 8302 10127 8330
rect 2233 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2375 8246
rect 17593 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17735 8246
rect 7625 8078 7630 8106
rect 7658 8078 8078 8106
rect 8106 8078 8111 8106
rect 2137 8022 2142 8050
rect 2170 8022 6062 8050
rect 6090 8022 7686 8050
rect 7714 8022 7719 8050
rect 13113 8022 13118 8050
rect 13146 8022 13566 8050
rect 13594 8022 14014 8050
rect 14042 8022 14047 8050
rect 11545 7966 11550 7994
rect 11578 7966 11942 7994
rect 11970 7966 11975 7994
rect 13281 7966 13286 7994
rect 13314 7966 14686 7994
rect 14714 7966 14719 7994
rect 7121 7910 7126 7938
rect 7154 7910 8078 7938
rect 8106 7910 8111 7938
rect 10089 7910 10094 7938
rect 10122 7910 10654 7938
rect 10682 7910 10687 7938
rect 10817 7910 10822 7938
rect 10850 7910 11998 7938
rect 12026 7910 12031 7938
rect 13393 7910 13398 7938
rect 13426 7910 13958 7938
rect 13986 7910 13991 7938
rect 9913 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10055 7854
rect 0 7770 400 7784
rect 20600 7770 21000 7784
rect 0 7742 966 7770
rect 994 7742 999 7770
rect 10313 7742 10318 7770
rect 10346 7742 11438 7770
rect 11466 7742 13734 7770
rect 13762 7742 14630 7770
rect 14658 7742 14663 7770
rect 20001 7742 20006 7770
rect 20034 7742 21000 7770
rect 0 7728 400 7742
rect 20600 7728 21000 7742
rect 7681 7686 7686 7714
rect 7714 7686 7719 7714
rect 9865 7686 9870 7714
rect 9898 7686 10430 7714
rect 10458 7686 10463 7714
rect 14289 7686 14294 7714
rect 14322 7686 14798 7714
rect 14826 7686 15974 7714
rect 7686 7602 7714 7686
rect 15946 7658 15974 7686
rect 8241 7630 8246 7658
rect 8274 7630 8974 7658
rect 9002 7630 9366 7658
rect 9394 7630 9590 7658
rect 9618 7630 9623 7658
rect 10481 7630 10486 7658
rect 10514 7630 10934 7658
rect 10962 7630 11746 7658
rect 15946 7630 18830 7658
rect 18858 7630 18863 7658
rect 6729 7574 6734 7602
rect 6762 7574 7518 7602
rect 7546 7574 7551 7602
rect 7686 7574 8862 7602
rect 8890 7574 8895 7602
rect 9081 7574 9086 7602
rect 9114 7574 9814 7602
rect 9842 7574 10542 7602
rect 10570 7574 10575 7602
rect 7686 7490 7714 7574
rect 11718 7546 11746 7630
rect 13617 7574 13622 7602
rect 13650 7574 14462 7602
rect 14490 7574 18942 7602
rect 18970 7574 18975 7602
rect 11718 7518 12110 7546
rect 12138 7518 12670 7546
rect 12698 7518 12894 7546
rect 12922 7518 12927 7546
rect 7681 7462 7686 7490
rect 7714 7462 7719 7490
rect 2233 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2375 7462
rect 17593 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17735 7462
rect 20600 7434 21000 7448
rect 20001 7406 20006 7434
rect 20034 7406 21000 7434
rect 20600 7392 21000 7406
rect 7961 7294 7966 7322
rect 7994 7294 8806 7322
rect 8834 7294 8839 7322
rect 10705 7294 10710 7322
rect 10738 7294 11046 7322
rect 11074 7294 11079 7322
rect 10257 7238 10262 7266
rect 10290 7238 10990 7266
rect 11018 7238 11023 7266
rect 10369 7182 10374 7210
rect 10402 7182 11214 7210
rect 11242 7182 11662 7210
rect 11690 7182 11695 7210
rect 9137 7126 9142 7154
rect 9170 7126 9758 7154
rect 9786 7126 9791 7154
rect 20600 7098 21000 7112
rect 20113 7070 20118 7098
rect 20146 7070 21000 7098
rect 9913 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10055 7070
rect 20600 7056 21000 7070
rect 8801 6958 8806 6986
rect 8834 6958 9030 6986
rect 9058 6958 9063 6986
rect 11097 6790 11102 6818
rect 11130 6790 11886 6818
rect 11914 6790 11919 6818
rect 6953 6734 6958 6762
rect 6986 6734 8246 6762
rect 8274 6734 8279 6762
rect 2233 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2375 6678
rect 17593 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17735 6678
rect 7793 6510 7798 6538
rect 7826 6510 8190 6538
rect 8218 6510 8750 6538
rect 8778 6510 9534 6538
rect 9562 6510 10374 6538
rect 10402 6510 10407 6538
rect 9913 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10055 6286
rect 2233 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2375 5894
rect 17593 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17735 5894
rect 9913 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10055 5502
rect 2233 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2375 5110
rect 17593 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17735 5110
rect 9913 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10055 4718
rect 2233 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2375 4326
rect 17593 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17735 4326
rect 9913 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10055 3934
rect 2233 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2375 3542
rect 17593 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17735 3542
rect 9913 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10055 3150
rect 2233 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2375 2758
rect 17593 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17735 2758
rect 8073 2590 8078 2618
rect 8106 2590 8694 2618
rect 8722 2590 8727 2618
rect 9913 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10055 2366
rect 9753 2030 9758 2058
rect 9786 2030 10374 2058
rect 10402 2030 10407 2058
rect 2233 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2375 1974
rect 17593 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17735 1974
rect 11881 1806 11886 1834
rect 11914 1806 12782 1834
rect 12810 1806 12815 1834
rect 9913 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10055 1582
<< via3 >>
rect 2238 19194 2266 19222
rect 2290 19194 2318 19222
rect 2342 19194 2370 19222
rect 17598 19194 17626 19222
rect 17650 19194 17678 19222
rect 17702 19194 17730 19222
rect 9918 18802 9946 18830
rect 9970 18802 9998 18830
rect 10022 18802 10050 18830
rect 2238 18410 2266 18438
rect 2290 18410 2318 18438
rect 2342 18410 2370 18438
rect 17598 18410 17626 18438
rect 17650 18410 17678 18438
rect 17702 18410 17730 18438
rect 9918 18018 9946 18046
rect 9970 18018 9998 18046
rect 10022 18018 10050 18046
rect 2238 17626 2266 17654
rect 2290 17626 2318 17654
rect 2342 17626 2370 17654
rect 17598 17626 17626 17654
rect 17650 17626 17678 17654
rect 17702 17626 17730 17654
rect 9918 17234 9946 17262
rect 9970 17234 9998 17262
rect 10022 17234 10050 17262
rect 2238 16842 2266 16870
rect 2290 16842 2318 16870
rect 2342 16842 2370 16870
rect 17598 16842 17626 16870
rect 17650 16842 17678 16870
rect 17702 16842 17730 16870
rect 9918 16450 9946 16478
rect 9970 16450 9998 16478
rect 10022 16450 10050 16478
rect 2238 16058 2266 16086
rect 2290 16058 2318 16086
rect 2342 16058 2370 16086
rect 17598 16058 17626 16086
rect 17650 16058 17678 16086
rect 17702 16058 17730 16086
rect 9918 15666 9946 15694
rect 9970 15666 9998 15694
rect 10022 15666 10050 15694
rect 2238 15274 2266 15302
rect 2290 15274 2318 15302
rect 2342 15274 2370 15302
rect 17598 15274 17626 15302
rect 17650 15274 17678 15302
rect 17702 15274 17730 15302
rect 9918 14882 9946 14910
rect 9970 14882 9998 14910
rect 10022 14882 10050 14910
rect 2238 14490 2266 14518
rect 2290 14490 2318 14518
rect 2342 14490 2370 14518
rect 17598 14490 17626 14518
rect 17650 14490 17678 14518
rect 17702 14490 17730 14518
rect 9918 14098 9946 14126
rect 9970 14098 9998 14126
rect 10022 14098 10050 14126
rect 2238 13706 2266 13734
rect 2290 13706 2318 13734
rect 2342 13706 2370 13734
rect 17598 13706 17626 13734
rect 17650 13706 17678 13734
rect 17702 13706 17730 13734
rect 9918 13314 9946 13342
rect 9970 13314 9998 13342
rect 10022 13314 10050 13342
rect 2238 12922 2266 12950
rect 2290 12922 2318 12950
rect 2342 12922 2370 12950
rect 17598 12922 17626 12950
rect 17650 12922 17678 12950
rect 17702 12922 17730 12950
rect 9918 12530 9946 12558
rect 9970 12530 9998 12558
rect 10022 12530 10050 12558
rect 2238 12138 2266 12166
rect 2290 12138 2318 12166
rect 2342 12138 2370 12166
rect 17598 12138 17626 12166
rect 17650 12138 17678 12166
rect 17702 12138 17730 12166
rect 9918 11746 9946 11774
rect 9970 11746 9998 11774
rect 10022 11746 10050 11774
rect 2238 11354 2266 11382
rect 2290 11354 2318 11382
rect 2342 11354 2370 11382
rect 17598 11354 17626 11382
rect 17650 11354 17678 11382
rect 17702 11354 17730 11382
rect 7854 10990 7882 11018
rect 9918 10962 9946 10990
rect 9970 10962 9998 10990
rect 10022 10962 10050 10990
rect 2238 10570 2266 10598
rect 2290 10570 2318 10598
rect 2342 10570 2370 10598
rect 17598 10570 17626 10598
rect 17650 10570 17678 10598
rect 17702 10570 17730 10598
rect 9918 10178 9946 10206
rect 9970 10178 9998 10206
rect 10022 10178 10050 10206
rect 2238 9786 2266 9814
rect 2290 9786 2318 9814
rect 2342 9786 2370 9814
rect 17598 9786 17626 9814
rect 17650 9786 17678 9814
rect 17702 9786 17730 9814
rect 7854 9422 7882 9450
rect 9918 9394 9946 9422
rect 9970 9394 9998 9422
rect 10022 9394 10050 9422
rect 2238 9002 2266 9030
rect 2290 9002 2318 9030
rect 2342 9002 2370 9030
rect 17598 9002 17626 9030
rect 17650 9002 17678 9030
rect 17702 9002 17730 9030
rect 9918 8610 9946 8638
rect 9970 8610 9998 8638
rect 10022 8610 10050 8638
rect 2238 8218 2266 8246
rect 2290 8218 2318 8246
rect 2342 8218 2370 8246
rect 17598 8218 17626 8246
rect 17650 8218 17678 8246
rect 17702 8218 17730 8246
rect 9918 7826 9946 7854
rect 9970 7826 9998 7854
rect 10022 7826 10050 7854
rect 2238 7434 2266 7462
rect 2290 7434 2318 7462
rect 2342 7434 2370 7462
rect 17598 7434 17626 7462
rect 17650 7434 17678 7462
rect 17702 7434 17730 7462
rect 9918 7042 9946 7070
rect 9970 7042 9998 7070
rect 10022 7042 10050 7070
rect 2238 6650 2266 6678
rect 2290 6650 2318 6678
rect 2342 6650 2370 6678
rect 17598 6650 17626 6678
rect 17650 6650 17678 6678
rect 17702 6650 17730 6678
rect 9918 6258 9946 6286
rect 9970 6258 9998 6286
rect 10022 6258 10050 6286
rect 2238 5866 2266 5894
rect 2290 5866 2318 5894
rect 2342 5866 2370 5894
rect 17598 5866 17626 5894
rect 17650 5866 17678 5894
rect 17702 5866 17730 5894
rect 9918 5474 9946 5502
rect 9970 5474 9998 5502
rect 10022 5474 10050 5502
rect 2238 5082 2266 5110
rect 2290 5082 2318 5110
rect 2342 5082 2370 5110
rect 17598 5082 17626 5110
rect 17650 5082 17678 5110
rect 17702 5082 17730 5110
rect 9918 4690 9946 4718
rect 9970 4690 9998 4718
rect 10022 4690 10050 4718
rect 2238 4298 2266 4326
rect 2290 4298 2318 4326
rect 2342 4298 2370 4326
rect 17598 4298 17626 4326
rect 17650 4298 17678 4326
rect 17702 4298 17730 4326
rect 9918 3906 9946 3934
rect 9970 3906 9998 3934
rect 10022 3906 10050 3934
rect 2238 3514 2266 3542
rect 2290 3514 2318 3542
rect 2342 3514 2370 3542
rect 17598 3514 17626 3542
rect 17650 3514 17678 3542
rect 17702 3514 17730 3542
rect 9918 3122 9946 3150
rect 9970 3122 9998 3150
rect 10022 3122 10050 3150
rect 2238 2730 2266 2758
rect 2290 2730 2318 2758
rect 2342 2730 2370 2758
rect 17598 2730 17626 2758
rect 17650 2730 17678 2758
rect 17702 2730 17730 2758
rect 9918 2338 9946 2366
rect 9970 2338 9998 2366
rect 10022 2338 10050 2366
rect 2238 1946 2266 1974
rect 2290 1946 2318 1974
rect 2342 1946 2370 1974
rect 17598 1946 17626 1974
rect 17650 1946 17678 1974
rect 17702 1946 17730 1974
rect 9918 1554 9946 1582
rect 9970 1554 9998 1582
rect 10022 1554 10050 1582
<< metal4 >>
rect 2224 19222 2384 19238
rect 2224 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2384 19222
rect 2224 18438 2384 19194
rect 2224 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2384 18438
rect 2224 17654 2384 18410
rect 2224 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2384 17654
rect 2224 16870 2384 17626
rect 2224 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2384 16870
rect 2224 16086 2384 16842
rect 2224 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2384 16086
rect 2224 15302 2384 16058
rect 2224 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2384 15302
rect 2224 14518 2384 15274
rect 2224 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2384 14518
rect 2224 13734 2384 14490
rect 2224 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2384 13734
rect 2224 12950 2384 13706
rect 2224 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2384 12950
rect 2224 12166 2384 12922
rect 2224 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2384 12166
rect 2224 11382 2384 12138
rect 2224 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2384 11382
rect 2224 10598 2384 11354
rect 9904 18830 10064 19238
rect 9904 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10064 18830
rect 9904 18046 10064 18802
rect 9904 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10064 18046
rect 9904 17262 10064 18018
rect 9904 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10064 17262
rect 9904 16478 10064 17234
rect 9904 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10064 16478
rect 9904 15694 10064 16450
rect 9904 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10064 15694
rect 9904 14910 10064 15666
rect 9904 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10064 14910
rect 9904 14126 10064 14882
rect 9904 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10064 14126
rect 9904 13342 10064 14098
rect 9904 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10064 13342
rect 9904 12558 10064 13314
rect 9904 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10064 12558
rect 9904 11774 10064 12530
rect 9904 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10064 11774
rect 2224 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2384 10598
rect 2224 9814 2384 10570
rect 2224 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2384 9814
rect 2224 9030 2384 9786
rect 7854 11018 7882 11023
rect 7854 9450 7882 10990
rect 7854 9417 7882 9422
rect 9904 10990 10064 11746
rect 9904 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10064 10990
rect 9904 10206 10064 10962
rect 9904 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10064 10206
rect 9904 9422 10064 10178
rect 2224 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2384 9030
rect 2224 8246 2384 9002
rect 2224 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2384 8246
rect 2224 7462 2384 8218
rect 2224 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2384 7462
rect 2224 6678 2384 7434
rect 2224 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2384 6678
rect 2224 5894 2384 6650
rect 2224 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2384 5894
rect 2224 5110 2384 5866
rect 2224 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2384 5110
rect 2224 4326 2384 5082
rect 2224 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2384 4326
rect 2224 3542 2384 4298
rect 2224 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2384 3542
rect 2224 2758 2384 3514
rect 2224 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2384 2758
rect 2224 1974 2384 2730
rect 2224 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2384 1974
rect 2224 1538 2384 1946
rect 9904 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10064 9422
rect 9904 8638 10064 9394
rect 9904 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10064 8638
rect 9904 7854 10064 8610
rect 9904 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10064 7854
rect 9904 7070 10064 7826
rect 9904 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10064 7070
rect 9904 6286 10064 7042
rect 9904 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10064 6286
rect 9904 5502 10064 6258
rect 9904 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10064 5502
rect 9904 4718 10064 5474
rect 9904 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10064 4718
rect 9904 3934 10064 4690
rect 9904 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10064 3934
rect 9904 3150 10064 3906
rect 9904 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10064 3150
rect 9904 2366 10064 3122
rect 9904 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10064 2366
rect 9904 1582 10064 2338
rect 9904 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10064 1582
rect 9904 1538 10064 1554
rect 17584 19222 17744 19238
rect 17584 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17744 19222
rect 17584 18438 17744 19194
rect 17584 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17744 18438
rect 17584 17654 17744 18410
rect 17584 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17744 17654
rect 17584 16870 17744 17626
rect 17584 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17744 16870
rect 17584 16086 17744 16842
rect 17584 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17744 16086
rect 17584 15302 17744 16058
rect 17584 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17744 15302
rect 17584 14518 17744 15274
rect 17584 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17744 14518
rect 17584 13734 17744 14490
rect 17584 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17744 13734
rect 17584 12950 17744 13706
rect 17584 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17744 12950
rect 17584 12166 17744 12922
rect 17584 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17744 12166
rect 17584 11382 17744 12138
rect 17584 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17744 11382
rect 17584 10598 17744 11354
rect 17584 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17744 10598
rect 17584 9814 17744 10570
rect 17584 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17744 9814
rect 17584 9030 17744 9786
rect 17584 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17744 9030
rect 17584 8246 17744 9002
rect 17584 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17744 8246
rect 17584 7462 17744 8218
rect 17584 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17744 7462
rect 17584 6678 17744 7434
rect 17584 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17744 6678
rect 17584 5894 17744 6650
rect 17584 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17744 5894
rect 17584 5110 17744 5866
rect 17584 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17744 5110
rect 17584 4326 17744 5082
rect 17584 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17744 4326
rect 17584 3542 17744 4298
rect 17584 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17744 3542
rect 17584 2758 17744 3514
rect 17584 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17744 2758
rect 17584 1974 17744 2730
rect 17584 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17744 1974
rect 17584 1538 17744 1946
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _101_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7952 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _102_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8736 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _103_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9912 0 -1 13328
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _104_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12096 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _105_
timestamp 1698175906
transform 1 0 10640 0 -1 13328
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _106_
timestamp 1698175906
transform 1 0 7784 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _107_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8904 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _108_
timestamp 1698175906
transform 1 0 9240 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _109_
timestamp 1698175906
transform 1 0 11480 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _110_
timestamp 1698175906
transform 1 0 8344 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _111_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9128 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _112_
timestamp 1698175906
transform -1 0 9968 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _113_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11424 0 1 11760
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _114_
timestamp 1698175906
transform -1 0 12824 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _115_
timestamp 1698175906
transform -1 0 10864 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _116_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10584 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _117_
timestamp 1698175906
transform -1 0 10360 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _118_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10024 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _119_
timestamp 1698175906
transform 1 0 6888 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _120_
timestamp 1698175906
transform 1 0 7224 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _121_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 7784 0 -1 10976
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _122_
timestamp 1698175906
transform -1 0 6496 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _123_
timestamp 1698175906
transform -1 0 9128 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _124_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10528 0 -1 10976
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _125_
timestamp 1698175906
transform -1 0 8232 0 1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _126_
timestamp 1698175906
transform 1 0 9576 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _127_
timestamp 1698175906
transform 1 0 10024 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _128_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10360 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _129_
timestamp 1698175906
transform -1 0 8008 0 -1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _130_
timestamp 1698175906
transform 1 0 9464 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _131_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9240 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _132_
timestamp 1698175906
transform -1 0 9128 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__mux2_2  _133_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7112 0 1 8624
box -43 -43 883 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _134_
timestamp 1698175906
transform -1 0 7000 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _135_
timestamp 1698175906
transform 1 0 9912 0 -1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _136_
timestamp 1698175906
transform 1 0 10584 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _137_
timestamp 1698175906
transform 1 0 10584 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _138_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 12096 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _139_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11200 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _140_
timestamp 1698175906
transform -1 0 11480 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _141_
timestamp 1698175906
transform -1 0 14336 0 1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _142_
timestamp 1698175906
transform -1 0 11144 0 -1 9408
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _143_
timestamp 1698175906
transform -1 0 8960 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__xnor2_1  _144_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7728 0 -1 10192
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _145_
timestamp 1698175906
transform -1 0 11424 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _146_
timestamp 1698175906
transform -1 0 13608 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _147_
timestamp 1698175906
transform 1 0 13496 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _148_
timestamp 1698175906
transform -1 0 13384 0 1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _149_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11760 0 -1 11760
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _150_
timestamp 1698175906
transform -1 0 12992 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _151_
timestamp 1698175906
transform 1 0 9240 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _152_
timestamp 1698175906
transform 1 0 9688 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _153_
timestamp 1698175906
transform 1 0 10920 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _154_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10248 0 -1 7840
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _155_
timestamp 1698175906
transform -1 0 8400 0 -1 14112
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _156_
timestamp 1698175906
transform -1 0 7896 0 1 12544
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _157_
timestamp 1698175906
transform -1 0 9856 0 1 11760
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _158_
timestamp 1698175906
transform -1 0 9240 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _159_
timestamp 1698175906
transform 1 0 8680 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__or4_1  _160_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9968 0 -1 9408
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _161_
timestamp 1698175906
transform -1 0 12824 0 -1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _162_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8680 0 1 9408
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _163_
timestamp 1698175906
transform 1 0 10584 0 1 10192
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _164_
timestamp 1698175906
transform -1 0 11872 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _165_
timestamp 1698175906
transform 1 0 11872 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _166_
timestamp 1698175906
transform 1 0 13160 0 1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _167_
timestamp 1698175906
transform 1 0 13272 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _168_
timestamp 1698175906
transform -1 0 15400 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _169_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 14952 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _170_
timestamp 1698175906
transform -1 0 14336 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _171_
timestamp 1698175906
transform -1 0 13832 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _172_
timestamp 1698175906
transform 1 0 13832 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _173_
timestamp 1698175906
transform 1 0 14560 0 -1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _174_
timestamp 1698175906
transform -1 0 13384 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _175_
timestamp 1698175906
transform -1 0 8176 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _176_
timestamp 1698175906
transform -1 0 8288 0 -1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _177_
timestamp 1698175906
transform 1 0 7560 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _178_
timestamp 1698175906
transform -1 0 7448 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _179_
timestamp 1698175906
transform 1 0 6664 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _180_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10584 0 1 10976
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _181_
timestamp 1698175906
transform 1 0 12544 0 -1 14112
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _182_
timestamp 1698175906
transform 1 0 11592 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _183_
timestamp 1698175906
transform -1 0 11312 0 1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _184_
timestamp 1698175906
transform 1 0 10584 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _185_
timestamp 1698175906
transform 1 0 12264 0 1 10976
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _186_
timestamp 1698175906
transform -1 0 12432 0 -1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _187_
timestamp 1698175906
transform -1 0 9856 0 -1 7840
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _188_
timestamp 1698175906
transform 1 0 7560 0 1 7840
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _189_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7840 0 1 7840
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _190_
timestamp 1698175906
transform -1 0 9184 0 -1 7056
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _191_
timestamp 1698175906
transform 1 0 8792 0 -1 7840
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _192_
timestamp 1698175906
transform 1 0 9128 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai31_1  _193_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8904 0 -1 11760
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _194_
timestamp 1698175906
transform 1 0 10696 0 1 11760
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _195_
timestamp 1698175906
transform -1 0 11760 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _196_
timestamp 1698175906
transform -1 0 10472 0 1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _197_
timestamp 1698175906
transform -1 0 9856 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _198_
timestamp 1698175906
transform -1 0 9632 0 -1 10192
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _199_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9520 0 1 7056
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _200_
timestamp 1698175906
transform 1 0 7616 0 1 7056
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _201_
timestamp 1698175906
transform 1 0 8120 0 -1 7056
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _202_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11424 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _203_
timestamp 1698175906
transform 1 0 8848 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _204_
timestamp 1698175906
transform 1 0 5488 0 -1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _205_
timestamp 1698175906
transform 1 0 6104 0 -1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _206_
timestamp 1698175906
transform 1 0 6048 0 -1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _207_
timestamp 1698175906
transform 1 0 10808 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _208_
timestamp 1698175906
transform 1 0 13272 0 -1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _209_
timestamp 1698175906
transform 1 0 12544 0 -1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _210_
timestamp 1698175906
transform 1 0 10360 0 -1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _211_
timestamp 1698175906
transform 1 0 6776 0 -1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _212_
timestamp 1698175906
transform 1 0 7224 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _213_
timestamp 1698175906
transform 1 0 10808 0 1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _214_
timestamp 1698175906
transform 1 0 12824 0 -1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _215_
timestamp 1698175906
transform 1 0 13608 0 -1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _216_
timestamp 1698175906
transform 1 0 12936 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _217_
timestamp 1698175906
transform 1 0 12768 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _218_
timestamp 1698175906
transform -1 0 7560 0 -1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _219_
timestamp 1698175906
transform 1 0 10808 0 -1 14112
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _220_
timestamp 1698175906
transform 1 0 9184 0 -1 14112
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _221_
timestamp 1698175906
transform 1 0 12152 0 1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _222_
timestamp 1698175906
transform -1 0 7616 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _223_
timestamp 1698175906
transform -1 0 9520 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _224_
timestamp 1698175906
transform 1 0 7840 0 1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _225_
timestamp 1698175906
transform -1 0 11312 0 -1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _226_
timestamp 1698175906
transform 1 0 8624 0 1 6272
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _227_
timestamp 1698175906
transform 1 0 6496 0 -1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _230_
timestamp 1698175906
transform 1 0 14672 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _231_
timestamp 1698175906
transform 1 0 13776 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__202__CLK dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13160 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__203__CLK
timestamp 1698175906
transform -1 0 8848 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__204__CLK
timestamp 1698175906
transform 1 0 6888 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__205__CLK
timestamp 1698175906
transform 1 0 8120 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__206__CLK
timestamp 1698175906
transform 1 0 7784 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__207__CLK
timestamp 1698175906
transform 1 0 12656 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__208__CLK
timestamp 1698175906
transform 1 0 15008 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__209__CLK
timestamp 1698175906
transform 1 0 14280 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__210__CLK
timestamp 1698175906
transform 1 0 12096 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__211__CLK
timestamp 1698175906
transform 1 0 8400 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__212__CLK
timestamp 1698175906
transform 1 0 8848 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__213__CLK
timestamp 1698175906
transform 1 0 12544 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__214__CLK
timestamp 1698175906
transform 1 0 14560 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__215__CLK
timestamp 1698175906
transform 1 0 13160 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__216__CLK
timestamp 1698175906
transform 1 0 15008 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__217__CLK
timestamp 1698175906
transform 1 0 14616 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__218__CLK
timestamp 1698175906
transform 1 0 7560 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__219__CLK
timestamp 1698175906
transform -1 0 13048 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__220__CLK
timestamp 1698175906
transform -1 0 9184 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__221__CLK
timestamp 1698175906
transform 1 0 14224 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__222__CLK
timestamp 1698175906
transform 1 0 7728 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__223__CLK
timestamp 1698175906
transform 1 0 9520 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__224__CLK
timestamp 1698175906
transform 1 0 9968 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__225__CLK
timestamp 1698175906
transform 1 0 11312 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__226__CLK
timestamp 1698175906
transform 1 0 10360 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__227__CLK
timestamp 1698175906
transform -1 0 8232 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform -1 0 9464 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9632 0 -1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 10472 0 1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 11592 0 1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 2688 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 4592 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 6496 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8400 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_172
timestamp 1698175906
transform 1 0 10304 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_176
timestamp 1698175906
transform 1 0 10528 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_232
timestamp 1698175906
transform 1 0 13664 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_236
timestamp 1698175906
transform 1 0 13888 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 14112 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 16016 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 17920 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 19824 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 20048 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20160 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 4368 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 4704 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 8288 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 -1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_158
timestamp 1698175906
transform 1 0 9520 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_162
timestamp 1698175906
transform 1 0 9744 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_1_189
timestamp 1698175906
transform 1 0 11256 0 -1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_205
timestamp 1698175906
transform 1 0 12152 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698175906
transform 1 0 12376 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_212
timestamp 1698175906
transform 1 0 12544 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_276
timestamp 1698175906
transform 1 0 16128 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 16464 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 20048 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 20160 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 784 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 2576 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 2744 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 6328 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_107
timestamp 1698175906
transform 1 0 6664 0 1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_2_123 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7560 0 1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_131
timestamp 1698175906
transform 1 0 8008 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_159
timestamp 1698175906
transform 1 0 9576 0 1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698175906
transform 1 0 10584 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 14168 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 14504 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 18088 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 18424 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 784 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 4368 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 4704 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 8288 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 8624 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 12208 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 12544 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 16128 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 16464 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 20048 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 20160 0 -1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 784 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 2576 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 2744 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 6328 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 6664 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 10248 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 10584 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 14168 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 14504 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 18088 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 18424 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 784 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 4368 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 4704 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 8288 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 8624 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 12208 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 12544 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 16128 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 16464 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 20048 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 20160 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 784 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 2576 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 2744 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 6328 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 6664 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 10248 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 10584 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 14168 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 14504 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 18088 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 18424 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 784 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 4368 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 4704 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 8288 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 8624 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 12208 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 12544 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 16128 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 16464 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 20048 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 20160 0 -1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 784 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 2576 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 2744 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 6328 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 6664 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 10248 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 10584 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 14168 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 14504 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 18088 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 18424 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 784 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 4368 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 4704 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 8288 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 8624 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 12208 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 12544 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 16128 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 16464 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 20048 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 20160 0 -1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 784 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 2576 0 1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 2744 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 6328 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 6664 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 10248 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 10584 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 14168 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 14504 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 18088 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 18424 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 784 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 4368 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 4704 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 8288 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 8624 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 12208 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 12544 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 16128 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 16464 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 20048 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 20160 0 -1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 784 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 2576 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 2744 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 6328 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_107
timestamp 1698175906
transform 1 0 6664 0 1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_123
timestamp 1698175906
transform 1 0 7560 0 1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_131
timestamp 1698175906
transform 1 0 8008 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_135
timestamp 1698175906
transform 1 0 8232 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_139
timestamp 1698175906
transform 1 0 8456 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_141
timestamp 1698175906
transform 1 0 8568 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_171
timestamp 1698175906
transform 1 0 10248 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_177
timestamp 1698175906
transform 1 0 10584 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698175906
transform 1 0 14168 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 14504 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 18088 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 18424 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 784 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 4368 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_72
timestamp 1698175906
transform 1 0 4704 0 -1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_138
timestamp 1698175906
transform 1 0 8400 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_142
timestamp 1698175906
transform 1 0 8624 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_146
timestamp 1698175906
transform 1 0 8848 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_152
timestamp 1698175906
transform 1 0 9184 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_156
timestamp 1698175906
transform 1 0 9408 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_164
timestamp 1698175906
transform 1 0 9856 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_172
timestamp 1698175906
transform 1 0 10304 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_202
timestamp 1698175906
transform 1 0 11984 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_206
timestamp 1698175906
transform 1 0 12208 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_212
timestamp 1698175906
transform 1 0 12544 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_276
timestamp 1698175906
transform 1 0 16128 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 16464 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 20048 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 20160 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 784 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 2576 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 2744 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 6328 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_107
timestamp 1698175906
transform 1 0 6664 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_123
timestamp 1698175906
transform 1 0 7560 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_177
timestamp 1698175906
transform 1 0 10584 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_181
timestamp 1698175906
transform 1 0 10808 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_191
timestamp 1698175906
transform 1 0 11368 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_207
timestamp 1698175906
transform 1 0 12264 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_215
timestamp 1698175906
transform 1 0 12712 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_247
timestamp 1698175906
transform 1 0 14504 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_251
timestamp 1698175906
transform 1 0 14728 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_317
timestamp 1698175906
transform 1 0 18424 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_333
timestamp 1698175906
transform 1 0 19320 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_341
timestamp 1698175906
transform 1 0 19768 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 784 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 4368 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_72
timestamp 1698175906
transform 1 0 4704 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_88
timestamp 1698175906
transform 1 0 5600 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_92
timestamp 1698175906
transform 1 0 5824 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_94
timestamp 1698175906
transform 1 0 5936 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_124
timestamp 1698175906
transform 1 0 7616 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_128
timestamp 1698175906
transform 1 0 7840 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_136
timestamp 1698175906
transform 1 0 8288 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_142
timestamp 1698175906
transform 1 0 8624 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_144
timestamp 1698175906
transform 1 0 8736 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_164
timestamp 1698175906
transform 1 0 9856 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_212
timestamp 1698175906
transform 1 0 12544 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_216
timestamp 1698175906
transform 1 0 12768 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_218
timestamp 1698175906
transform 1 0 12880 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_254
timestamp 1698175906
transform 1 0 14896 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_258
timestamp 1698175906
transform 1 0 15120 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_274
timestamp 1698175906
transform 1 0 16016 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_278
timestamp 1698175906
transform 1 0 16240 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_282
timestamp 1698175906
transform 1 0 16464 0 -1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_314
timestamp 1698175906
transform 1 0 18256 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_322
timestamp 1698175906
transform 1 0 18704 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_28
timestamp 1698175906
transform 1 0 2240 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_32
timestamp 1698175906
transform 1 0 2464 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 2576 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 2744 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 6328 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_107
timestamp 1698175906
transform 1 0 6664 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_137
timestamp 1698175906
transform 1 0 8344 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_151
timestamp 1698175906
transform 1 0 9128 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_173
timestamp 1698175906
transform 1 0 10360 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_183
timestamp 1698175906
transform 1 0 10920 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_187
timestamp 1698175906
transform 1 0 11144 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_204
timestamp 1698175906
transform 1 0 12096 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_220
timestamp 1698175906
transform 1 0 12992 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_241
timestamp 1698175906
transform 1 0 14168 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 14504 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 18088 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_317
timestamp 1698175906
transform 1 0 18424 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_321
timestamp 1698175906
transform 1 0 18648 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698175906
transform 1 0 784 0 -1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698175906
transform 1 0 4368 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_72
timestamp 1698175906
transform 1 0 4704 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_88
timestamp 1698175906
transform 1 0 5600 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_125
timestamp 1698175906
transform 1 0 7672 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_129
timestamp 1698175906
transform 1 0 7896 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_137
timestamp 1698175906
transform 1 0 8344 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_139
timestamp 1698175906
transform 1 0 8456 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_142
timestamp 1698175906
transform 1 0 8624 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_146
timestamp 1698175906
transform 1 0 8848 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_163
timestamp 1698175906
transform 1 0 9800 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_195
timestamp 1698175906
transform 1 0 11592 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_203
timestamp 1698175906
transform 1 0 12040 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_207
timestamp 1698175906
transform 1 0 12264 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1698175906
transform 1 0 12376 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_212
timestamp 1698175906
transform 1 0 12544 0 -1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_276
timestamp 1698175906
transform 1 0 16128 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_282
timestamp 1698175906
transform 1 0 16464 0 -1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_346
timestamp 1698175906
transform 1 0 20048 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_348
timestamp 1698175906
transform 1 0 20160 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698175906
transform 1 0 784 0 1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 2576 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698175906
transform 1 0 2744 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698175906
transform 1 0 6328 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_113
timestamp 1698175906
transform 1 0 7000 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_135
timestamp 1698175906
transform 1 0 8232 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_143
timestamp 1698175906
transform 1 0 8680 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_157
timestamp 1698175906
transform 1 0 9464 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_173
timestamp 1698175906
transform 1 0 10360 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_183
timestamp 1698175906
transform 1 0 10920 0 1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_215
timestamp 1698175906
transform 1 0 12712 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_223
timestamp 1698175906
transform 1 0 13160 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_233
timestamp 1698175906
transform 1 0 13720 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_241
timestamp 1698175906
transform 1 0 14168 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698175906
transform 1 0 14504 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698175906
transform 1 0 18088 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_317
timestamp 1698175906
transform 1 0 18424 0 1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698175906
transform 1 0 784 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698175906
transform 1 0 4368 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_72
timestamp 1698175906
transform 1 0 4704 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_88
timestamp 1698175906
transform 1 0 5600 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_96
timestamp 1698175906
transform 1 0 6048 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_131
timestamp 1698175906
transform 1 0 8008 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_135
timestamp 1698175906
transform 1 0 8232 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_139
timestamp 1698175906
transform 1 0 8456 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_142
timestamp 1698175906
transform 1 0 8624 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_152
timestamp 1698175906
transform 1 0 9184 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_156
timestamp 1698175906
transform 1 0 9408 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_163
timestamp 1698175906
transform 1 0 9800 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_165
timestamp 1698175906
transform 1 0 9912 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_199
timestamp 1698175906
transform 1 0 11816 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_207
timestamp 1698175906
transform 1 0 12264 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_209
timestamp 1698175906
transform 1 0 12376 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_212
timestamp 1698175906
transform 1 0 12544 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_216
timestamp 1698175906
transform 1 0 12768 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_246
timestamp 1698175906
transform 1 0 14448 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_250
timestamp 1698175906
transform 1 0 14672 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_266
timestamp 1698175906
transform 1 0 15568 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_274
timestamp 1698175906
transform 1 0 16016 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_278
timestamp 1698175906
transform 1 0 16240 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_282
timestamp 1698175906
transform 1 0 16464 0 -1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_314
timestamp 1698175906
transform 1 0 18256 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_322
timestamp 1698175906
transform 1 0 18704 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 784 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 2576 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698175906
transform 1 0 2744 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698175906
transform 1 0 6328 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_107
timestamp 1698175906
transform 1 0 6664 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_123
timestamp 1698175906
transform 1 0 7560 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_127
timestamp 1698175906
transform 1 0 7784 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_129
timestamp 1698175906
transform 1 0 7896 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_136
timestamp 1698175906
transform 1 0 8288 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_153
timestamp 1698175906
transform 1 0 9240 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_173
timestamp 1698175906
transform 1 0 10360 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_210
timestamp 1698175906
transform 1 0 12432 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_214
timestamp 1698175906
transform 1 0 12656 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_222
timestamp 1698175906
transform 1 0 13104 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_228
timestamp 1698175906
transform 1 0 13440 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_237
timestamp 1698175906
transform 1 0 13944 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_244
timestamp 1698175906
transform 1 0 14336 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698175906
transform 1 0 14504 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698175906
transform 1 0 18088 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_317
timestamp 1698175906
transform 1 0 18424 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_321
timestamp 1698175906
transform 1 0 18648 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698175906
transform 1 0 784 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698175906
transform 1 0 4368 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_72
timestamp 1698175906
transform 1 0 4704 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_104
timestamp 1698175906
transform 1 0 6496 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_120
timestamp 1698175906
transform 1 0 7392 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_124
timestamp 1698175906
transform 1 0 7616 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_139
timestamp 1698175906
transform 1 0 8456 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_148
timestamp 1698175906
transform 1 0 8960 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_217
timestamp 1698175906
transform 1 0 12824 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_254
timestamp 1698175906
transform 1 0 14896 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_258
timestamp 1698175906
transform 1 0 15120 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_274
timestamp 1698175906
transform 1 0 16016 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_278
timestamp 1698175906
transform 1 0 16240 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_282
timestamp 1698175906
transform 1 0 16464 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_314
timestamp 1698175906
transform 1 0 18256 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_322
timestamp 1698175906
transform 1 0 18704 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 784 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 2576 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_37
timestamp 1698175906
transform 1 0 2744 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_69
timestamp 1698175906
transform 1 0 4536 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_85
timestamp 1698175906
transform 1 0 5432 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_93
timestamp 1698175906
transform 1 0 5880 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_97
timestamp 1698175906
transform 1 0 6104 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_104
timestamp 1698175906
transform 1 0 6496 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_107
timestamp 1698175906
transform 1 0 6664 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_192
timestamp 1698175906
transform 1 0 11424 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_194
timestamp 1698175906
transform 1 0 11536 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_263
timestamp 1698175906
transform 1 0 15400 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_295
timestamp 1698175906
transform 1 0 17192 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698175906
transform 1 0 18088 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_317
timestamp 1698175906
transform 1 0 18424 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698175906
transform 1 0 784 0 -1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698175906
transform 1 0 4368 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_72
timestamp 1698175906
transform 1 0 4704 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_80
timestamp 1698175906
transform 1 0 5152 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_84
timestamp 1698175906
transform 1 0 5376 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_133
timestamp 1698175906
transform 1 0 8120 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_137
timestamp 1698175906
transform 1 0 8344 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_139
timestamp 1698175906
transform 1 0 8456 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_142
timestamp 1698175906
transform 1 0 8624 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_150
timestamp 1698175906
transform 1 0 9072 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_152
timestamp 1698175906
transform 1 0 9184 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_182
timestamp 1698175906
transform 1 0 10864 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_190
timestamp 1698175906
transform 1 0 11312 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_208
timestamp 1698175906
transform 1 0 12320 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_212
timestamp 1698175906
transform 1 0 12544 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_220
timestamp 1698175906
transform 1 0 12992 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_222
timestamp 1698175906
transform 1 0 13104 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_260
timestamp 1698175906
transform 1 0 15232 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_276
timestamp 1698175906
transform 1 0 16128 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698175906
transform 1 0 16464 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_314
timestamp 1698175906
transform 1 0 18256 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_322
timestamp 1698175906
transform 1 0 18704 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698175906
transform 1 0 784 0 1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 2576 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698175906
transform 1 0 2744 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698175906
transform 1 0 6328 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_107
timestamp 1698175906
transform 1 0 6664 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_121
timestamp 1698175906
transform 1 0 7448 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_125
timestamp 1698175906
transform 1 0 7672 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_134
timestamp 1698175906
transform 1 0 8176 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_142
timestamp 1698175906
transform 1 0 8624 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_146
timestamp 1698175906
transform 1 0 8848 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_159
timestamp 1698175906
transform 1 0 9576 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_166
timestamp 1698175906
transform 1 0 9968 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_174
timestamp 1698175906
transform 1 0 10416 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_190
timestamp 1698175906
transform 1 0 11312 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_206
timestamp 1698175906
transform 1 0 12208 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_214
timestamp 1698175906
transform 1 0 12656 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_227
timestamp 1698175906
transform 1 0 13384 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_235
timestamp 1698175906
transform 1 0 13832 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_237
timestamp 1698175906
transform 1 0 13944 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_244
timestamp 1698175906
transform 1 0 14336 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_247
timestamp 1698175906
transform 1 0 14504 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_249
timestamp 1698175906
transform 1 0 14616 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_256
timestamp 1698175906
transform 1 0 15008 0 1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_288
timestamp 1698175906
transform 1 0 16800 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_304
timestamp 1698175906
transform 1 0 17696 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_312
timestamp 1698175906
transform 1 0 18144 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_314
timestamp 1698175906
transform 1 0 18256 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_317
timestamp 1698175906
transform 1 0 18424 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698175906
transform 1 0 18648 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2
timestamp 1698175906
transform 1 0 784 0 -1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_66
timestamp 1698175906
transform 1 0 4368 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_72
timestamp 1698175906
transform 1 0 4704 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_88
timestamp 1698175906
transform 1 0 5600 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_92
timestamp 1698175906
transform 1 0 5824 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_136
timestamp 1698175906
transform 1 0 8288 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_142
timestamp 1698175906
transform 1 0 8624 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_146
timestamp 1698175906
transform 1 0 8848 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_158
timestamp 1698175906
transform 1 0 9520 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_160
timestamp 1698175906
transform 1 0 9632 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_241
timestamp 1698175906
transform 1 0 14168 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_245
timestamp 1698175906
transform 1 0 14392 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_277
timestamp 1698175906
transform 1 0 16184 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_279
timestamp 1698175906
transform 1 0 16296 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_282
timestamp 1698175906
transform 1 0 16464 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_314
timestamp 1698175906
transform 1 0 18256 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_322
timestamp 1698175906
transform 1 0 18704 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_28
timestamp 1698175906
transform 1 0 2240 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_32
timestamp 1698175906
transform 1 0 2464 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 2576 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698175906
transform 1 0 2744 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698175906
transform 1 0 6328 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_113
timestamp 1698175906
transform 1 0 7000 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_121
timestamp 1698175906
transform 1 0 7448 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_125
timestamp 1698175906
transform 1 0 7672 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_127
timestamp 1698175906
transform 1 0 7784 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_164
timestamp 1698175906
transform 1 0 9856 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_168
timestamp 1698175906
transform 1 0 10080 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_172
timestamp 1698175906
transform 1 0 10304 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_174
timestamp 1698175906
transform 1 0 10416 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_177
timestamp 1698175906
transform 1 0 10584 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_188
timestamp 1698175906
transform 1 0 11200 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_201
timestamp 1698175906
transform 1 0 11928 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_240
timestamp 1698175906
transform 1 0 14112 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_244
timestamp 1698175906
transform 1 0 14336 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 14504 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 18088 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_317
timestamp 1698175906
transform 1 0 18424 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_321
timestamp 1698175906
transform 1 0 18648 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698175906
transform 1 0 784 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698175906
transform 1 0 4368 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_72
timestamp 1698175906
transform 1 0 4704 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_136
timestamp 1698175906
transform 1 0 8288 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_142
timestamp 1698175906
transform 1 0 8624 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_206
timestamp 1698175906
transform 1 0 12208 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_220
timestamp 1698175906
transform 1 0 12992 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_252
timestamp 1698175906
transform 1 0 14784 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_268
timestamp 1698175906
transform 1 0 15680 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_276
timestamp 1698175906
transform 1 0 16128 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_282
timestamp 1698175906
transform 1 0 16464 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_314
timestamp 1698175906
transform 1 0 18256 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_322
timestamp 1698175906
transform 1 0 18704 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698175906
transform 1 0 784 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 2576 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 2744 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 6328 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_107
timestamp 1698175906
transform 1 0 6664 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_123
timestamp 1698175906
transform 1 0 7560 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_129
timestamp 1698175906
transform 1 0 7896 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_137
timestamp 1698175906
transform 1 0 8344 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_140
timestamp 1698175906
transform 1 0 8512 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_142
timestamp 1698175906
transform 1 0 8624 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_151
timestamp 1698175906
transform 1 0 9128 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_167
timestamp 1698175906
transform 1 0 10024 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_177
timestamp 1698175906
transform 1 0 10584 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_241
timestamp 1698175906
transform 1 0 14168 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 14504 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 18088 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_317
timestamp 1698175906
transform 1 0 18424 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2
timestamp 1698175906
transform 1 0 784 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_66
timestamp 1698175906
transform 1 0 4368 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_72
timestamp 1698175906
transform 1 0 4704 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_104
timestamp 1698175906
transform 1 0 6496 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_108
timestamp 1698175906
transform 1 0 6720 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_138
timestamp 1698175906
transform 1 0 8400 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_142
timestamp 1698175906
transform 1 0 8624 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_153
timestamp 1698175906
transform 1 0 9240 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_157
timestamp 1698175906
transform 1 0 9464 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_165
timestamp 1698175906
transform 1 0 9912 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_173
timestamp 1698175906
transform 1 0 10360 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_177
timestamp 1698175906
transform 1 0 10584 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_184
timestamp 1698175906
transform 1 0 10976 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_192
timestamp 1698175906
transform 1 0 11424 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_194
timestamp 1698175906
transform 1 0 11536 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_203
timestamp 1698175906
transform 1 0 12040 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_209
timestamp 1698175906
transform 1 0 12376 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_217
timestamp 1698175906
transform 1 0 12824 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_249
timestamp 1698175906
transform 1 0 14616 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_265
timestamp 1698175906
transform 1 0 15512 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_273
timestamp 1698175906
transform 1 0 15960 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_277
timestamp 1698175906
transform 1 0 16184 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_279
timestamp 1698175906
transform 1 0 16296 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_282
timestamp 1698175906
transform 1 0 16464 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_346
timestamp 1698175906
transform 1 0 20048 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_348
timestamp 1698175906
transform 1 0 20160 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698175906
transform 1 0 784 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 2576 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 2744 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 6328 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_107
timestamp 1698175906
transform 1 0 6664 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_115
timestamp 1698175906
transform 1 0 7112 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_190
timestamp 1698175906
transform 1 0 11312 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_221
timestamp 1698175906
transform 1 0 13048 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_225
timestamp 1698175906
transform 1 0 13272 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_241
timestamp 1698175906
transform 1 0 14168 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 14504 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 18088 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_317
timestamp 1698175906
transform 1 0 18424 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 784 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 4368 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_72
timestamp 1698175906
transform 1 0 4704 0 -1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_104
timestamp 1698175906
transform 1 0 6496 0 -1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_120
timestamp 1698175906
transform 1 0 7392 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_128
timestamp 1698175906
transform 1 0 7840 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_132
timestamp 1698175906
transform 1 0 8064 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_138
timestamp 1698175906
transform 1 0 8400 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_142
timestamp 1698175906
transform 1 0 8624 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_146
timestamp 1698175906
transform 1 0 8848 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_217
timestamp 1698175906
transform 1 0 12824 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_221
timestamp 1698175906
transform 1 0 13048 0 -1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_253
timestamp 1698175906
transform 1 0 14840 0 -1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_269
timestamp 1698175906
transform 1 0 15736 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_277
timestamp 1698175906
transform 1 0 16184 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_279
timestamp 1698175906
transform 1 0 16296 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 16464 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 20048 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 20160 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 784 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 2576 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 2744 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 6328 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698175906
transform 1 0 6664 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698175906
transform 1 0 10248 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698175906
transform 1 0 10584 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698175906
transform 1 0 14168 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 14504 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 18088 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 18424 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 784 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 4368 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 4704 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 8288 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 8624 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 12208 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 12544 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 16128 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 16464 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 20048 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 20160 0 -1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 784 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 2576 0 1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 2744 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 6328 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 6664 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 10248 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 10584 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 14168 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 14504 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 18088 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 18424 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 784 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 4368 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 4704 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 8288 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 8624 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 12208 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 12544 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 16128 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 16464 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 20048 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 20160 0 -1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 784 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 2576 0 1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 2744 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 6328 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 6664 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 10248 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 10584 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 14168 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 14504 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 18088 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 18424 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 784 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 4368 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 4704 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 8288 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 8624 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 12208 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 12544 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 16128 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 16464 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 20048 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 20160 0 -1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 784 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 2576 0 1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 2744 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 6328 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 6664 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 10248 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 10584 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 14168 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 14504 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 18088 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 18424 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 784 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 4368 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 4704 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 8288 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 8624 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 12208 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 12544 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 16128 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 16464 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 20048 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 20160 0 -1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 784 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 2576 0 1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 2744 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 6328 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 6664 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 10248 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 10584 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 14168 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 14504 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 18088 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 18424 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 784 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 4368 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 4704 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 8288 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 8624 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 12208 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 12544 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 16128 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 16464 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 20048 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 20160 0 -1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 784 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 2576 0 1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 2744 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 6328 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_107
timestamp 1698175906
transform 1 0 6664 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_165
timestamp 1698175906
transform 1 0 9912 0 1 18032
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_173
timestamp 1698175906
transform 1 0 10360 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698175906
transform 1 0 10584 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 14168 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 14504 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 18088 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 18424 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 784 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 4368 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 4704 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 8288 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_142
timestamp 1698175906
transform 1 0 8624 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_150
timestamp 1698175906
transform 1 0 9072 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_154
timestamp 1698175906
transform 1 0 9296 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_207
timestamp 1698175906
transform 1 0 12264 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 12376 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_212
timestamp 1698175906
transform 1 0 12544 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_216
timestamp 1698175906
transform 1 0 12768 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_243
timestamp 1698175906
transform 1 0 14280 0 -1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_275
timestamp 1698175906
transform 1 0 16072 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_279
timestamp 1698175906
transform 1 0 16296 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 16464 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 20048 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 20160 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 784 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 2688 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 4592 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 6496 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_138
timestamp 1698175906
transform 1 0 8400 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_142
timestamp 1698175906
transform 1 0 8624 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_172
timestamp 1698175906
transform 1 0 10304 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_176
timestamp 1698175906
transform 1 0 10528 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_206
timestamp 1698175906
transform 1 0 12208 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_210
timestamp 1698175906
transform 1 0 12432 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_237
timestamp 1698175906
transform 1 0 13944 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_240
timestamp 1698175906
transform 1 0 14112 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_245
timestamp 1698175906
transform 1 0 14392 0 1 18816
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_261
timestamp 1698175906
transform 1 0 15288 0 1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_269
timestamp 1698175906
transform 1 0 15736 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_271
timestamp 1698175906
transform 1 0 15848 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 16016 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 17920 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 19824 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 20048 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 20160 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita7_25 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19992 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita7_26
timestamp 1698175906
transform -1 0 14392 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18760 0 1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform 1 0 9352 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform 1 0 10640 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform 1 0 9800 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform 1 0 8120 0 1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform 1 0 18760 0 -1 12544
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform 1 0 18760 0 -1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform 1 0 18760 0 1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform 1 0 18760 0 1 7840
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform 1 0 18760 0 -1 7840
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform -1 0 2240 0 1 7840
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform 1 0 8736 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform 1 0 18760 0 -1 9408
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform 1 0 12488 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform 1 0 10808 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform 1 0 18760 0 -1 10192
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform 1 0 8736 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform 1 0 8456 0 1 18032
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform -1 0 12096 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform 1 0 18760 0 -1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform 1 0 18760 0 1 9408
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform 1 0 12208 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform -1 0 2240 0 1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698175906
transform 1 0 12824 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 20328 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 20328 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 20328 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 20328 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 20328 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 20328 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 20328 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 672 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 20328 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 672 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 20328 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 672 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 20328 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 672 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 20328 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 672 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 20328 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 672 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 20328 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 672 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 20328 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 672 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 20328 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 672 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 20328 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 672 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 20328 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 672 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 20328 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 672 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 20328 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 672 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 20328 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 672 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 20328 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 672 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 20328 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 672 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 20328 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 672 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 20328 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 672 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 20328 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 672 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 20328 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 672 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 20328 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 672 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 20328 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 672 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 20328 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 672 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 20328 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 672 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 20328 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 672 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 20328 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 672 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 20328 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 672 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 20328 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 672 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 20328 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 672 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 20328 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 672 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 20328 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 672 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 20328 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 672 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 20328 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 672 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 20328 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 672 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 20328 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 672 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 20328 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 672 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 20328 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 672 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 20328 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 672 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 20328 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 2576 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 4480 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 6384 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 8288 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 10192 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 12096 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 14000 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 15904 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 17808 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 19712 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 4592 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 8512 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 12432 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 16352 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 6552 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 10472 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 14392 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 18312 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 4592 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 8512 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 12432 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 16352 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 6552 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 10472 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 14392 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 18312 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 4592 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 8512 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 12432 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 16352 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 6552 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 10472 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 14392 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 18312 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 4592 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 8512 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 12432 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 16352 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 2632 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 6552 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 10472 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 14392 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 18312 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 4592 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 8512 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 12432 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 16352 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 2632 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 6552 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 10472 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 14392 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 18312 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 4592 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 8512 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 12432 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 16352 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 2632 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 6552 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 10472 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 14392 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 18312 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 4592 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 8512 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 12432 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 16352 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 2632 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 6552 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 10472 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 14392 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 18312 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 4592 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 8512 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 12432 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 16352 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 2632 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 6552 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 10472 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 14392 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 18312 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 4592 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 8512 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 12432 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 16352 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 2632 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 6552 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 10472 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 14392 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 18312 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 4592 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 8512 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 12432 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 16352 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 2632 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 6552 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 10472 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 14392 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 18312 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 4592 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 8512 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 12432 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 16352 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 2632 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 6552 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 10472 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 14392 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 18312 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 4592 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 8512 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 12432 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 16352 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 2632 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 6552 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 10472 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 14392 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 18312 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 4592 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 8512 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 12432 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 16352 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 2632 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 6552 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 10472 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 14392 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 18312 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 4592 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 8512 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 12432 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 16352 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 2632 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 6552 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 10472 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 14392 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 18312 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 4592 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 8512 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 12432 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 16352 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 2632 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 6552 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 10472 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 14392 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 18312 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 4592 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 8512 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 12432 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 16352 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 2632 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 6552 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 10472 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 14392 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 18312 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 4592 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 8512 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 12432 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 16352 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 2632 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 6552 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 10472 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 14392 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 18312 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 4592 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 8512 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 12432 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 16352 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 2632 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 6552 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 10472 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 14392 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 18312 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 4592 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 8512 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 12432 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 16352 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 2632 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 6552 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 10472 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 14392 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 18312 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 4592 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 8512 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 12432 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 16352 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 2632 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 6552 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 10472 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 14392 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 18312 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 4592 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 8512 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 12432 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 16352 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 2632 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 6552 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 10472 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 14392 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 18312 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 4592 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 8512 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 12432 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 16352 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 2576 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 4480 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 6384 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 8288 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 10192 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 12096 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 14000 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 15904 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 17808 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 19712 0 1 18816
box -43 -43 155 435
<< labels >>
flabel metal3 s 0 13440 400 13496 0 FreeSans 224 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 20600 11088 21000 11144 0 FreeSans 224 0 0 0 segm[0]
port 1 nsew signal tristate
flabel metal2 s 9408 20600 9464 21000 0 FreeSans 224 90 0 0 segm[10]
port 2 nsew signal tristate
flabel metal2 s 11088 20600 11144 21000 0 FreeSans 224 90 0 0 segm[11]
port 3 nsew signal tristate
flabel metal2 s 9744 0 9800 400 0 FreeSans 224 90 0 0 segm[12]
port 4 nsew signal tristate
flabel metal2 s 8064 0 8120 400 0 FreeSans 224 90 0 0 segm[13]
port 5 nsew signal tristate
flabel metal3 s 20600 7056 21000 7112 0 FreeSans 224 0 0 0 segm[1]
port 6 nsew signal tristate
flabel metal3 s 20600 12096 21000 12152 0 FreeSans 224 0 0 0 segm[2]
port 7 nsew signal tristate
flabel metal3 s 20600 10752 21000 10808 0 FreeSans 224 0 0 0 segm[3]
port 8 nsew signal tristate
flabel metal2 s 14112 20600 14168 21000 0 FreeSans 224 90 0 0 segm[4]
port 9 nsew signal tristate
flabel metal3 s 20600 11760 21000 11816 0 FreeSans 224 0 0 0 segm[5]
port 10 nsew signal tristate
flabel metal3 s 20600 7728 21000 7784 0 FreeSans 224 0 0 0 segm[6]
port 11 nsew signal tristate
flabel metal3 s 20600 7392 21000 7448 0 FreeSans 224 0 0 0 segm[7]
port 12 nsew signal tristate
flabel metal3 s 0 7728 400 7784 0 FreeSans 224 0 0 0 segm[8]
port 13 nsew signal tristate
flabel metal2 s 9072 0 9128 400 0 FreeSans 224 90 0 0 segm[9]
port 14 nsew signal tristate
flabel metal3 s 20600 9072 21000 9128 0 FreeSans 224 0 0 0 sel[0]
port 15 nsew signal tristate
flabel metal2 s 12432 20600 12488 21000 0 FreeSans 224 90 0 0 sel[10]
port 16 nsew signal tristate
flabel metal2 s 10752 20600 10808 21000 0 FreeSans 224 90 0 0 sel[11]
port 17 nsew signal tristate
flabel metal3 s 20600 9744 21000 9800 0 FreeSans 224 0 0 0 sel[1]
port 18 nsew signal tristate
flabel metal2 s 9072 20600 9128 21000 0 FreeSans 224 90 0 0 sel[2]
port 19 nsew signal tristate
flabel metal2 s 8400 20600 8456 21000 0 FreeSans 224 90 0 0 sel[3]
port 20 nsew signal tristate
flabel metal2 s 11088 0 11144 400 0 FreeSans 224 90 0 0 sel[4]
port 21 nsew signal tristate
flabel metal3 s 20600 11424 21000 11480 0 FreeSans 224 0 0 0 sel[5]
port 22 nsew signal tristate
flabel metal3 s 20600 9408 21000 9464 0 FreeSans 224 0 0 0 sel[6]
port 23 nsew signal tristate
flabel metal2 s 11760 0 11816 400 0 FreeSans 224 90 0 0 sel[7]
port 24 nsew signal tristate
flabel metal3 s 0 11760 400 11816 0 FreeSans 224 0 0 0 sel[8]
port 25 nsew signal tristate
flabel metal2 s 12768 20600 12824 21000 0 FreeSans 224 90 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 2224 1538 2384 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 17584 1538 17744 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 9904 1538 10064 19238 0 FreeSans 640 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 10500 19208 10500 19208 0 vdd
rlabel metal1 10500 18816 10500 18816 0 vss
rlabel metal2 7084 11732 7084 11732 0 _000_
rlabel metal3 11508 13244 11508 13244 0 _001_
rlabel metal2 9660 13720 9660 13720 0 _002_
rlabel metal2 12180 11788 12180 11788 0 _003_
rlabel metal2 7140 7812 7140 7812 0 _004_
rlabel metal2 9044 7448 9044 7448 0 _005_
rlabel metal2 8316 11760 8316 11760 0 _006_
rlabel metal3 11228 11508 11228 11508 0 _007_
rlabel metal2 9128 6524 9128 6524 0 _008_
rlabel metal2 6972 6776 6972 6776 0 _009_
rlabel metal2 12572 13272 12572 13272 0 _010_
rlabel metal3 9436 13468 9436 13468 0 _011_
rlabel metal2 6244 10528 6244 10528 0 _012_
rlabel metal3 7168 9212 7168 9212 0 _013_
rlabel metal2 6524 8596 6524 8596 0 _014_
rlabel metal2 11312 7700 11312 7700 0 _015_
rlabel metal2 13636 9800 13636 9800 0 _016_
rlabel metal2 12936 11620 12936 11620 0 _017_
rlabel metal2 10780 7756 10780 7756 0 _018_
rlabel metal2 7644 12908 7644 12908 0 _019_
rlabel metal3 8260 12796 8260 12796 0 _020_
rlabel metal2 11284 9884 11284 9884 0 _021_
rlabel metal2 13356 8708 13356 8708 0 _022_
rlabel metal2 14084 10948 14084 10948 0 _023_
rlabel metal2 13412 7812 13412 7812 0 _024_
rlabel metal2 13244 7616 13244 7616 0 _025_
rlabel metal2 13132 11340 13132 11340 0 _026_
rlabel metal2 12124 12012 12124 12012 0 _027_
rlabel metal2 9968 7196 9968 7196 0 _028_
rlabel metal2 9100 7616 9100 7616 0 _029_
rlabel metal3 10892 7308 10892 7308 0 _030_
rlabel metal2 7980 13916 7980 13916 0 _031_
rlabel metal3 9128 12068 9128 12068 0 _032_
rlabel metal2 9100 12880 9100 12880 0 _033_
rlabel metal2 13468 8932 13468 8932 0 _034_
rlabel metal2 12572 10080 12572 10080 0 _035_
rlabel metal2 9520 11116 9520 11116 0 _036_
rlabel metal2 10892 10472 10892 10472 0 _037_
rlabel metal3 11956 10780 11956 10780 0 _038_
rlabel metal2 13384 8820 13384 8820 0 _039_
rlabel metal2 14896 10444 14896 10444 0 _040_
rlabel metal3 14420 10500 14420 10500 0 _041_
rlabel metal2 13804 8036 13804 8036 0 _042_
rlabel metal2 14700 7868 14700 7868 0 _043_
rlabel metal2 7812 11200 7812 11200 0 _044_
rlabel metal2 8036 11592 8036 11592 0 _045_
rlabel metal2 7252 11396 7252 11396 0 _046_
rlabel metal2 7084 11368 7084 11368 0 _047_
rlabel metal3 11592 11620 11592 11620 0 _048_
rlabel metal3 12348 13804 12348 13804 0 _049_
rlabel metal2 11004 13524 11004 13524 0 _050_
rlabel metal2 12376 11284 12376 11284 0 _051_
rlabel metal2 9716 7336 9716 7336 0 _052_
rlabel metal2 7868 7980 7868 7980 0 _053_
rlabel metal2 8932 7308 8932 7308 0 _054_
rlabel metal2 9240 11228 9240 11228 0 _055_
rlabel metal2 11340 11508 11340 11508 0 _056_
rlabel metal2 10080 7308 10080 7308 0 _057_
rlabel metal2 9688 6972 9688 6972 0 _058_
rlabel metal2 9800 7364 9800 7364 0 _059_
rlabel metal2 8204 7028 8204 7028 0 _060_
rlabel metal2 8820 9828 8820 9828 0 _061_
rlabel metal2 9128 11172 9128 11172 0 _062_
rlabel metal2 12180 13272 12180 13272 0 _063_
rlabel metal3 12516 13188 12516 13188 0 _064_
rlabel metal3 11340 13188 11340 13188 0 _065_
rlabel metal2 9324 10752 9324 10752 0 _066_
rlabel metal2 8988 11564 8988 11564 0 _067_
rlabel metal2 9548 8876 9548 8876 0 _068_
rlabel metal2 11732 9436 11732 9436 0 _069_
rlabel metal3 8904 8876 8904 8876 0 _070_
rlabel metal3 10276 11116 10276 11116 0 _071_
rlabel metal2 11564 12012 11564 12012 0 _072_
rlabel metal3 12320 13132 12320 13132 0 _073_
rlabel metal3 10276 10836 10276 10836 0 _074_
rlabel metal2 10724 9380 10724 9380 0 _075_
rlabel metal2 7476 10752 7476 10752 0 _076_
rlabel metal2 7252 10276 7252 10276 0 _077_
rlabel metal2 7532 10584 7532 10584 0 _078_
rlabel metal2 6412 10556 6412 10556 0 _079_
rlabel metal2 8988 6860 8988 6860 0 _080_
rlabel metal2 11340 9828 11340 9828 0 _081_
rlabel metal2 7924 8820 7924 8820 0 _082_
rlabel metal2 10108 8176 10108 8176 0 _083_
rlabel metal3 10640 7252 10640 7252 0 _084_
rlabel metal2 7812 12628 7812 12628 0 _085_
rlabel metal2 9716 9240 9716 9240 0 _086_
rlabel metal2 8204 8176 8204 8176 0 _087_
rlabel metal2 7364 11060 7364 11060 0 _088_
rlabel metal2 7084 8764 7084 8764 0 _089_
rlabel metal2 13748 7840 13748 7840 0 _090_
rlabel metal3 11424 7924 11424 7924 0 _091_
rlabel metal3 10808 7196 10808 7196 0 _092_
rlabel metal3 11760 7980 11760 7980 0 _093_
rlabel metal2 14252 9688 14252 9688 0 _094_
rlabel metal2 13748 9632 13748 9632 0 _095_
rlabel metal2 13524 9408 13524 9408 0 _096_
rlabel metal3 10360 10052 10360 10052 0 _097_
rlabel metal3 9716 10332 9716 10332 0 _098_
rlabel metal2 13468 10612 13468 10612 0 _099_
rlabel metal2 13580 9450 13580 9450 0 _100_
rlabel metal3 1239 13468 1239 13468 0 clk
rlabel metal2 11676 10220 11676 10220 0 clknet_0_clk
rlabel metal3 6272 11060 6272 11060 0 clknet_1_0__leaf_clk
rlabel metal2 11508 13720 11508 13720 0 clknet_1_1__leaf_clk
rlabel metal2 10500 13580 10500 13580 0 dut7.count\[0\]
rlabel metal2 7028 10752 7028 10752 0 dut7.count\[1\]
rlabel metal2 8036 9436 8036 9436 0 dut7.count\[2\]
rlabel metal3 8456 9212 8456 9212 0 dut7.count\[3\]
rlabel metal3 15442 11060 15442 11060 0 net1
rlabel metal2 14812 7672 14812 7672 0 net10
rlabel metal2 6076 7812 6076 7812 0 net11
rlabel metal3 8932 6972 8932 6972 0 net12
rlabel metal3 14364 9212 14364 9212 0 net13
rlabel metal2 12348 13944 12348 13944 0 net14
rlabel metal3 10920 13860 10920 13860 0 net15
rlabel metal3 15960 10024 15960 10024 0 net16
rlabel metal2 8820 18326 8820 18326 0 net17
rlabel metal2 8400 18228 8400 18228 0 net18
rlabel metal2 11788 2982 11788 2982 0 net19
rlabel metal2 9408 15960 9408 15960 0 net2
rlabel metal3 15022 11508 15022 11508 0 net20
rlabel metal2 14196 9744 14196 9744 0 net21
rlabel metal2 12292 4662 12292 4662 0 net22
rlabel metal2 6020 11732 6020 11732 0 net23
rlabel metal2 12964 16100 12964 16100 0 net24
rlabel metal2 20132 7112 20132 7112 0 net25
rlabel metal2 14196 18956 14196 18956 0 net26
rlabel metal2 9772 11592 9772 11592 0 net3
rlabel metal2 9856 2156 9856 2156 0 net4
rlabel metal2 8204 3374 8204 3374 0 net5
rlabel metal2 18956 12096 18956 12096 0 net6
rlabel metal2 15148 10696 15148 10696 0 net7
rlabel metal2 13916 11984 13916 11984 0 net8
rlabel metal2 13636 7756 13636 7756 0 net9
rlabel metal2 20020 11172 20020 11172 0 segm[0]
rlabel metal3 9688 18732 9688 18732 0 segm[10]
rlabel metal2 11116 19873 11116 19873 0 segm[11]
rlabel metal2 9772 1211 9772 1211 0 segm[12]
rlabel metal2 8092 1491 8092 1491 0 segm[13]
rlabel metal2 20020 12180 20020 12180 0 segm[2]
rlabel metal2 20020 10752 20020 10752 0 segm[3]
rlabel metal2 20020 11900 20020 11900 0 segm[5]
rlabel metal2 20020 7924 20020 7924 0 segm[6]
rlabel metal2 20020 7504 20020 7504 0 segm[7]
rlabel metal3 679 7756 679 7756 0 segm[8]
rlabel metal2 9100 1099 9100 1099 0 segm[9]
rlabel metal3 20321 9100 20321 9100 0 sel[0]
rlabel metal2 12460 19873 12460 19873 0 sel[10]
rlabel metal2 10780 19677 10780 19677 0 sel[11]
rlabel metal2 20020 9828 20020 9828 0 sel[1]
rlabel metal2 9100 19873 9100 19873 0 sel[2]
rlabel metal2 8428 19481 8428 19481 0 sel[3]
rlabel metal2 11116 1043 11116 1043 0 sel[4]
rlabel metal3 20321 11452 20321 11452 0 sel[5]
rlabel metal2 20020 9548 20020 9548 0 sel[6]
rlabel metal2 11788 427 11788 427 0 sel[7]
rlabel metal3 679 11788 679 11788 0 sel[8]
rlabel metal2 12796 19677 12796 19677 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 21000 21000
<< end >>
