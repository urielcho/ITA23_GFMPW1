magic
tech gf180mcuD
magscale 1 10
timestamp 1699642542
<< metal1 >>
rect 1344 38442 40656 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 40656 38442
rect 1344 38356 40656 38390
rect 18622 38274 18674 38286
rect 18622 38210 18674 38222
rect 22430 38274 22482 38286
rect 22430 38210 22482 38222
rect 25566 38274 25618 38286
rect 25566 38210 25618 38222
rect 27470 38274 27522 38286
rect 27470 38210 27522 38222
rect 17602 37998 17614 38050
rect 17666 37998 17678 38050
rect 21746 37998 21758 38050
rect 21810 37998 21822 38050
rect 24546 37998 24558 38050
rect 24610 37998 24622 38050
rect 5630 37938 5682 37950
rect 5630 37874 5682 37886
rect 34526 37938 34578 37950
rect 34526 37874 34578 37886
rect 1344 37658 40656 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 40656 37658
rect 1344 37572 40656 37606
rect 18398 37490 18450 37502
rect 18398 37426 18450 37438
rect 22094 37490 22146 37502
rect 22094 37426 22146 37438
rect 26238 37490 26290 37502
rect 26238 37426 26290 37438
rect 17378 37214 17390 37266
rect 17442 37214 17454 37266
rect 21074 37214 21086 37266
rect 21138 37214 21150 37266
rect 25218 37214 25230 37266
rect 25282 37214 25294 37266
rect 1344 36874 40656 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 40656 36874
rect 1344 36788 40656 36822
rect 17390 36706 17442 36718
rect 17390 36642 17442 36654
rect 16370 36430 16382 36482
rect 16434 36430 16446 36482
rect 1344 36090 40656 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 40656 36090
rect 1344 36004 40656 36038
rect 1344 35306 40656 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 40656 35306
rect 1344 35220 40656 35254
rect 1344 34522 40656 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 40656 34522
rect 1344 34436 40656 34470
rect 1344 33738 40656 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 40656 33738
rect 1344 33652 40656 33686
rect 1344 32954 40656 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 40656 32954
rect 1344 32868 40656 32902
rect 1344 32170 40656 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 40656 32170
rect 1344 32084 40656 32118
rect 1344 31386 40656 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 40656 31386
rect 1344 31300 40656 31334
rect 1710 31106 1762 31118
rect 1710 31042 1762 31054
rect 1344 30602 40656 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 40656 30602
rect 1344 30516 40656 30550
rect 1344 29818 40656 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 40656 29818
rect 1344 29732 40656 29766
rect 1344 29034 40656 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 40656 29034
rect 1344 28948 40656 28982
rect 1344 28250 40656 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 40656 28250
rect 1344 28164 40656 28198
rect 16270 28082 16322 28094
rect 16594 28030 16606 28082
rect 16658 28030 16670 28082
rect 16270 28018 16322 28030
rect 15934 27970 15986 27982
rect 15934 27906 15986 27918
rect 19730 27806 19742 27858
rect 19794 27806 19806 27858
rect 23214 27746 23266 27758
rect 20514 27694 20526 27746
rect 20578 27694 20590 27746
rect 22642 27694 22654 27746
rect 22706 27694 22718 27746
rect 23214 27682 23266 27694
rect 15822 27634 15874 27646
rect 15822 27570 15874 27582
rect 1344 27466 40656 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 40656 27466
rect 1344 27380 40656 27414
rect 21646 27186 21698 27198
rect 18498 27134 18510 27186
rect 18562 27134 18574 27186
rect 25218 27134 25230 27186
rect 25282 27134 25294 27186
rect 21646 27122 21698 27134
rect 15698 27022 15710 27074
rect 15762 27022 15774 27074
rect 22306 27022 22318 27074
rect 22370 27022 22382 27074
rect 21310 26962 21362 26974
rect 16370 26910 16382 26962
rect 16434 26910 16446 26962
rect 21310 26898 21362 26910
rect 21534 26962 21586 26974
rect 25678 26962 25730 26974
rect 23090 26910 23102 26962
rect 23154 26910 23166 26962
rect 21534 26898 21586 26910
rect 25678 26898 25730 26910
rect 18958 26850 19010 26862
rect 18958 26786 19010 26798
rect 21758 26850 21810 26862
rect 21758 26786 21810 26798
rect 21870 26850 21922 26862
rect 21870 26786 21922 26798
rect 40238 26850 40290 26862
rect 40238 26786 40290 26798
rect 1344 26682 40656 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 40656 26682
rect 1344 26596 40656 26630
rect 17614 26514 17666 26526
rect 17614 26450 17666 26462
rect 22766 26514 22818 26526
rect 22766 26450 22818 26462
rect 23550 26514 23602 26526
rect 23550 26450 23602 26462
rect 24110 26514 24162 26526
rect 24110 26450 24162 26462
rect 17838 26402 17890 26414
rect 17838 26338 17890 26350
rect 22990 26402 23042 26414
rect 22990 26338 23042 26350
rect 17390 26290 17442 26302
rect 23102 26290 23154 26302
rect 13794 26238 13806 26290
rect 13858 26238 13870 26290
rect 18610 26238 18622 26290
rect 18674 26238 18686 26290
rect 19618 26238 19630 26290
rect 19682 26238 19694 26290
rect 17390 26226 17442 26238
rect 23102 26226 23154 26238
rect 23886 26290 23938 26302
rect 23886 26226 23938 26238
rect 24222 26290 24274 26302
rect 24222 26226 24274 26238
rect 17502 26178 17554 26190
rect 14466 26126 14478 26178
rect 14530 26126 14542 26178
rect 16594 26126 16606 26178
rect 16658 26126 16670 26178
rect 18498 26126 18510 26178
rect 18562 26126 18574 26178
rect 20290 26126 20302 26178
rect 20354 26126 20366 26178
rect 22418 26126 22430 26178
rect 22482 26126 22494 26178
rect 17502 26114 17554 26126
rect 18286 26066 18338 26078
rect 18286 26002 18338 26014
rect 1344 25898 40656 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 40656 25898
rect 1344 25812 40656 25846
rect 22430 25730 22482 25742
rect 20626 25678 20638 25730
rect 20690 25727 20702 25730
rect 20850 25727 20862 25730
rect 20690 25681 20862 25727
rect 20690 25678 20702 25681
rect 20850 25678 20862 25681
rect 20914 25678 20926 25730
rect 22430 25666 22482 25678
rect 22542 25618 22594 25630
rect 27918 25618 27970 25630
rect 27458 25566 27470 25618
rect 27522 25566 27534 25618
rect 22542 25554 22594 25566
rect 27918 25554 27970 25566
rect 40014 25618 40066 25630
rect 40014 25554 40066 25566
rect 15598 25506 15650 25518
rect 15598 25442 15650 25454
rect 15822 25506 15874 25518
rect 15822 25442 15874 25454
rect 16270 25506 16322 25518
rect 16270 25442 16322 25454
rect 21198 25506 21250 25518
rect 21198 25442 21250 25454
rect 22094 25506 22146 25518
rect 24546 25454 24558 25506
rect 24610 25454 24622 25506
rect 37650 25454 37662 25506
rect 37714 25454 37726 25506
rect 22094 25442 22146 25454
rect 21534 25394 21586 25406
rect 21534 25330 21586 25342
rect 21758 25394 21810 25406
rect 25330 25342 25342 25394
rect 25394 25342 25406 25394
rect 21758 25330 21810 25342
rect 15934 25282 15986 25294
rect 15934 25218 15986 25230
rect 16830 25282 16882 25294
rect 16830 25218 16882 25230
rect 21422 25282 21474 25294
rect 21422 25218 21474 25230
rect 21982 25282 22034 25294
rect 21982 25218 22034 25230
rect 1344 25114 40656 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 40656 25114
rect 1344 25028 40656 25062
rect 21758 24946 21810 24958
rect 25566 24946 25618 24958
rect 23650 24894 23662 24946
rect 23714 24894 23726 24946
rect 21758 24882 21810 24894
rect 25566 24882 25618 24894
rect 21422 24834 21474 24846
rect 21422 24770 21474 24782
rect 21534 24834 21586 24846
rect 21534 24770 21586 24782
rect 25678 24834 25730 24846
rect 25678 24770 25730 24782
rect 26462 24834 26514 24846
rect 26462 24770 26514 24782
rect 25454 24722 25506 24734
rect 4274 24670 4286 24722
rect 4338 24670 4350 24722
rect 23874 24670 23886 24722
rect 23938 24670 23950 24722
rect 25218 24670 25230 24722
rect 25282 24670 25294 24722
rect 25454 24658 25506 24670
rect 25790 24722 25842 24734
rect 25790 24658 25842 24670
rect 1934 24498 1986 24510
rect 1934 24434 1986 24446
rect 26350 24498 26402 24510
rect 26350 24434 26402 24446
rect 1344 24330 40656 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 40656 24330
rect 1344 24244 40656 24278
rect 1934 24050 1986 24062
rect 13458 23998 13470 24050
rect 13522 23998 13534 24050
rect 17826 23998 17838 24050
rect 17890 23998 17902 24050
rect 1934 23986 1986 23998
rect 18398 23938 18450 23950
rect 4274 23886 4286 23938
rect 4338 23886 4350 23938
rect 14914 23886 14926 23938
rect 14978 23886 14990 23938
rect 18398 23874 18450 23886
rect 13806 23826 13858 23838
rect 15698 23774 15710 23826
rect 15762 23774 15774 23826
rect 13806 23762 13858 23774
rect 13582 23714 13634 23726
rect 13582 23650 13634 23662
rect 18062 23714 18114 23726
rect 18062 23650 18114 23662
rect 18286 23714 18338 23726
rect 18286 23650 18338 23662
rect 18846 23714 18898 23726
rect 18846 23650 18898 23662
rect 24222 23714 24274 23726
rect 24222 23650 24274 23662
rect 1344 23546 40656 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 40656 23546
rect 1344 23460 40656 23494
rect 15038 23378 15090 23390
rect 15038 23314 15090 23326
rect 16270 23378 16322 23390
rect 16270 23314 16322 23326
rect 16606 23378 16658 23390
rect 16606 23314 16658 23326
rect 24334 23266 24386 23278
rect 24334 23202 24386 23214
rect 24446 23266 24498 23278
rect 24446 23202 24498 23214
rect 15262 23154 15314 23166
rect 4274 23102 4286 23154
rect 4338 23102 4350 23154
rect 14690 23102 14702 23154
rect 14754 23102 14766 23154
rect 15262 23090 15314 23102
rect 15710 23154 15762 23166
rect 15710 23090 15762 23102
rect 16158 23154 16210 23166
rect 16158 23090 16210 23102
rect 16382 23154 16434 23166
rect 24670 23154 24722 23166
rect 17826 23102 17838 23154
rect 17890 23102 17902 23154
rect 21186 23102 21198 23154
rect 21250 23102 21262 23154
rect 37650 23102 37662 23154
rect 37714 23102 37726 23154
rect 16382 23090 16434 23102
rect 24670 23090 24722 23102
rect 15150 23042 15202 23054
rect 11778 22990 11790 23042
rect 11842 22990 11854 23042
rect 13906 22990 13918 23042
rect 13970 22990 13982 23042
rect 15150 22978 15202 22990
rect 17502 23042 17554 23054
rect 18610 22990 18622 23042
rect 18674 22990 18686 23042
rect 20738 22990 20750 23042
rect 20802 22990 20814 23042
rect 21858 22990 21870 23042
rect 21922 22990 21934 23042
rect 23986 22990 23998 23042
rect 24050 22990 24062 23042
rect 17502 22978 17554 22990
rect 1934 22930 1986 22942
rect 1934 22866 1986 22878
rect 40014 22930 40066 22942
rect 40014 22866 40066 22878
rect 1344 22762 40656 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 40656 22762
rect 1344 22676 40656 22710
rect 14030 22594 14082 22606
rect 14030 22530 14082 22542
rect 14366 22594 14418 22606
rect 14366 22530 14418 22542
rect 14702 22594 14754 22606
rect 14702 22530 14754 22542
rect 15150 22482 15202 22494
rect 13794 22430 13806 22482
rect 13858 22430 13870 22482
rect 15150 22418 15202 22430
rect 17838 22482 17890 22494
rect 17838 22418 17890 22430
rect 21646 22482 21698 22494
rect 40014 22482 40066 22494
rect 23202 22430 23214 22482
rect 23266 22430 23278 22482
rect 21646 22418 21698 22430
rect 40014 22418 40066 22430
rect 19742 22370 19794 22382
rect 20862 22370 20914 22382
rect 13682 22318 13694 22370
rect 13746 22318 13758 22370
rect 17602 22318 17614 22370
rect 17666 22318 17678 22370
rect 20290 22318 20302 22370
rect 20354 22318 20366 22370
rect 19742 22306 19794 22318
rect 20862 22306 20914 22318
rect 22990 22370 23042 22382
rect 26114 22318 26126 22370
rect 26178 22318 26190 22370
rect 37874 22318 37886 22370
rect 37938 22318 37950 22370
rect 22990 22306 23042 22318
rect 17950 22258 18002 22270
rect 18958 22258 19010 22270
rect 16930 22206 16942 22258
rect 16994 22206 17006 22258
rect 18274 22206 18286 22258
rect 18338 22206 18350 22258
rect 17950 22194 18002 22206
rect 18958 22194 19010 22206
rect 19854 22258 19906 22270
rect 19854 22194 19906 22206
rect 20078 22258 20130 22270
rect 20078 22194 20130 22206
rect 21310 22258 21362 22270
rect 21310 22194 21362 22206
rect 21534 22258 21586 22270
rect 28142 22258 28194 22270
rect 25330 22206 25342 22258
rect 25394 22206 25406 22258
rect 21534 22194 21586 22206
rect 28142 22194 28194 22206
rect 14478 22146 14530 22158
rect 14478 22082 14530 22094
rect 17278 22146 17330 22158
rect 17278 22082 17330 22094
rect 18622 22146 18674 22158
rect 20526 22146 20578 22158
rect 19282 22094 19294 22146
rect 19346 22094 19358 22146
rect 18622 22082 18674 22094
rect 20526 22082 20578 22094
rect 20750 22146 20802 22158
rect 20750 22082 20802 22094
rect 21758 22146 21810 22158
rect 21758 22082 21810 22094
rect 21870 22146 21922 22158
rect 21870 22082 21922 22094
rect 22318 22146 22370 22158
rect 22318 22082 22370 22094
rect 22430 22146 22482 22158
rect 22430 22082 22482 22094
rect 22542 22146 22594 22158
rect 22542 22082 22594 22094
rect 26574 22146 26626 22158
rect 26574 22082 26626 22094
rect 28030 22146 28082 22158
rect 28030 22082 28082 22094
rect 1344 21978 40656 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 40656 21978
rect 1344 21892 40656 21926
rect 14478 21810 14530 21822
rect 14478 21746 14530 21758
rect 17838 21810 17890 21822
rect 17838 21746 17890 21758
rect 17950 21810 18002 21822
rect 17950 21746 18002 21758
rect 18286 21810 18338 21822
rect 18286 21746 18338 21758
rect 25342 21810 25394 21822
rect 25342 21746 25394 21758
rect 25678 21810 25730 21822
rect 25678 21746 25730 21758
rect 14926 21698 14978 21710
rect 13234 21646 13246 21698
rect 13298 21646 13310 21698
rect 14926 21634 14978 21646
rect 15038 21586 15090 21598
rect 14018 21534 14030 21586
rect 14082 21534 14094 21586
rect 15038 21522 15090 21534
rect 17278 21586 17330 21598
rect 17278 21522 17330 21534
rect 17726 21586 17778 21598
rect 17726 21522 17778 21534
rect 18846 21586 18898 21598
rect 25230 21586 25282 21598
rect 19170 21534 19182 21586
rect 19234 21534 19246 21586
rect 18846 21522 18898 21534
rect 25230 21522 25282 21534
rect 25454 21586 25506 21598
rect 26226 21534 26238 21586
rect 26290 21534 26302 21586
rect 37650 21534 37662 21586
rect 37714 21534 37726 21586
rect 25454 21522 25506 21534
rect 18398 21474 18450 21486
rect 29486 21474 29538 21486
rect 11106 21422 11118 21474
rect 11170 21422 11182 21474
rect 23090 21422 23102 21474
rect 23154 21422 23166 21474
rect 26898 21422 26910 21474
rect 26962 21422 26974 21474
rect 29026 21422 29038 21474
rect 29090 21422 29102 21474
rect 18398 21410 18450 21422
rect 29486 21410 29538 21422
rect 29934 21474 29986 21486
rect 29934 21410 29986 21422
rect 40014 21474 40066 21486
rect 40014 21410 40066 21422
rect 14926 21362 14978 21374
rect 14926 21298 14978 21310
rect 29374 21362 29426 21374
rect 29374 21298 29426 21310
rect 1344 21194 40656 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 40656 21194
rect 1344 21108 40656 21142
rect 29710 20914 29762 20926
rect 17490 20862 17502 20914
rect 17554 20862 17566 20914
rect 21970 20862 21982 20914
rect 22034 20862 22046 20914
rect 29710 20850 29762 20862
rect 40014 20914 40066 20926
rect 40014 20850 40066 20862
rect 14478 20802 14530 20814
rect 21422 20802 21474 20814
rect 29262 20802 29314 20814
rect 20066 20750 20078 20802
rect 20130 20750 20142 20802
rect 22418 20750 22430 20802
rect 22482 20750 22494 20802
rect 23090 20750 23102 20802
rect 23154 20750 23166 20802
rect 14478 20738 14530 20750
rect 21422 20738 21474 20750
rect 29262 20738 29314 20750
rect 29934 20802 29986 20814
rect 29934 20738 29986 20750
rect 30158 20802 30210 20814
rect 30158 20738 30210 20750
rect 30606 20802 30658 20814
rect 37650 20750 37662 20802
rect 37714 20750 37726 20802
rect 30606 20738 30658 20750
rect 21982 20690 22034 20702
rect 26562 20638 26574 20690
rect 26626 20638 26638 20690
rect 21982 20626 22034 20638
rect 21534 20578 21586 20590
rect 14130 20526 14142 20578
rect 14194 20526 14206 20578
rect 21534 20514 21586 20526
rect 21758 20578 21810 20590
rect 21758 20514 21810 20526
rect 22206 20578 22258 20590
rect 22206 20514 22258 20526
rect 29374 20578 29426 20590
rect 29374 20514 29426 20526
rect 29486 20578 29538 20590
rect 29486 20514 29538 20526
rect 1344 20410 40656 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 40656 20410
rect 1344 20324 40656 20358
rect 18062 20242 18114 20254
rect 18062 20178 18114 20190
rect 26126 20242 26178 20254
rect 26126 20178 26178 20190
rect 15150 20130 15202 20142
rect 15150 20066 15202 20078
rect 15374 20130 15426 20142
rect 15374 20066 15426 20078
rect 16270 20130 16322 20142
rect 16270 20066 16322 20078
rect 16382 20130 16434 20142
rect 16382 20066 16434 20078
rect 17390 20130 17442 20142
rect 17390 20066 17442 20078
rect 18174 20130 18226 20142
rect 18174 20066 18226 20078
rect 19406 20130 19458 20142
rect 19406 20066 19458 20078
rect 20414 20130 20466 20142
rect 20414 20066 20466 20078
rect 20638 20130 20690 20142
rect 26014 20130 26066 20142
rect 23090 20078 23102 20130
rect 23154 20078 23166 20130
rect 24658 20078 24670 20130
rect 24722 20078 24734 20130
rect 20638 20066 20690 20078
rect 26014 20066 26066 20078
rect 26238 20130 26290 20142
rect 30046 20130 30098 20142
rect 27458 20078 27470 20130
rect 27522 20078 27534 20130
rect 26238 20066 26290 20078
rect 30046 20066 30098 20078
rect 15486 20018 15538 20030
rect 16942 20018 16994 20030
rect 20302 20018 20354 20030
rect 11218 19966 11230 20018
rect 11282 19966 11294 20018
rect 16594 19966 16606 20018
rect 16658 19966 16670 20018
rect 17602 19966 17614 20018
rect 17666 19966 17678 20018
rect 15486 19954 15538 19966
rect 16942 19954 16994 19966
rect 20302 19954 20354 19966
rect 22766 20018 22818 20030
rect 25566 20018 25618 20030
rect 24434 19966 24446 20018
rect 24498 19966 24510 20018
rect 26674 19966 26686 20018
rect 26738 19966 26750 20018
rect 22766 19954 22818 19966
rect 25566 19954 25618 19966
rect 14702 19906 14754 19918
rect 11890 19854 11902 19906
rect 11954 19854 11966 19906
rect 14018 19854 14030 19906
rect 14082 19854 14094 19906
rect 14702 19842 14754 19854
rect 14926 19906 14978 19918
rect 14926 19842 14978 19854
rect 19966 19906 20018 19918
rect 19966 19842 20018 19854
rect 25790 19906 25842 19918
rect 29586 19854 29598 19906
rect 29650 19854 29662 19906
rect 25790 19842 25842 19854
rect 19630 19794 19682 19806
rect 14354 19742 14366 19794
rect 14418 19742 14430 19794
rect 19630 19730 19682 19742
rect 25342 19794 25394 19806
rect 25342 19730 25394 19742
rect 1344 19626 40656 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 40656 19626
rect 1344 19540 40656 19574
rect 18062 19458 18114 19470
rect 18062 19394 18114 19406
rect 14254 19346 14306 19358
rect 14254 19282 14306 19294
rect 17502 19346 17554 19358
rect 25006 19346 25058 19358
rect 21410 19294 21422 19346
rect 21474 19294 21486 19346
rect 17502 19282 17554 19294
rect 25006 19282 25058 19294
rect 25902 19346 25954 19358
rect 25902 19282 25954 19294
rect 12686 19234 12738 19246
rect 12686 19170 12738 19182
rect 15934 19234 15986 19246
rect 15934 19170 15986 19182
rect 16382 19234 16434 19246
rect 16382 19170 16434 19182
rect 17278 19234 17330 19246
rect 23214 19234 23266 19246
rect 18050 19182 18062 19234
rect 18114 19182 18126 19234
rect 21858 19182 21870 19234
rect 21922 19182 21934 19234
rect 22194 19182 22206 19234
rect 22258 19182 22270 19234
rect 17278 19170 17330 19182
rect 23214 19170 23266 19182
rect 12350 19122 12402 19134
rect 12350 19058 12402 19070
rect 14926 19122 14978 19134
rect 14926 19058 14978 19070
rect 15262 19122 15314 19134
rect 15262 19058 15314 19070
rect 16606 19122 16658 19134
rect 16606 19058 16658 19070
rect 18398 19122 18450 19134
rect 22878 19122 22930 19134
rect 20402 19070 20414 19122
rect 20466 19070 20478 19122
rect 18398 19058 18450 19070
rect 22878 19058 22930 19070
rect 16158 19010 16210 19022
rect 20750 19010 20802 19022
rect 22990 19010 23042 19022
rect 16930 18958 16942 19010
rect 16994 18958 17006 19010
rect 21746 18958 21758 19010
rect 21810 18958 21822 19010
rect 16158 18946 16210 18958
rect 20750 18946 20802 18958
rect 22990 18946 23042 18958
rect 1344 18842 40656 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 40656 18842
rect 1344 18756 40656 18790
rect 15262 18674 15314 18686
rect 21534 18674 21586 18686
rect 22990 18674 23042 18686
rect 20066 18622 20078 18674
rect 20130 18622 20142 18674
rect 20850 18622 20862 18674
rect 20914 18622 20926 18674
rect 22642 18622 22654 18674
rect 22706 18622 22718 18674
rect 15262 18610 15314 18622
rect 21534 18610 21586 18622
rect 22990 18610 23042 18622
rect 23438 18674 23490 18686
rect 23438 18610 23490 18622
rect 26910 18674 26962 18686
rect 26910 18610 26962 18622
rect 15598 18562 15650 18574
rect 14914 18510 14926 18562
rect 14978 18510 14990 18562
rect 15598 18498 15650 18510
rect 15710 18562 15762 18574
rect 23550 18562 23602 18574
rect 21970 18510 21982 18562
rect 22034 18510 22046 18562
rect 15710 18498 15762 18510
rect 23550 18498 23602 18510
rect 15934 18450 15986 18462
rect 18174 18450 18226 18462
rect 16146 18398 16158 18450
rect 16210 18398 16222 18450
rect 15934 18386 15986 18398
rect 18174 18386 18226 18398
rect 18286 18450 18338 18462
rect 20526 18450 20578 18462
rect 18498 18398 18510 18450
rect 18562 18398 18574 18450
rect 19394 18398 19406 18450
rect 19458 18398 19470 18450
rect 19730 18398 19742 18450
rect 19794 18398 19806 18450
rect 18286 18386 18338 18398
rect 20526 18386 20578 18398
rect 21198 18450 21250 18462
rect 21198 18386 21250 18398
rect 22318 18450 22370 18462
rect 22318 18386 22370 18398
rect 23886 18450 23938 18462
rect 23886 18386 23938 18398
rect 25230 18450 25282 18462
rect 25230 18386 25282 18398
rect 25454 18450 25506 18462
rect 25454 18386 25506 18398
rect 25790 18450 25842 18462
rect 25790 18386 25842 18398
rect 26238 18450 26290 18462
rect 26238 18386 26290 18398
rect 27134 18450 27186 18462
rect 37650 18398 37662 18450
rect 37714 18398 37726 18450
rect 27134 18386 27186 18398
rect 25342 18338 25394 18350
rect 19058 18286 19070 18338
rect 19122 18286 19134 18338
rect 25342 18274 25394 18286
rect 26686 18338 26738 18350
rect 27010 18286 27022 18338
rect 27074 18286 27086 18338
rect 26686 18274 26738 18286
rect 23438 18226 23490 18238
rect 16146 18174 16158 18226
rect 16210 18174 16222 18226
rect 17714 18174 17726 18226
rect 17778 18174 17790 18226
rect 23438 18162 23490 18174
rect 23998 18226 24050 18238
rect 23998 18162 24050 18174
rect 26462 18226 26514 18238
rect 26462 18162 26514 18174
rect 40014 18226 40066 18238
rect 40014 18162 40066 18174
rect 1344 18058 40656 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 40656 18058
rect 1344 17972 40656 18006
rect 16270 17890 16322 17902
rect 16270 17826 16322 17838
rect 22654 17890 22706 17902
rect 22654 17826 22706 17838
rect 24222 17890 24274 17902
rect 28366 17890 28418 17902
rect 27682 17838 27694 17890
rect 27746 17887 27758 17890
rect 28130 17887 28142 17890
rect 27746 17841 28142 17887
rect 27746 17838 27758 17841
rect 28130 17838 28142 17841
rect 28194 17838 28206 17890
rect 24222 17826 24274 17838
rect 28366 17826 28418 17838
rect 1934 17778 1986 17790
rect 27918 17778 27970 17790
rect 22978 17726 22990 17778
rect 23042 17726 23054 17778
rect 27458 17726 27470 17778
rect 27522 17726 27534 17778
rect 1934 17714 1986 17726
rect 27918 17714 27970 17726
rect 40014 17778 40066 17790
rect 40014 17714 40066 17726
rect 14366 17666 14418 17678
rect 4274 17614 4286 17666
rect 4338 17614 4350 17666
rect 13682 17614 13694 17666
rect 13746 17614 13758 17666
rect 14366 17602 14418 17614
rect 14702 17666 14754 17678
rect 14702 17602 14754 17614
rect 18622 17666 18674 17678
rect 18622 17602 18674 17614
rect 21982 17666 22034 17678
rect 21982 17602 22034 17614
rect 23550 17666 23602 17678
rect 28478 17666 28530 17678
rect 23874 17614 23886 17666
rect 23938 17614 23950 17666
rect 24658 17614 24670 17666
rect 24722 17614 24734 17666
rect 37650 17614 37662 17666
rect 37714 17614 37726 17666
rect 23550 17602 23602 17614
rect 28478 17602 28530 17614
rect 14590 17554 14642 17566
rect 14590 17490 14642 17502
rect 16046 17554 16098 17566
rect 16046 17490 16098 17502
rect 17390 17554 17442 17566
rect 17390 17490 17442 17502
rect 17726 17554 17778 17566
rect 17726 17490 17778 17502
rect 18062 17554 18114 17566
rect 18062 17490 18114 17502
rect 18286 17554 18338 17566
rect 18286 17490 18338 17502
rect 18846 17554 18898 17566
rect 18846 17490 18898 17502
rect 18958 17554 19010 17566
rect 22878 17554 22930 17566
rect 19730 17502 19742 17554
rect 19794 17502 19806 17554
rect 18958 17490 19010 17502
rect 22878 17490 22930 17502
rect 23662 17554 23714 17566
rect 25330 17502 25342 17554
rect 25394 17502 25406 17554
rect 23662 17490 23714 17502
rect 13918 17442 13970 17454
rect 13918 17378 13970 17390
rect 14142 17442 14194 17454
rect 14142 17378 14194 17390
rect 14254 17442 14306 17454
rect 14254 17378 14306 17390
rect 15150 17442 15202 17454
rect 15150 17378 15202 17390
rect 16158 17442 16210 17454
rect 16158 17378 16210 17390
rect 16606 17442 16658 17454
rect 18174 17442 18226 17454
rect 16930 17390 16942 17442
rect 16994 17390 17006 17442
rect 16606 17378 16658 17390
rect 18174 17378 18226 17390
rect 19406 17442 19458 17454
rect 19406 17378 19458 17390
rect 21758 17442 21810 17454
rect 21758 17378 21810 17390
rect 21870 17442 21922 17454
rect 21870 17378 21922 17390
rect 23774 17442 23826 17454
rect 23774 17378 23826 17390
rect 1344 17274 40656 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 40656 17274
rect 1344 17188 40656 17222
rect 17838 17106 17890 17118
rect 20414 17106 20466 17118
rect 19730 17054 19742 17106
rect 19794 17054 19806 17106
rect 17838 17042 17890 17054
rect 20414 17042 20466 17054
rect 23326 17106 23378 17118
rect 23326 17042 23378 17054
rect 29822 17106 29874 17118
rect 29822 17042 29874 17054
rect 21758 16994 21810 17006
rect 13010 16942 13022 16994
rect 13074 16942 13086 16994
rect 27234 16942 27246 16994
rect 27298 16942 27310 16994
rect 21758 16930 21810 16942
rect 17614 16882 17666 16894
rect 12226 16830 12238 16882
rect 12290 16830 12302 16882
rect 17378 16830 17390 16882
rect 17442 16830 17454 16882
rect 17614 16818 17666 16830
rect 17950 16882 18002 16894
rect 21982 16882 22034 16894
rect 19170 16830 19182 16882
rect 19234 16830 19246 16882
rect 19394 16830 19406 16882
rect 19458 16830 19470 16882
rect 17950 16818 18002 16830
rect 21982 16818 22034 16830
rect 22318 16882 22370 16894
rect 22318 16818 22370 16830
rect 22654 16882 22706 16894
rect 22654 16818 22706 16830
rect 22878 16882 22930 16894
rect 22878 16818 22930 16830
rect 23550 16882 23602 16894
rect 26450 16830 26462 16882
rect 26514 16830 26526 16882
rect 23550 16818 23602 16830
rect 15598 16770 15650 16782
rect 20190 16770 20242 16782
rect 15138 16718 15150 16770
rect 15202 16718 15214 16770
rect 17490 16718 17502 16770
rect 17554 16718 17566 16770
rect 18834 16718 18846 16770
rect 18898 16718 18910 16770
rect 15598 16706 15650 16718
rect 20190 16706 20242 16718
rect 21870 16770 21922 16782
rect 21870 16706 21922 16718
rect 23102 16770 23154 16782
rect 23426 16718 23438 16770
rect 23490 16718 23502 16770
rect 29362 16718 29374 16770
rect 29426 16718 29438 16770
rect 23102 16706 23154 16718
rect 20526 16658 20578 16670
rect 20526 16594 20578 16606
rect 1344 16490 40656 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 40656 16490
rect 1344 16404 40656 16438
rect 21310 16322 21362 16334
rect 21310 16258 21362 16270
rect 21646 16322 21698 16334
rect 21646 16258 21698 16270
rect 22990 16322 23042 16334
rect 22990 16258 23042 16270
rect 23326 16322 23378 16334
rect 23326 16258 23378 16270
rect 22766 16210 22818 16222
rect 13458 16158 13470 16210
rect 13522 16158 13534 16210
rect 15586 16158 15598 16210
rect 15650 16158 15662 16210
rect 22766 16146 22818 16158
rect 23214 16210 23266 16222
rect 23214 16146 23266 16158
rect 16942 16098 16994 16110
rect 16258 16046 16270 16098
rect 16322 16046 16334 16098
rect 16942 16034 16994 16046
rect 17278 16098 17330 16110
rect 19282 16046 19294 16098
rect 19346 16046 19358 16098
rect 21298 16046 21310 16098
rect 21362 16046 21374 16098
rect 17278 16034 17330 16046
rect 19070 15986 19122 15998
rect 19070 15922 19122 15934
rect 17054 15874 17106 15886
rect 17054 15810 17106 15822
rect 17614 15874 17666 15886
rect 17614 15810 17666 15822
rect 22878 15874 22930 15886
rect 22878 15810 22930 15822
rect 1344 15706 40656 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 40656 15706
rect 1344 15620 40656 15654
rect 25230 15538 25282 15550
rect 25230 15474 25282 15486
rect 19854 15426 19906 15438
rect 14690 15374 14702 15426
rect 14754 15374 14766 15426
rect 19854 15362 19906 15374
rect 19966 15426 20018 15438
rect 19966 15362 20018 15374
rect 20862 15426 20914 15438
rect 20862 15362 20914 15374
rect 21198 15426 21250 15438
rect 22766 15426 22818 15438
rect 21522 15374 21534 15426
rect 21586 15374 21598 15426
rect 21198 15362 21250 15374
rect 22766 15362 22818 15374
rect 14018 15262 14030 15314
rect 14082 15262 14094 15314
rect 22978 15262 22990 15314
rect 23042 15262 23054 15314
rect 17502 15202 17554 15214
rect 16818 15150 16830 15202
rect 16882 15150 16894 15202
rect 17502 15138 17554 15150
rect 20638 15202 20690 15214
rect 20638 15138 20690 15150
rect 25342 15202 25394 15214
rect 25342 15138 25394 15150
rect 20302 15090 20354 15102
rect 20302 15026 20354 15038
rect 1344 14922 40656 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 40656 14922
rect 1344 14836 40656 14870
rect 19518 14642 19570 14654
rect 26126 14642 26178 14654
rect 16930 14590 16942 14642
rect 16994 14590 17006 14642
rect 19058 14590 19070 14642
rect 19122 14590 19134 14642
rect 23538 14590 23550 14642
rect 23602 14590 23614 14642
rect 25666 14590 25678 14642
rect 25730 14590 25742 14642
rect 19518 14578 19570 14590
rect 26126 14578 26178 14590
rect 16258 14478 16270 14530
rect 16322 14478 16334 14530
rect 20178 14478 20190 14530
rect 20242 14478 20254 14530
rect 22866 14478 22878 14530
rect 22930 14478 22942 14530
rect 20414 14306 20466 14318
rect 20414 14242 20466 14254
rect 1344 14138 40656 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 40656 14138
rect 1344 14052 40656 14086
rect 25342 13970 25394 13982
rect 25342 13906 25394 13918
rect 20626 13806 20638 13858
rect 20690 13806 20702 13858
rect 22530 13806 22542 13858
rect 22594 13806 22606 13858
rect 21410 13694 21422 13746
rect 21474 13694 21486 13746
rect 21858 13694 21870 13746
rect 21922 13694 21934 13746
rect 18498 13582 18510 13634
rect 18562 13582 18574 13634
rect 24658 13582 24670 13634
rect 24722 13582 24734 13634
rect 1344 13354 40656 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 40656 13354
rect 1344 13268 40656 13302
rect 21758 13074 21810 13086
rect 21758 13010 21810 13022
rect 1344 12570 40656 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 40656 12570
rect 1344 12484 40656 12518
rect 1344 11786 40656 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 40656 11786
rect 1344 11700 40656 11734
rect 1344 11002 40656 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 40656 11002
rect 1344 10916 40656 10950
rect 1344 10218 40656 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 40656 10218
rect 1344 10132 40656 10166
rect 1344 9434 40656 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 40656 9434
rect 1344 9348 40656 9382
rect 1344 8650 40656 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 40656 8650
rect 1344 8564 40656 8598
rect 1344 7866 40656 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 40656 7866
rect 1344 7780 40656 7814
rect 1344 7082 40656 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 40656 7082
rect 1344 6996 40656 7030
rect 1344 6298 40656 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 40656 6298
rect 1344 6212 40656 6246
rect 1344 5514 40656 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 40656 5514
rect 1344 5428 40656 5462
rect 1344 4730 40656 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 40656 4730
rect 1344 4644 40656 4678
rect 25218 4286 25230 4338
rect 25282 4286 25294 4338
rect 26238 4114 26290 4126
rect 26238 4050 26290 4062
rect 1344 3946 40656 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 40656 3946
rect 1344 3860 40656 3894
rect 25566 3666 25618 3678
rect 25566 3602 25618 3614
rect 17042 3502 17054 3554
rect 17106 3502 17118 3554
rect 24546 3502 24558 3554
rect 24610 3502 24622 3554
rect 18062 3330 18114 3342
rect 18062 3266 18114 3278
rect 1344 3162 40656 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 40656 3162
rect 1344 3076 40656 3110
<< via1 >>
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 18622 38222 18674 38274
rect 22430 38222 22482 38274
rect 25566 38222 25618 38274
rect 27470 38222 27522 38274
rect 17614 37998 17666 38050
rect 21758 37998 21810 38050
rect 24558 37998 24610 38050
rect 5630 37886 5682 37938
rect 34526 37886 34578 37938
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 18398 37438 18450 37490
rect 22094 37438 22146 37490
rect 26238 37438 26290 37490
rect 17390 37214 17442 37266
rect 21086 37214 21138 37266
rect 25230 37214 25282 37266
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 17390 36654 17442 36706
rect 16382 36430 16434 36482
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 1710 31054 1762 31106
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 16270 28030 16322 28082
rect 16606 28030 16658 28082
rect 15934 27918 15986 27970
rect 19742 27806 19794 27858
rect 20526 27694 20578 27746
rect 22654 27694 22706 27746
rect 23214 27694 23266 27746
rect 15822 27582 15874 27634
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 18510 27134 18562 27186
rect 21646 27134 21698 27186
rect 25230 27134 25282 27186
rect 15710 27022 15762 27074
rect 22318 27022 22370 27074
rect 16382 26910 16434 26962
rect 21310 26910 21362 26962
rect 21534 26910 21586 26962
rect 23102 26910 23154 26962
rect 25678 26910 25730 26962
rect 18958 26798 19010 26850
rect 21758 26798 21810 26850
rect 21870 26798 21922 26850
rect 40238 26798 40290 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 17614 26462 17666 26514
rect 22766 26462 22818 26514
rect 23550 26462 23602 26514
rect 24110 26462 24162 26514
rect 17838 26350 17890 26402
rect 22990 26350 23042 26402
rect 13806 26238 13858 26290
rect 17390 26238 17442 26290
rect 18622 26238 18674 26290
rect 19630 26238 19682 26290
rect 23102 26238 23154 26290
rect 23886 26238 23938 26290
rect 24222 26238 24274 26290
rect 14478 26126 14530 26178
rect 16606 26126 16658 26178
rect 17502 26126 17554 26178
rect 18510 26126 18562 26178
rect 20302 26126 20354 26178
rect 22430 26126 22482 26178
rect 18286 26014 18338 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 20638 25678 20690 25730
rect 20862 25678 20914 25730
rect 22430 25678 22482 25730
rect 22542 25566 22594 25618
rect 27470 25566 27522 25618
rect 27918 25566 27970 25618
rect 40014 25566 40066 25618
rect 15598 25454 15650 25506
rect 15822 25454 15874 25506
rect 16270 25454 16322 25506
rect 21198 25454 21250 25506
rect 22094 25454 22146 25506
rect 24558 25454 24610 25506
rect 37662 25454 37714 25506
rect 21534 25342 21586 25394
rect 21758 25342 21810 25394
rect 25342 25342 25394 25394
rect 15934 25230 15986 25282
rect 16830 25230 16882 25282
rect 21422 25230 21474 25282
rect 21982 25230 22034 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 21758 24894 21810 24946
rect 23662 24894 23714 24946
rect 25566 24894 25618 24946
rect 21422 24782 21474 24834
rect 21534 24782 21586 24834
rect 25678 24782 25730 24834
rect 26462 24782 26514 24834
rect 4286 24670 4338 24722
rect 23886 24670 23938 24722
rect 25230 24670 25282 24722
rect 25454 24670 25506 24722
rect 25790 24670 25842 24722
rect 1934 24446 1986 24498
rect 26350 24446 26402 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 1934 23998 1986 24050
rect 13470 23998 13522 24050
rect 17838 23998 17890 24050
rect 4286 23886 4338 23938
rect 14926 23886 14978 23938
rect 18398 23886 18450 23938
rect 13806 23774 13858 23826
rect 15710 23774 15762 23826
rect 13582 23662 13634 23714
rect 18062 23662 18114 23714
rect 18286 23662 18338 23714
rect 18846 23662 18898 23714
rect 24222 23662 24274 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 15038 23326 15090 23378
rect 16270 23326 16322 23378
rect 16606 23326 16658 23378
rect 24334 23214 24386 23266
rect 24446 23214 24498 23266
rect 4286 23102 4338 23154
rect 14702 23102 14754 23154
rect 15262 23102 15314 23154
rect 15710 23102 15762 23154
rect 16158 23102 16210 23154
rect 16382 23102 16434 23154
rect 17838 23102 17890 23154
rect 21198 23102 21250 23154
rect 24670 23102 24722 23154
rect 37662 23102 37714 23154
rect 11790 22990 11842 23042
rect 13918 22990 13970 23042
rect 15150 22990 15202 23042
rect 17502 22990 17554 23042
rect 18622 22990 18674 23042
rect 20750 22990 20802 23042
rect 21870 22990 21922 23042
rect 23998 22990 24050 23042
rect 1934 22878 1986 22930
rect 40014 22878 40066 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 14030 22542 14082 22594
rect 14366 22542 14418 22594
rect 14702 22542 14754 22594
rect 13806 22430 13858 22482
rect 15150 22430 15202 22482
rect 17838 22430 17890 22482
rect 21646 22430 21698 22482
rect 23214 22430 23266 22482
rect 40014 22430 40066 22482
rect 13694 22318 13746 22370
rect 17614 22318 17666 22370
rect 19742 22318 19794 22370
rect 20302 22318 20354 22370
rect 20862 22318 20914 22370
rect 22990 22318 23042 22370
rect 26126 22318 26178 22370
rect 37886 22318 37938 22370
rect 16942 22206 16994 22258
rect 17950 22206 18002 22258
rect 18286 22206 18338 22258
rect 18958 22206 19010 22258
rect 19854 22206 19906 22258
rect 20078 22206 20130 22258
rect 21310 22206 21362 22258
rect 21534 22206 21586 22258
rect 25342 22206 25394 22258
rect 28142 22206 28194 22258
rect 14478 22094 14530 22146
rect 17278 22094 17330 22146
rect 18622 22094 18674 22146
rect 19294 22094 19346 22146
rect 20526 22094 20578 22146
rect 20750 22094 20802 22146
rect 21758 22094 21810 22146
rect 21870 22094 21922 22146
rect 22318 22094 22370 22146
rect 22430 22094 22482 22146
rect 22542 22094 22594 22146
rect 26574 22094 26626 22146
rect 28030 22094 28082 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 14478 21758 14530 21810
rect 17838 21758 17890 21810
rect 17950 21758 18002 21810
rect 18286 21758 18338 21810
rect 25342 21758 25394 21810
rect 25678 21758 25730 21810
rect 13246 21646 13298 21698
rect 14926 21646 14978 21698
rect 14030 21534 14082 21586
rect 15038 21534 15090 21586
rect 17278 21534 17330 21586
rect 17726 21534 17778 21586
rect 18846 21534 18898 21586
rect 19182 21534 19234 21586
rect 25230 21534 25282 21586
rect 25454 21534 25506 21586
rect 26238 21534 26290 21586
rect 37662 21534 37714 21586
rect 11118 21422 11170 21474
rect 18398 21422 18450 21474
rect 23102 21422 23154 21474
rect 26910 21422 26962 21474
rect 29038 21422 29090 21474
rect 29486 21422 29538 21474
rect 29934 21422 29986 21474
rect 40014 21422 40066 21474
rect 14926 21310 14978 21362
rect 29374 21310 29426 21362
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 17502 20862 17554 20914
rect 21982 20862 22034 20914
rect 29710 20862 29762 20914
rect 40014 20862 40066 20914
rect 14478 20750 14530 20802
rect 20078 20750 20130 20802
rect 21422 20750 21474 20802
rect 22430 20750 22482 20802
rect 23102 20750 23154 20802
rect 29262 20750 29314 20802
rect 29934 20750 29986 20802
rect 30158 20750 30210 20802
rect 30606 20750 30658 20802
rect 37662 20750 37714 20802
rect 21982 20638 22034 20690
rect 26574 20638 26626 20690
rect 14142 20526 14194 20578
rect 21534 20526 21586 20578
rect 21758 20526 21810 20578
rect 22206 20526 22258 20578
rect 29374 20526 29426 20578
rect 29486 20526 29538 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 18062 20190 18114 20242
rect 26126 20190 26178 20242
rect 15150 20078 15202 20130
rect 15374 20078 15426 20130
rect 16270 20078 16322 20130
rect 16382 20078 16434 20130
rect 17390 20078 17442 20130
rect 18174 20078 18226 20130
rect 19406 20078 19458 20130
rect 20414 20078 20466 20130
rect 20638 20078 20690 20130
rect 23102 20078 23154 20130
rect 24670 20078 24722 20130
rect 26014 20078 26066 20130
rect 26238 20078 26290 20130
rect 27470 20078 27522 20130
rect 30046 20078 30098 20130
rect 11230 19966 11282 20018
rect 15486 19966 15538 20018
rect 16606 19966 16658 20018
rect 16942 19966 16994 20018
rect 17614 19966 17666 20018
rect 20302 19966 20354 20018
rect 22766 19966 22818 20018
rect 24446 19966 24498 20018
rect 25566 19966 25618 20018
rect 26686 19966 26738 20018
rect 11902 19854 11954 19906
rect 14030 19854 14082 19906
rect 14702 19854 14754 19906
rect 14926 19854 14978 19906
rect 19966 19854 20018 19906
rect 25790 19854 25842 19906
rect 29598 19854 29650 19906
rect 14366 19742 14418 19794
rect 19630 19742 19682 19794
rect 25342 19742 25394 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 18062 19406 18114 19458
rect 14254 19294 14306 19346
rect 17502 19294 17554 19346
rect 21422 19294 21474 19346
rect 25006 19294 25058 19346
rect 25902 19294 25954 19346
rect 12686 19182 12738 19234
rect 15934 19182 15986 19234
rect 16382 19182 16434 19234
rect 17278 19182 17330 19234
rect 18062 19182 18114 19234
rect 21870 19182 21922 19234
rect 22206 19182 22258 19234
rect 23214 19182 23266 19234
rect 12350 19070 12402 19122
rect 14926 19070 14978 19122
rect 15262 19070 15314 19122
rect 16606 19070 16658 19122
rect 18398 19070 18450 19122
rect 20414 19070 20466 19122
rect 22878 19070 22930 19122
rect 16158 18958 16210 19010
rect 16942 18958 16994 19010
rect 20750 18958 20802 19010
rect 21758 18958 21810 19010
rect 22990 18958 23042 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 15262 18622 15314 18674
rect 20078 18622 20130 18674
rect 20862 18622 20914 18674
rect 21534 18622 21586 18674
rect 22654 18622 22706 18674
rect 22990 18622 23042 18674
rect 23438 18622 23490 18674
rect 26910 18622 26962 18674
rect 14926 18510 14978 18562
rect 15598 18510 15650 18562
rect 15710 18510 15762 18562
rect 21982 18510 22034 18562
rect 23550 18510 23602 18562
rect 15934 18398 15986 18450
rect 16158 18398 16210 18450
rect 18174 18398 18226 18450
rect 18286 18398 18338 18450
rect 18510 18398 18562 18450
rect 19406 18398 19458 18450
rect 19742 18398 19794 18450
rect 20526 18398 20578 18450
rect 21198 18398 21250 18450
rect 22318 18398 22370 18450
rect 23886 18398 23938 18450
rect 25230 18398 25282 18450
rect 25454 18398 25506 18450
rect 25790 18398 25842 18450
rect 26238 18398 26290 18450
rect 27134 18398 27186 18450
rect 37662 18398 37714 18450
rect 19070 18286 19122 18338
rect 25342 18286 25394 18338
rect 26686 18286 26738 18338
rect 27022 18286 27074 18338
rect 16158 18174 16210 18226
rect 17726 18174 17778 18226
rect 23438 18174 23490 18226
rect 23998 18174 24050 18226
rect 26462 18174 26514 18226
rect 40014 18174 40066 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 16270 17838 16322 17890
rect 22654 17838 22706 17890
rect 24222 17838 24274 17890
rect 27694 17838 27746 17890
rect 28142 17838 28194 17890
rect 28366 17838 28418 17890
rect 1934 17726 1986 17778
rect 22990 17726 23042 17778
rect 27470 17726 27522 17778
rect 27918 17726 27970 17778
rect 40014 17726 40066 17778
rect 4286 17614 4338 17666
rect 13694 17614 13746 17666
rect 14366 17614 14418 17666
rect 14702 17614 14754 17666
rect 18622 17614 18674 17666
rect 21982 17614 22034 17666
rect 23550 17614 23602 17666
rect 23886 17614 23938 17666
rect 24670 17614 24722 17666
rect 28478 17614 28530 17666
rect 37662 17614 37714 17666
rect 14590 17502 14642 17554
rect 16046 17502 16098 17554
rect 17390 17502 17442 17554
rect 17726 17502 17778 17554
rect 18062 17502 18114 17554
rect 18286 17502 18338 17554
rect 18846 17502 18898 17554
rect 18958 17502 19010 17554
rect 19742 17502 19794 17554
rect 22878 17502 22930 17554
rect 23662 17502 23714 17554
rect 25342 17502 25394 17554
rect 13918 17390 13970 17442
rect 14142 17390 14194 17442
rect 14254 17390 14306 17442
rect 15150 17390 15202 17442
rect 16158 17390 16210 17442
rect 16606 17390 16658 17442
rect 16942 17390 16994 17442
rect 18174 17390 18226 17442
rect 19406 17390 19458 17442
rect 21758 17390 21810 17442
rect 21870 17390 21922 17442
rect 23774 17390 23826 17442
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 17838 17054 17890 17106
rect 19742 17054 19794 17106
rect 20414 17054 20466 17106
rect 23326 17054 23378 17106
rect 29822 17054 29874 17106
rect 13022 16942 13074 16994
rect 21758 16942 21810 16994
rect 27246 16942 27298 16994
rect 12238 16830 12290 16882
rect 17390 16830 17442 16882
rect 17614 16830 17666 16882
rect 17950 16830 18002 16882
rect 19182 16830 19234 16882
rect 19406 16830 19458 16882
rect 21982 16830 22034 16882
rect 22318 16830 22370 16882
rect 22654 16830 22706 16882
rect 22878 16830 22930 16882
rect 23550 16830 23602 16882
rect 26462 16830 26514 16882
rect 15150 16718 15202 16770
rect 15598 16718 15650 16770
rect 17502 16718 17554 16770
rect 18846 16718 18898 16770
rect 20190 16718 20242 16770
rect 21870 16718 21922 16770
rect 23102 16718 23154 16770
rect 23438 16718 23490 16770
rect 29374 16718 29426 16770
rect 20526 16606 20578 16658
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 21310 16270 21362 16322
rect 21646 16270 21698 16322
rect 22990 16270 23042 16322
rect 23326 16270 23378 16322
rect 13470 16158 13522 16210
rect 15598 16158 15650 16210
rect 22766 16158 22818 16210
rect 23214 16158 23266 16210
rect 16270 16046 16322 16098
rect 16942 16046 16994 16098
rect 17278 16046 17330 16098
rect 19294 16046 19346 16098
rect 21310 16046 21362 16098
rect 19070 15934 19122 15986
rect 17054 15822 17106 15874
rect 17614 15822 17666 15874
rect 22878 15822 22930 15874
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 25230 15486 25282 15538
rect 14702 15374 14754 15426
rect 19854 15374 19906 15426
rect 19966 15374 20018 15426
rect 20862 15374 20914 15426
rect 21198 15374 21250 15426
rect 21534 15374 21586 15426
rect 22766 15374 22818 15426
rect 14030 15262 14082 15314
rect 22990 15262 23042 15314
rect 16830 15150 16882 15202
rect 17502 15150 17554 15202
rect 20638 15150 20690 15202
rect 25342 15150 25394 15202
rect 20302 15038 20354 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 16942 14590 16994 14642
rect 19070 14590 19122 14642
rect 19518 14590 19570 14642
rect 23550 14590 23602 14642
rect 25678 14590 25730 14642
rect 26126 14590 26178 14642
rect 16270 14478 16322 14530
rect 20190 14478 20242 14530
rect 22878 14478 22930 14530
rect 20414 14254 20466 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 25342 13918 25394 13970
rect 20638 13806 20690 13858
rect 22542 13806 22594 13858
rect 21422 13694 21474 13746
rect 21870 13694 21922 13746
rect 18510 13582 18562 13634
rect 24670 13582 24722 13634
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 21758 13022 21810 13074
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 25230 4286 25282 4338
rect 26238 4062 26290 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 25566 3614 25618 3666
rect 17054 3502 17106 3554
rect 24558 3502 24610 3554
rect 18062 3278 18114 3330
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 5376 41200 5488 42000
rect 16128 41200 16240 42000
rect 16800 41200 16912 42000
rect 18144 41200 18256 42000
rect 20832 41200 20944 42000
rect 22176 41200 22288 42000
rect 22848 41200 22960 42000
rect 24864 41200 24976 42000
rect 26208 41200 26320 42000
rect 34272 41200 34384 42000
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 5404 37940 5460 41200
rect 5628 37940 5684 37950
rect 5404 37938 5684 37940
rect 5404 37886 5630 37938
rect 5682 37886 5684 37938
rect 5404 37884 5684 37886
rect 5628 37874 5684 37884
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 16156 36708 16212 41200
rect 16828 37492 16884 41200
rect 18172 38276 18228 41200
rect 18620 38276 18676 38286
rect 18172 38274 18676 38276
rect 18172 38222 18622 38274
rect 18674 38222 18676 38274
rect 18172 38220 18676 38222
rect 18620 38210 18676 38220
rect 16828 37426 16884 37436
rect 17612 38050 17668 38062
rect 17612 37998 17614 38050
rect 17666 37998 17668 38050
rect 17388 37268 17444 37278
rect 16156 36642 16212 36652
rect 17276 37266 17444 37268
rect 17276 37214 17390 37266
rect 17442 37214 17444 37266
rect 17276 37212 17444 37214
rect 16380 36482 16436 36494
rect 16380 36430 16382 36482
rect 16434 36430 16436 36482
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 16380 31948 16436 36430
rect 16268 31892 16436 31948
rect 1708 31106 1764 31118
rect 1708 31054 1710 31106
rect 1762 31054 1764 31106
rect 1708 30324 1764 31054
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 1708 30258 1764 30268
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 16268 28084 16324 31892
rect 16604 28084 16660 28094
rect 15932 28082 16548 28084
rect 15932 28030 16270 28082
rect 16322 28030 16548 28082
rect 15932 28028 16548 28030
rect 15932 27970 15988 28028
rect 16268 28018 16324 28028
rect 15932 27918 15934 27970
rect 15986 27918 15988 27970
rect 15932 27906 15988 27918
rect 15820 27634 15876 27646
rect 15820 27582 15822 27634
rect 15874 27582 15876 27634
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 15708 27074 15764 27086
rect 15708 27022 15710 27074
rect 15762 27022 15764 27074
rect 4172 26964 4228 26974
rect 1932 24500 1988 24510
rect 1932 24406 1988 24444
rect 1932 24050 1988 24062
rect 1932 23998 1934 24050
rect 1986 23998 1988 24050
rect 1932 23604 1988 23998
rect 1932 23538 1988 23548
rect 1932 22932 1988 22942
rect 1932 22838 1988 22876
rect 4172 21476 4228 26908
rect 13804 26290 13860 26302
rect 13804 26238 13806 26290
rect 13858 26238 13860 26290
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 13804 25284 13860 26238
rect 15596 26292 15652 26302
rect 14476 26180 14532 26190
rect 14476 26086 14532 26124
rect 15596 25508 15652 26236
rect 15148 25506 15652 25508
rect 15148 25454 15598 25506
rect 15650 25454 15652 25506
rect 15148 25452 15652 25454
rect 15036 25284 15092 25294
rect 13804 25218 13860 25228
rect 14924 25228 15036 25284
rect 4284 24724 4340 24734
rect 4284 24630 4340 24668
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 13468 24050 13524 24062
rect 13468 23998 13470 24050
rect 13522 23998 13524 24050
rect 4284 23940 4340 23950
rect 4284 23846 4340 23884
rect 11116 23940 11172 23950
rect 4284 23156 4340 23166
rect 4284 23062 4340 23100
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 4172 21410 4228 21420
rect 11116 22372 11172 23884
rect 11788 23156 11844 23166
rect 11788 23042 11844 23100
rect 11788 22990 11790 23042
rect 11842 22990 11844 23042
rect 11788 22978 11844 22990
rect 13468 22596 13524 23998
rect 14924 23940 14980 25228
rect 15036 25218 15092 25228
rect 15148 23940 15204 25452
rect 15596 25442 15652 25452
rect 15708 25284 15764 27022
rect 15820 25506 15876 27582
rect 16380 26962 16436 26974
rect 16380 26910 16382 26962
rect 16434 26910 16436 26962
rect 16268 26404 16324 26414
rect 15820 25454 15822 25506
rect 15874 25454 15876 25506
rect 15820 25442 15876 25454
rect 15932 26180 15988 26190
rect 15708 25218 15764 25228
rect 15932 25282 15988 26124
rect 16268 25508 16324 26348
rect 16380 26180 16436 26910
rect 16492 26908 16548 28028
rect 16604 27990 16660 28028
rect 17276 28084 17332 37212
rect 17388 37202 17444 37212
rect 17388 36708 17444 36718
rect 17388 36614 17444 36652
rect 17276 28018 17332 28028
rect 17612 27188 17668 37998
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 18396 37492 18452 37502
rect 18396 37398 18452 37436
rect 20860 37492 20916 41200
rect 22204 38276 22260 41200
rect 22428 38276 22484 38286
rect 22204 38274 22484 38276
rect 22204 38222 22430 38274
rect 22482 38222 22484 38274
rect 22204 38220 22484 38222
rect 22428 38210 22484 38220
rect 22876 38276 22932 41200
rect 22876 38210 22932 38220
rect 21756 38052 21812 38062
rect 21756 37958 21812 37996
rect 22428 38052 22484 38062
rect 20860 37426 20916 37436
rect 22092 37492 22148 37502
rect 22092 37398 22148 37436
rect 21084 37266 21140 37278
rect 21084 37214 21086 37266
rect 21138 37214 21140 37266
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 21084 31948 21140 37214
rect 20748 31892 21140 31948
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 19740 27860 19796 27870
rect 19628 27858 19796 27860
rect 19628 27806 19742 27858
rect 19794 27806 19796 27858
rect 19628 27804 19796 27806
rect 16492 26852 16660 26908
rect 16380 26114 16436 26124
rect 16604 26178 16660 26852
rect 17612 26514 17668 27132
rect 18508 27188 18564 27198
rect 18508 27094 18564 27132
rect 19628 27076 19684 27804
rect 19740 27794 19796 27804
rect 20524 27748 20580 27758
rect 20524 27654 20580 27692
rect 17612 26462 17614 26514
rect 17666 26462 17668 26514
rect 17612 26450 17668 26462
rect 18956 26850 19012 26862
rect 18956 26798 18958 26850
rect 19010 26798 19012 26850
rect 17836 26404 17892 26414
rect 17836 26310 17892 26348
rect 17388 26292 17444 26302
rect 17388 26198 17444 26236
rect 18620 26290 18676 26302
rect 18620 26238 18622 26290
rect 18674 26238 18676 26290
rect 16604 26126 16606 26178
rect 16658 26126 16660 26178
rect 16604 26114 16660 26126
rect 17500 26180 17556 26190
rect 18508 26180 18564 26190
rect 17500 26178 17892 26180
rect 17500 26126 17502 26178
rect 17554 26126 17892 26178
rect 17500 26124 17892 26126
rect 17500 26114 17556 26124
rect 17836 26068 17892 26124
rect 18508 26086 18564 26124
rect 18284 26068 18340 26078
rect 17836 26066 18340 26068
rect 17836 26014 18286 26066
rect 18338 26014 18340 26066
rect 17836 26012 18340 26014
rect 18284 26002 18340 26012
rect 17164 25956 17220 25966
rect 16268 25506 16436 25508
rect 16268 25454 16270 25506
rect 16322 25454 16436 25506
rect 16268 25452 16436 25454
rect 16268 25442 16324 25452
rect 15932 25230 15934 25282
rect 15986 25230 15988 25282
rect 15932 25218 15988 25230
rect 14700 23938 14980 23940
rect 14700 23886 14926 23938
rect 14978 23886 14980 23938
rect 14700 23884 14980 23886
rect 13804 23826 13860 23838
rect 13804 23774 13806 23826
rect 13858 23774 13860 23826
rect 11116 21474 11172 22316
rect 13244 22540 13524 22596
rect 13580 23714 13636 23726
rect 13580 23662 13582 23714
rect 13634 23662 13636 23714
rect 13244 21698 13300 22540
rect 13244 21646 13246 21698
rect 13298 21646 13300 21698
rect 13244 21634 13300 21646
rect 11116 21422 11118 21474
rect 11170 21422 11172 21474
rect 11116 21410 11172 21422
rect 13580 21364 13636 23662
rect 13804 22482 13860 23774
rect 14588 23380 14644 23390
rect 13916 23044 13972 23054
rect 13916 23042 14420 23044
rect 13916 22990 13918 23042
rect 13970 22990 14420 23042
rect 13916 22988 14420 22990
rect 13916 22978 13972 22988
rect 14028 22596 14084 22606
rect 14028 22502 14084 22540
rect 14364 22594 14420 22988
rect 14364 22542 14366 22594
rect 14418 22542 14420 22594
rect 14364 22530 14420 22542
rect 14588 22596 14644 23324
rect 14700 23156 14756 23884
rect 14924 23874 14980 23884
rect 15036 23884 15204 23940
rect 15036 23380 15092 23884
rect 15708 23828 15764 23838
rect 15708 23826 16324 23828
rect 15708 23774 15710 23826
rect 15762 23774 16324 23826
rect 15708 23772 16324 23774
rect 15708 23762 15764 23772
rect 15036 23286 15092 23324
rect 16268 23378 16324 23772
rect 16268 23326 16270 23378
rect 16322 23326 16324 23378
rect 16268 23314 16324 23326
rect 15260 23156 15316 23166
rect 14700 23154 15092 23156
rect 14700 23102 14702 23154
rect 14754 23102 15092 23154
rect 14700 23100 15092 23102
rect 14700 23090 14756 23100
rect 14588 22530 14644 22540
rect 14700 22932 14756 22942
rect 14700 22594 14756 22876
rect 14700 22542 14702 22594
rect 14754 22542 14756 22594
rect 14700 22530 14756 22542
rect 13804 22430 13806 22482
rect 13858 22430 13860 22482
rect 13804 22418 13860 22430
rect 13692 22372 13748 22382
rect 13692 22278 13748 22316
rect 14476 22148 14532 22158
rect 14476 22054 14532 22092
rect 14476 21812 14532 21822
rect 14812 21812 14868 23100
rect 15036 22484 15092 23100
rect 15260 23062 15316 23100
rect 15708 23154 15764 23166
rect 15708 23102 15710 23154
rect 15762 23102 15764 23154
rect 15148 23044 15204 23054
rect 15148 22950 15204 22988
rect 15148 22484 15204 22494
rect 15036 22482 15204 22484
rect 15036 22430 15150 22482
rect 15202 22430 15204 22482
rect 15036 22428 15204 22430
rect 15148 22418 15204 22428
rect 14028 21810 14868 21812
rect 14028 21758 14478 21810
rect 14530 21758 14868 21810
rect 14028 21756 14868 21758
rect 15484 22148 15540 22158
rect 14028 21586 14084 21756
rect 14028 21534 14030 21586
rect 14082 21534 14084 21586
rect 14028 21522 14084 21534
rect 13580 21298 13636 21308
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 14140 20578 14196 20590
rect 14140 20526 14142 20578
rect 14194 20526 14196 20578
rect 11228 20020 11284 20030
rect 11228 19926 11284 19964
rect 11676 20020 11732 20030
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 11676 18452 11732 19964
rect 11900 19908 11956 19918
rect 11900 19906 12404 19908
rect 11900 19854 11902 19906
rect 11954 19854 12404 19906
rect 11900 19852 12404 19854
rect 11900 19842 11956 19852
rect 12348 19122 12404 19852
rect 14028 19906 14084 19918
rect 14028 19854 14030 19906
rect 14082 19854 14084 19906
rect 12684 19796 12740 19806
rect 12684 19234 12740 19740
rect 12684 19182 12686 19234
rect 12738 19182 12740 19234
rect 12684 19170 12740 19182
rect 12348 19070 12350 19122
rect 12402 19070 12404 19122
rect 12348 19058 12404 19070
rect 14028 19124 14084 19854
rect 14140 19348 14196 20526
rect 14140 19282 14196 19292
rect 14252 20020 14308 21756
rect 14476 21746 14532 21756
rect 14924 21700 14980 21710
rect 14588 21698 14980 21700
rect 14588 21646 14926 21698
rect 14978 21646 14980 21698
rect 14588 21644 14980 21646
rect 14476 20804 14532 20814
rect 14588 20804 14644 21644
rect 14924 21634 14980 21644
rect 15036 21586 15092 21598
rect 15036 21534 15038 21586
rect 15090 21534 15092 21586
rect 14700 21364 14756 21374
rect 14924 21364 14980 21374
rect 14756 21362 14980 21364
rect 14756 21310 14926 21362
rect 14978 21310 14980 21362
rect 14756 21308 14980 21310
rect 14700 21298 14756 21308
rect 14924 21298 14980 21308
rect 14476 20802 14644 20804
rect 14476 20750 14478 20802
rect 14530 20750 14644 20802
rect 14476 20748 14644 20750
rect 14476 20132 14532 20748
rect 14476 20066 14532 20076
rect 14252 19346 14308 19964
rect 14700 19908 14756 19918
rect 14700 19814 14756 19852
rect 14924 19908 14980 19918
rect 15036 19908 15092 21534
rect 15148 20132 15204 20142
rect 15372 20132 15428 20142
rect 15148 20038 15204 20076
rect 15260 20130 15428 20132
rect 15260 20078 15374 20130
rect 15426 20078 15428 20130
rect 15260 20076 15428 20078
rect 14924 19906 15092 19908
rect 14924 19854 14926 19906
rect 14978 19854 15092 19906
rect 14924 19852 15092 19854
rect 14924 19842 14980 19852
rect 14364 19796 14420 19806
rect 14364 19702 14420 19740
rect 14252 19294 14254 19346
rect 14306 19294 14308 19346
rect 14252 19282 14308 19294
rect 14028 19058 14084 19068
rect 14924 19124 14980 19134
rect 14924 19030 14980 19068
rect 13020 18564 13076 18574
rect 11676 18396 12292 18452
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 1932 17778 1988 17790
rect 1932 17726 1934 17778
rect 1986 17726 1988 17778
rect 1932 16884 1988 17726
rect 4284 17668 4340 17678
rect 4284 17574 4340 17612
rect 1932 16818 1988 16828
rect 12236 16882 12292 18396
rect 13020 16994 13076 18508
rect 14924 18562 14980 18574
rect 14924 18510 14926 18562
rect 14978 18510 14980 18562
rect 14924 18340 14980 18510
rect 14700 18284 14924 18340
rect 13020 16942 13022 16994
rect 13074 16942 13076 16994
rect 13020 16930 13076 16942
rect 13468 17668 13524 17678
rect 12236 16830 12238 16882
rect 12290 16830 12292 16882
rect 12236 16772 12292 16830
rect 12236 16706 12292 16716
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 13468 16210 13524 17612
rect 13692 17668 13748 17678
rect 14364 17668 14420 17678
rect 13692 17666 14420 17668
rect 13692 17614 13694 17666
rect 13746 17614 14366 17666
rect 14418 17614 14420 17666
rect 13692 17612 14420 17614
rect 13692 17602 13748 17612
rect 14364 17602 14420 17612
rect 14588 17668 14644 17678
rect 14588 17554 14644 17612
rect 14700 17666 14756 18284
rect 14924 18274 14980 18284
rect 14700 17614 14702 17666
rect 14754 17614 14756 17666
rect 14700 17602 14756 17614
rect 14588 17502 14590 17554
rect 14642 17502 14644 17554
rect 14588 17490 14644 17502
rect 13916 17444 13972 17454
rect 13916 17350 13972 17388
rect 14140 17442 14196 17454
rect 14140 17390 14142 17442
rect 14194 17390 14196 17442
rect 14140 17332 14196 17390
rect 14140 17266 14196 17276
rect 14252 17442 14308 17454
rect 14252 17390 14254 17442
rect 14306 17390 14308 17442
rect 13468 16158 13470 16210
rect 13522 16158 13524 16210
rect 13468 16146 13524 16158
rect 14028 16772 14084 16782
rect 14028 15314 14084 16716
rect 14252 16212 14308 17390
rect 14924 17444 14980 17454
rect 15036 17444 15092 19852
rect 14980 17388 15092 17444
rect 15148 19348 15204 19358
rect 15148 17444 15204 19292
rect 15260 19236 15316 20076
rect 15372 20066 15428 20076
rect 15484 20020 15540 22092
rect 15708 21812 15764 23102
rect 15708 21746 15764 21756
rect 16156 23154 16212 23166
rect 16156 23102 16158 23154
rect 16210 23102 16212 23154
rect 16156 20132 16212 23102
rect 16380 23154 16436 25452
rect 16828 25284 16884 25294
rect 16604 23716 16660 23726
rect 16604 23378 16660 23660
rect 16604 23326 16606 23378
rect 16658 23326 16660 23378
rect 16604 23314 16660 23326
rect 16380 23102 16382 23154
rect 16434 23102 16436 23154
rect 16380 22372 16436 23102
rect 16828 23156 16884 25228
rect 16828 23090 16884 23100
rect 16940 23380 16996 23390
rect 16380 22306 16436 22316
rect 16940 22258 16996 23324
rect 16940 22206 16942 22258
rect 16994 22206 16996 22258
rect 16940 22194 16996 22206
rect 16268 20132 16324 20142
rect 16212 20130 16324 20132
rect 16212 20078 16270 20130
rect 16322 20078 16324 20130
rect 16212 20076 16324 20078
rect 16156 20038 16212 20076
rect 16268 20066 16324 20076
rect 16380 20130 16436 20142
rect 16380 20078 16382 20130
rect 16434 20078 16436 20130
rect 15484 20018 15652 20020
rect 15484 19966 15486 20018
rect 15538 19966 15652 20018
rect 15484 19964 15652 19966
rect 15484 19954 15540 19964
rect 15260 19122 15316 19180
rect 15260 19070 15262 19122
rect 15314 19070 15316 19122
rect 15260 18674 15316 19070
rect 15260 18622 15262 18674
rect 15314 18622 15316 18674
rect 15260 18610 15316 18622
rect 15596 18676 15652 19964
rect 15932 19796 15988 19806
rect 15932 19234 15988 19740
rect 15932 19182 15934 19234
rect 15986 19182 15988 19234
rect 15932 19170 15988 19182
rect 16380 19234 16436 20078
rect 16604 20020 16660 20030
rect 16604 19926 16660 19964
rect 16940 20018 16996 20030
rect 16940 19966 16942 20018
rect 16994 19966 16996 20018
rect 16380 19182 16382 19234
rect 16434 19182 16436 19234
rect 15596 18562 15652 18620
rect 16156 19010 16212 19022
rect 16156 18958 16158 19010
rect 16210 18958 16212 19010
rect 15596 18510 15598 18562
rect 15650 18510 15652 18562
rect 15596 18498 15652 18510
rect 15708 18564 15764 18574
rect 15708 18470 15764 18508
rect 15932 18450 15988 18462
rect 15932 18398 15934 18450
rect 15986 18398 15988 18450
rect 15932 18340 15988 18398
rect 16156 18450 16212 18958
rect 16156 18398 16158 18450
rect 16210 18398 16212 18450
rect 16156 18386 16212 18398
rect 15148 17442 15316 17444
rect 15148 17390 15150 17442
rect 15202 17390 15316 17442
rect 15148 17388 15316 17390
rect 14924 17378 14980 17388
rect 15148 17378 15204 17388
rect 15260 17332 15316 17388
rect 15260 17266 15316 17276
rect 15148 17220 15204 17230
rect 15148 16770 15204 17164
rect 15932 16884 15988 18284
rect 16156 18228 16212 18238
rect 16156 18134 16212 18172
rect 16268 18004 16324 18014
rect 16268 17890 16324 17948
rect 16268 17838 16270 17890
rect 16322 17838 16324 17890
rect 16268 17826 16324 17838
rect 16044 17668 16100 17678
rect 16044 17554 16100 17612
rect 16044 17502 16046 17554
rect 16098 17502 16100 17554
rect 16044 17490 16100 17502
rect 16380 17556 16436 19182
rect 16940 19236 16996 19966
rect 17164 19572 17220 25900
rect 18508 25956 18564 25966
rect 18620 25956 18676 26238
rect 18564 25900 18676 25956
rect 18508 25890 18564 25900
rect 17836 24724 17892 24734
rect 17836 24050 17892 24668
rect 17836 23998 17838 24050
rect 17890 23998 17892 24050
rect 17836 23604 17892 23998
rect 18396 23940 18452 23950
rect 17836 23538 17892 23548
rect 17948 23938 18452 23940
rect 17948 23886 18398 23938
rect 18450 23886 18452 23938
rect 17948 23884 18452 23886
rect 17948 23380 18004 23884
rect 18396 23874 18452 23884
rect 18060 23716 18116 23726
rect 18060 23622 18116 23660
rect 18284 23714 18340 23726
rect 18284 23662 18286 23714
rect 18338 23662 18340 23714
rect 18284 23604 18340 23662
rect 18844 23716 18900 23726
rect 18956 23716 19012 26798
rect 19628 26290 19684 27020
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19628 26238 19630 26290
rect 19682 26238 19684 26290
rect 19628 26226 19684 26238
rect 20300 26180 20356 26190
rect 20300 26178 20692 26180
rect 20300 26126 20302 26178
rect 20354 26126 20692 26178
rect 20300 26124 20692 26126
rect 20300 26114 20356 26124
rect 20636 25730 20692 26124
rect 20636 25678 20638 25730
rect 20690 25678 20692 25730
rect 20636 25666 20692 25678
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 19836 25050 20100 25060
rect 18844 23714 19012 23716
rect 18844 23662 18846 23714
rect 18898 23662 19012 23714
rect 18844 23660 19012 23662
rect 20300 24836 20356 24846
rect 18844 23604 18900 23660
rect 18284 23538 18340 23548
rect 18396 23548 18900 23604
rect 19836 23548 20100 23558
rect 17836 23156 17892 23166
rect 17500 23044 17556 23054
rect 17836 23044 17892 23100
rect 17500 23042 17892 23044
rect 17500 22990 17502 23042
rect 17554 22990 17892 23042
rect 17500 22988 17892 22990
rect 17276 22148 17332 22158
rect 17276 21586 17332 22092
rect 17276 21534 17278 21586
rect 17330 21534 17332 21586
rect 17276 20244 17332 21534
rect 17500 20914 17556 22988
rect 17836 22484 17892 22494
rect 17948 22484 18004 23324
rect 18396 23156 18452 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 18396 23090 18452 23100
rect 17836 22482 18004 22484
rect 17836 22430 17838 22482
rect 17890 22430 18004 22482
rect 17836 22428 18004 22430
rect 18620 23042 18676 23054
rect 18620 22990 18622 23042
rect 18674 22990 18676 23042
rect 18620 22484 18676 22990
rect 17836 22418 17892 22428
rect 18620 22418 18676 22428
rect 19852 23044 19908 23054
rect 17612 22370 17668 22382
rect 17612 22318 17614 22370
rect 17666 22318 17668 22370
rect 17612 22148 17668 22318
rect 18284 22372 18340 22382
rect 17948 22260 18004 22270
rect 17948 22166 18004 22204
rect 18284 22258 18340 22316
rect 19740 22372 19796 22382
rect 19740 22278 19796 22316
rect 18284 22206 18286 22258
rect 18338 22206 18340 22258
rect 18284 22194 18340 22206
rect 18396 22260 18452 22270
rect 17612 22082 17668 22092
rect 17836 21812 17892 21822
rect 17836 21718 17892 21756
rect 17948 21812 18004 21822
rect 18172 21812 18228 21822
rect 17948 21810 18172 21812
rect 17948 21758 17950 21810
rect 18002 21758 18172 21810
rect 17948 21756 18172 21758
rect 17948 21746 18004 21756
rect 17500 20862 17502 20914
rect 17554 20862 17556 20914
rect 17500 20850 17556 20862
rect 17724 21586 17780 21598
rect 17724 21534 17726 21586
rect 17778 21534 17780 21586
rect 17724 20692 17780 21534
rect 17724 20626 17780 20636
rect 18172 20356 18228 21756
rect 18284 21812 18340 21822
rect 18396 21812 18452 22204
rect 18956 22260 19012 22270
rect 18956 22166 19012 22204
rect 19852 22258 19908 22988
rect 20300 22372 20356 24780
rect 20748 23044 20804 31892
rect 21644 27748 21700 27758
rect 21644 27186 21700 27692
rect 21644 27134 21646 27186
rect 21698 27134 21700 27186
rect 21644 27122 21700 27134
rect 22316 27076 22372 27086
rect 22316 26982 22372 27020
rect 21308 26962 21364 26974
rect 21308 26910 21310 26962
rect 21362 26910 21364 26962
rect 21308 25956 21364 26910
rect 21532 26964 21588 26974
rect 21532 26962 21700 26964
rect 21532 26910 21534 26962
rect 21586 26910 21700 26962
rect 21532 26908 21700 26910
rect 21532 26898 21588 26908
rect 21644 26404 21700 26908
rect 21644 25956 21700 26348
rect 21756 26850 21812 26862
rect 21756 26798 21758 26850
rect 21810 26798 21812 26850
rect 21756 26180 21812 26798
rect 21868 26852 21924 26862
rect 21868 26850 22148 26852
rect 21868 26798 21870 26850
rect 21922 26798 22148 26850
rect 21868 26796 22148 26798
rect 21868 26786 21924 26796
rect 21756 26114 21812 26124
rect 21644 25900 21924 25956
rect 21308 25890 21364 25900
rect 20860 25732 20916 25742
rect 20860 25730 21252 25732
rect 20860 25678 20862 25730
rect 20914 25678 21252 25730
rect 20860 25676 21252 25678
rect 20860 25666 20916 25676
rect 21196 25506 21252 25676
rect 21196 25454 21198 25506
rect 21250 25454 21252 25506
rect 21196 25442 21252 25454
rect 21532 25396 21588 25406
rect 21756 25396 21812 25406
rect 21532 25394 21812 25396
rect 21532 25342 21534 25394
rect 21586 25342 21758 25394
rect 21810 25342 21812 25394
rect 21532 25340 21812 25342
rect 21532 25330 21588 25340
rect 21756 25330 21812 25340
rect 21420 25284 21476 25294
rect 20748 22950 20804 22988
rect 21084 25282 21476 25284
rect 21084 25230 21422 25282
rect 21474 25230 21476 25282
rect 21084 25228 21476 25230
rect 20188 22370 20356 22372
rect 20188 22318 20302 22370
rect 20354 22318 20356 22370
rect 20188 22316 20356 22318
rect 19852 22206 19854 22258
rect 19906 22206 19908 22258
rect 19852 22194 19908 22206
rect 20076 22260 20132 22270
rect 20076 22166 20132 22204
rect 18284 21810 18452 21812
rect 18284 21758 18286 21810
rect 18338 21758 18452 21810
rect 18284 21756 18452 21758
rect 18620 22146 18676 22158
rect 18620 22094 18622 22146
rect 18674 22094 18676 22146
rect 18284 21746 18340 21756
rect 18396 21474 18452 21486
rect 18396 21422 18398 21474
rect 18450 21422 18452 21474
rect 18172 20300 18340 20356
rect 17276 20178 17332 20188
rect 18060 20244 18116 20254
rect 18060 20150 18116 20188
rect 17388 20132 17444 20142
rect 18172 20132 18228 20142
rect 17444 20076 17556 20132
rect 17388 20038 17444 20076
rect 17276 19572 17332 19582
rect 17164 19516 17276 19572
rect 17276 19506 17332 19516
rect 17500 19346 17556 20076
rect 18172 20038 18228 20076
rect 17500 19294 17502 19346
rect 17554 19294 17556 19346
rect 17500 19282 17556 19294
rect 17612 20018 17668 20030
rect 17612 19966 17614 20018
rect 17666 19966 17668 20018
rect 16940 19170 16996 19180
rect 17276 19234 17332 19246
rect 17276 19182 17278 19234
rect 17330 19182 17332 19234
rect 16604 19122 16660 19134
rect 16604 19070 16606 19122
rect 16658 19070 16660 19122
rect 16604 18116 16660 19070
rect 16604 18050 16660 18060
rect 16940 19010 16996 19022
rect 16940 18958 16942 19010
rect 16994 18958 16996 19010
rect 16940 17668 16996 18958
rect 17276 18228 17332 19182
rect 17276 18162 17332 18172
rect 17612 19124 17668 19966
rect 18284 20020 18340 20300
rect 18284 19954 18340 19964
rect 18172 19796 18228 19806
rect 18396 19796 18452 21422
rect 18228 19740 18452 19796
rect 18060 19572 18116 19582
rect 18060 19458 18116 19516
rect 18060 19406 18062 19458
rect 18114 19406 18116 19458
rect 18060 19394 18116 19406
rect 18060 19236 18116 19246
rect 18060 19142 18116 19180
rect 16940 17602 16996 17612
rect 17052 18116 17108 18126
rect 16380 17490 16436 17500
rect 16156 17444 16212 17454
rect 16156 17350 16212 17388
rect 16604 17442 16660 17454
rect 16604 17390 16606 17442
rect 16658 17390 16660 17442
rect 16604 17220 16660 17390
rect 16604 17154 16660 17164
rect 16940 17444 16996 17454
rect 17052 17444 17108 18060
rect 17612 17668 17668 19068
rect 18172 18450 18228 19740
rect 18396 19122 18452 19134
rect 18396 19070 18398 19122
rect 18450 19070 18452 19122
rect 18396 18564 18452 19070
rect 18396 18498 18452 18508
rect 18172 18398 18174 18450
rect 18226 18398 18228 18450
rect 17724 18228 17780 18238
rect 17724 18134 17780 18172
rect 18172 18004 18228 18398
rect 18284 18450 18340 18462
rect 18284 18398 18286 18450
rect 18338 18398 18340 18450
rect 18284 18340 18340 18398
rect 18508 18452 18564 18462
rect 18508 18358 18564 18396
rect 18284 18274 18340 18284
rect 18620 18116 18676 22094
rect 19292 22146 19348 22158
rect 19292 22094 19294 22146
rect 19346 22094 19348 22146
rect 18844 21588 18900 21598
rect 19180 21588 19236 21598
rect 18844 21586 19236 21588
rect 18844 21534 18846 21586
rect 18898 21534 19182 21586
rect 19234 21534 19236 21586
rect 18844 21532 19236 21534
rect 18844 21476 18900 21532
rect 19180 21522 19236 21532
rect 18844 21410 18900 21420
rect 19068 18676 19124 18686
rect 19292 18676 19348 22094
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 19836 21914 20100 21924
rect 20076 20804 20132 20814
rect 20076 20710 20132 20748
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 19404 20132 19460 20142
rect 19404 20038 19460 20076
rect 19964 20020 20020 20030
rect 19964 19906 20020 19964
rect 19964 19854 19966 19906
rect 20018 19854 20020 19906
rect 19964 19842 20020 19854
rect 19628 19796 19684 19806
rect 19628 19702 19684 19740
rect 20188 18900 20244 22316
rect 20300 22306 20356 22316
rect 20860 22372 20916 22382
rect 20860 22278 20916 22316
rect 20524 22146 20580 22158
rect 20524 22094 20526 22146
rect 20578 22094 20580 22146
rect 20524 21812 20580 22094
rect 20748 22148 20804 22158
rect 20748 22146 20916 22148
rect 20748 22094 20750 22146
rect 20802 22094 20916 22146
rect 20748 22092 20916 22094
rect 20748 22082 20804 22092
rect 20412 20132 20468 20142
rect 20412 20038 20468 20076
rect 20300 20018 20356 20030
rect 20300 19966 20302 20018
rect 20354 19966 20356 20018
rect 20300 19796 20356 19966
rect 20300 19730 20356 19740
rect 20412 19124 20468 19134
rect 20524 19124 20580 21756
rect 20636 20132 20692 20142
rect 20636 20038 20692 20076
rect 20412 19122 20580 19124
rect 20412 19070 20414 19122
rect 20466 19070 20580 19122
rect 20412 19068 20580 19070
rect 20412 19058 20468 19068
rect 20748 19012 20804 19022
rect 20748 18918 20804 18956
rect 19836 18844 20100 18854
rect 20188 18844 20692 18900
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19124 18620 19348 18676
rect 20076 18674 20132 18686
rect 20076 18622 20078 18674
rect 20130 18622 20132 18674
rect 19068 18338 19124 18620
rect 20076 18564 20132 18622
rect 20076 18498 20132 18508
rect 19068 18286 19070 18338
rect 19122 18286 19124 18338
rect 19068 18274 19124 18286
rect 19404 18452 19460 18462
rect 18676 18060 18900 18116
rect 18620 18050 18676 18060
rect 17612 17602 17668 17612
rect 17724 17948 18228 18004
rect 16940 17442 17108 17444
rect 16940 17390 16942 17442
rect 16994 17390 17108 17442
rect 16940 17388 17108 17390
rect 17388 17554 17444 17566
rect 17388 17502 17390 17554
rect 17442 17502 17444 17554
rect 15932 16818 15988 16828
rect 15148 16718 15150 16770
rect 15202 16718 15204 16770
rect 15148 16706 15204 16718
rect 15596 16772 15652 16782
rect 15596 16678 15652 16716
rect 16268 16772 16324 16782
rect 14252 16146 14308 16156
rect 15596 16212 15652 16222
rect 15596 16118 15652 16156
rect 14700 16100 14756 16110
rect 14700 15426 14756 16044
rect 14700 15374 14702 15426
rect 14754 15374 14756 15426
rect 14700 15362 14756 15374
rect 16268 16098 16324 16716
rect 16268 16046 16270 16098
rect 16322 16046 16324 16098
rect 14028 15262 14030 15314
rect 14082 15262 14084 15314
rect 14028 15250 14084 15262
rect 16268 15204 16324 16046
rect 16940 16098 16996 17388
rect 17388 17220 17444 17502
rect 17724 17554 17780 17948
rect 18732 17892 18788 17902
rect 18620 17836 18732 17892
rect 18284 17668 18340 17678
rect 17724 17502 17726 17554
rect 17778 17502 17780 17554
rect 17724 17490 17780 17502
rect 18060 17554 18116 17566
rect 18060 17502 18062 17554
rect 18114 17502 18116 17554
rect 17388 17154 17444 17164
rect 17836 17444 17892 17454
rect 17836 17106 17892 17388
rect 17836 17054 17838 17106
rect 17890 17054 17892 17106
rect 17836 17042 17892 17054
rect 17948 17332 18004 17342
rect 17388 16884 17444 16894
rect 16940 16046 16942 16098
rect 16994 16046 16996 16098
rect 16940 16034 16996 16046
rect 17276 16882 17444 16884
rect 17276 16830 17390 16882
rect 17442 16830 17444 16882
rect 17276 16828 17444 16830
rect 17276 16098 17332 16828
rect 17388 16818 17444 16828
rect 17612 16884 17668 16894
rect 17276 16046 17278 16098
rect 17330 16046 17332 16098
rect 17276 16034 17332 16046
rect 17500 16770 17556 16782
rect 17500 16718 17502 16770
rect 17554 16718 17556 16770
rect 17500 16100 17556 16718
rect 17612 16660 17668 16828
rect 17948 16882 18004 17276
rect 18060 17220 18116 17502
rect 18284 17554 18340 17612
rect 18284 17502 18286 17554
rect 18338 17502 18340 17554
rect 18284 17490 18340 17502
rect 18620 17666 18676 17836
rect 18732 17826 18788 17836
rect 18620 17614 18622 17666
rect 18674 17614 18676 17666
rect 18060 17154 18116 17164
rect 18172 17442 18228 17454
rect 18172 17390 18174 17442
rect 18226 17390 18228 17442
rect 18172 16996 18228 17390
rect 18620 17332 18676 17614
rect 18732 17668 18788 17678
rect 18732 17332 18788 17612
rect 18844 17554 18900 18060
rect 18844 17502 18846 17554
rect 18898 17502 18900 17554
rect 18844 17490 18900 17502
rect 18956 17554 19012 17566
rect 18956 17502 18958 17554
rect 19010 17502 19012 17554
rect 18956 17444 19012 17502
rect 19404 17444 19460 18396
rect 19740 18452 19796 18462
rect 20524 18452 20580 18462
rect 19740 18450 19908 18452
rect 19740 18398 19742 18450
rect 19794 18398 19908 18450
rect 19740 18396 19908 18398
rect 19740 18386 19796 18396
rect 18956 17378 19012 17388
rect 19068 17442 19460 17444
rect 19068 17390 19406 17442
rect 19458 17390 19460 17442
rect 19068 17388 19460 17390
rect 18732 17276 18900 17332
rect 18620 17266 18676 17276
rect 18172 16930 18228 16940
rect 17948 16830 17950 16882
rect 18002 16830 18004 16882
rect 17948 16818 18004 16830
rect 18732 16884 18788 16894
rect 17612 16594 17668 16604
rect 17500 16034 17556 16044
rect 17052 15874 17108 15886
rect 17052 15822 17054 15874
rect 17106 15822 17108 15874
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 16268 14530 16324 15148
rect 16268 14478 16270 14530
rect 16322 14478 16324 14530
rect 16268 14466 16324 14478
rect 16828 15202 16884 15214
rect 16828 15150 16830 15202
rect 16882 15150 16884 15202
rect 16828 15148 16884 15150
rect 17052 15148 17108 15822
rect 17612 15874 17668 15886
rect 17612 15822 17614 15874
rect 17666 15822 17668 15874
rect 16828 15092 17108 15148
rect 17500 15204 17556 15242
rect 17612 15204 17668 15822
rect 17556 15148 17668 15204
rect 17500 15138 17556 15148
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 16828 8428 16884 15092
rect 16940 14644 16996 14654
rect 16940 14550 16996 14588
rect 18508 13636 18564 13646
rect 18732 13636 18788 16828
rect 18844 16770 18900 17276
rect 18844 16718 18846 16770
rect 18898 16718 18900 16770
rect 18844 16706 18900 16718
rect 19068 15986 19124 17388
rect 19404 17378 19460 17388
rect 19516 18340 19572 18350
rect 19068 15934 19070 15986
rect 19122 15934 19124 15986
rect 19068 15922 19124 15934
rect 19180 16882 19236 16894
rect 19180 16830 19182 16882
rect 19234 16830 19236 16882
rect 19180 16100 19236 16830
rect 19404 16884 19460 16894
rect 19516 16884 19572 18284
rect 19852 18004 19908 18396
rect 20636 18452 20692 18844
rect 20860 18674 20916 22092
rect 20860 18622 20862 18674
rect 20914 18622 20916 18674
rect 20748 18452 20804 18462
rect 20636 18396 20748 18452
rect 20524 18358 20580 18396
rect 20748 18386 20804 18396
rect 20860 18228 20916 18622
rect 20860 18162 20916 18172
rect 21084 18676 21140 25228
rect 21420 25218 21476 25228
rect 21868 25172 21924 25900
rect 22092 25508 22148 26796
rect 22428 26180 22484 37996
rect 24556 38050 24612 38062
rect 24556 37998 24558 38050
rect 24610 37998 24612 38050
rect 22652 27748 22708 27758
rect 22092 25414 22148 25452
rect 22316 26178 22484 26180
rect 22316 26126 22430 26178
rect 22482 26126 22484 26178
rect 22316 26124 22484 26126
rect 21980 25284 22036 25294
rect 22316 25284 22372 26124
rect 22428 26114 22484 26124
rect 22540 27692 22652 27748
rect 22428 25844 22484 25854
rect 22428 25730 22484 25788
rect 22428 25678 22430 25730
rect 22482 25678 22484 25730
rect 22428 25666 22484 25678
rect 22540 25618 22596 27692
rect 22652 27654 22708 27692
rect 23212 27746 23268 27758
rect 23212 27694 23214 27746
rect 23266 27694 23268 27746
rect 23212 27076 23268 27694
rect 24556 27748 24612 37998
rect 24892 37492 24948 41200
rect 25564 38276 25620 38286
rect 25564 38182 25620 38220
rect 26236 38276 26292 41200
rect 26236 38210 26292 38220
rect 27468 38276 27524 38286
rect 27468 38182 27524 38220
rect 34300 37940 34356 41200
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 34524 37940 34580 37950
rect 34300 37938 34580 37940
rect 34300 37886 34526 37938
rect 34578 37886 34580 37938
rect 34300 37884 34580 37886
rect 34524 37874 34580 37884
rect 24892 37426 24948 37436
rect 26236 37492 26292 37502
rect 26236 37398 26292 37436
rect 24556 27682 24612 27692
rect 25228 37266 25284 37278
rect 25228 37214 25230 37266
rect 25282 37214 25284 37266
rect 25228 27186 25284 37214
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 25228 27134 25230 27186
rect 25282 27134 25284 27186
rect 23268 27020 23604 27076
rect 23212 27010 23268 27020
rect 23100 26964 23156 26974
rect 22764 26962 23156 26964
rect 22764 26910 23102 26962
rect 23154 26910 23156 26962
rect 22764 26908 23156 26910
rect 22764 26514 22820 26908
rect 23100 26898 23156 26908
rect 22764 26462 22766 26514
rect 22818 26462 22820 26514
rect 22764 26450 22820 26462
rect 23548 26516 23604 27020
rect 23548 26422 23604 26460
rect 24108 26628 24164 26638
rect 24108 26514 24164 26572
rect 25228 26628 25284 27134
rect 25228 26562 25284 26572
rect 25676 26962 25732 26974
rect 25676 26910 25678 26962
rect 25730 26910 25732 26962
rect 24108 26462 24110 26514
rect 24162 26462 24164 26514
rect 24108 26450 24164 26462
rect 24556 26516 24612 26526
rect 22988 26404 23044 26414
rect 22988 26310 23044 26348
rect 23100 26292 23156 26302
rect 23100 26198 23156 26236
rect 23884 26292 23940 26302
rect 23884 26198 23940 26236
rect 24220 26290 24276 26302
rect 24220 26238 24222 26290
rect 24274 26238 24276 26290
rect 22540 25566 22542 25618
rect 22594 25566 22596 25618
rect 22540 25554 22596 25566
rect 21980 25282 22372 25284
rect 21980 25230 21982 25282
rect 22034 25230 22372 25282
rect 21980 25228 22372 25230
rect 23660 25508 23716 25518
rect 21980 25218 22036 25228
rect 21756 25116 21924 25172
rect 21756 24946 21812 25116
rect 21756 24894 21758 24946
rect 21810 24894 21812 24946
rect 21756 24882 21812 24894
rect 23660 24946 23716 25452
rect 24220 25508 24276 26238
rect 24220 25442 24276 25452
rect 24556 25506 24612 26460
rect 25676 26516 25732 26910
rect 40236 26852 40292 26862
rect 40236 26758 40292 26796
rect 25676 26450 25732 26460
rect 27916 26516 27972 26526
rect 27468 25620 27524 25630
rect 24556 25454 24558 25506
rect 24610 25454 24612 25506
rect 23660 24894 23662 24946
rect 23714 24894 23716 24946
rect 23660 24882 23716 24894
rect 21420 24836 21476 24846
rect 21420 24742 21476 24780
rect 21532 24834 21588 24846
rect 21532 24782 21534 24834
rect 21586 24782 21588 24834
rect 21196 23156 21252 23166
rect 21196 23062 21252 23100
rect 21532 22708 21588 24782
rect 23884 24722 23940 24734
rect 23884 24670 23886 24722
rect 23938 24670 23940 24722
rect 23884 23380 23940 24670
rect 23884 23314 23940 23324
rect 24220 23716 24276 23726
rect 24556 23716 24612 25454
rect 25116 25508 25172 25518
rect 25116 24724 25172 25452
rect 25340 25396 25396 25406
rect 25340 25394 25620 25396
rect 25340 25342 25342 25394
rect 25394 25342 25620 25394
rect 25340 25340 25620 25342
rect 25340 25330 25396 25340
rect 25564 24946 25620 25340
rect 25564 24894 25566 24946
rect 25618 24894 25620 24946
rect 25564 24882 25620 24894
rect 25676 24836 25732 24846
rect 25676 24742 25732 24780
rect 26460 24836 26516 24846
rect 26460 24742 26516 24780
rect 27468 24836 27524 25564
rect 27916 25618 27972 26460
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 27916 25566 27918 25618
rect 27970 25566 27972 25618
rect 27916 25554 27972 25566
rect 40012 25618 40068 25630
rect 40012 25566 40014 25618
rect 40066 25566 40068 25618
rect 37660 25508 37716 25518
rect 37660 25414 37716 25452
rect 40012 24948 40068 25566
rect 40012 24882 40068 24892
rect 27468 24770 27524 24780
rect 25228 24724 25284 24734
rect 25116 24722 25284 24724
rect 25116 24670 25230 24722
rect 25282 24670 25284 24722
rect 25116 24668 25284 24670
rect 25228 24658 25284 24668
rect 25340 24724 25396 24734
rect 24220 23714 24612 23716
rect 24220 23662 24222 23714
rect 24274 23662 24612 23714
rect 24220 23660 24612 23662
rect 25340 23716 25396 24668
rect 25452 24724 25508 24734
rect 25788 24724 25844 24734
rect 25452 24722 25620 24724
rect 25452 24670 25454 24722
rect 25506 24670 25620 24722
rect 25452 24668 25620 24670
rect 25452 24658 25508 24668
rect 25564 24500 25620 24668
rect 25788 24630 25844 24668
rect 26348 24500 26404 24510
rect 25564 24498 26404 24500
rect 25564 24446 26350 24498
rect 26402 24446 26404 24498
rect 25564 24444 26404 24446
rect 26348 24434 26404 24444
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 25340 23660 25620 23716
rect 23212 23268 23268 23278
rect 21868 23044 21924 23054
rect 22988 23044 23044 23054
rect 21868 23042 22036 23044
rect 21868 22990 21870 23042
rect 21922 22990 22036 23042
rect 21868 22988 22036 22990
rect 21868 22978 21924 22988
rect 21196 22652 21588 22708
rect 21196 18676 21252 22652
rect 21644 22484 21700 22494
rect 21644 22390 21700 22428
rect 21420 22372 21476 22382
rect 21476 22316 21588 22372
rect 21420 22306 21476 22316
rect 21308 22260 21364 22270
rect 21308 22166 21364 22204
rect 21532 22258 21588 22316
rect 21532 22206 21534 22258
rect 21586 22206 21588 22258
rect 21532 22194 21588 22206
rect 21756 22146 21812 22158
rect 21756 22094 21758 22146
rect 21810 22094 21812 22146
rect 21756 21140 21812 22094
rect 21308 21084 21812 21140
rect 21868 22148 21924 22158
rect 21308 19908 21364 21084
rect 21868 20916 21924 22092
rect 21308 19842 21364 19852
rect 21420 20860 21924 20916
rect 21980 20914 22036 22988
rect 22988 22370 23044 22988
rect 23212 22482 23268 23212
rect 24220 23156 24276 23660
rect 24332 23380 24388 23390
rect 24332 23266 24388 23324
rect 24332 23214 24334 23266
rect 24386 23214 24388 23266
rect 24332 23202 24388 23214
rect 24444 23268 24500 23278
rect 24444 23174 24500 23212
rect 23996 23044 24052 23054
rect 23996 22950 24052 22988
rect 23212 22430 23214 22482
rect 23266 22430 23268 22482
rect 23212 22418 23268 22430
rect 22988 22318 22990 22370
rect 23042 22318 23044 22370
rect 22988 22306 23044 22318
rect 24220 22372 24276 23100
rect 24220 22306 24276 22316
rect 24668 23154 24724 23166
rect 24668 23102 24670 23154
rect 24722 23102 24724 23154
rect 22316 22148 22372 22158
rect 22316 22054 22372 22092
rect 22428 22146 22484 22158
rect 22428 22094 22430 22146
rect 22482 22094 22484 22146
rect 21980 20862 21982 20914
rect 22034 20862 22036 20914
rect 21420 20802 21476 20860
rect 21980 20850 22036 20862
rect 22092 21700 22148 21710
rect 21420 20750 21422 20802
rect 21474 20750 21476 20802
rect 21420 20020 21476 20750
rect 21868 20692 21924 20702
rect 21532 20578 21588 20590
rect 21532 20526 21534 20578
rect 21586 20526 21588 20578
rect 21532 20132 21588 20526
rect 21756 20580 21812 20590
rect 21756 20486 21812 20524
rect 21532 20066 21588 20076
rect 21420 19346 21476 19964
rect 21420 19294 21422 19346
rect 21474 19294 21476 19346
rect 21420 19282 21476 19294
rect 21868 19572 21924 20636
rect 21980 20692 22036 20702
rect 22092 20692 22148 21644
rect 22428 20802 22484 22094
rect 22428 20750 22430 20802
rect 22482 20750 22484 20802
rect 22428 20738 22484 20750
rect 22540 22146 22596 22158
rect 22540 22094 22542 22146
rect 22594 22094 22596 22146
rect 21980 20690 22148 20692
rect 21980 20638 21982 20690
rect 22034 20638 22148 20690
rect 21980 20636 22148 20638
rect 21980 20626 22036 20636
rect 22204 20580 22260 20590
rect 21868 19236 21924 19516
rect 21644 19234 21924 19236
rect 21644 19182 21870 19234
rect 21922 19182 21924 19234
rect 21644 19180 21924 19182
rect 21532 19012 21588 19022
rect 21196 18620 21364 18676
rect 20188 18004 20244 18014
rect 19852 17948 20188 18004
rect 19740 17556 19796 17566
rect 19740 17462 19796 17500
rect 19628 17444 19684 17454
rect 19628 17108 19684 17388
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 19740 17108 19796 17118
rect 19628 17106 19796 17108
rect 19628 17054 19742 17106
rect 19794 17054 19796 17106
rect 19628 17052 19796 17054
rect 19740 17042 19796 17052
rect 19460 16828 19572 16884
rect 19404 16790 19460 16828
rect 20188 16770 20244 17948
rect 21084 17892 21140 18620
rect 21196 18450 21252 18462
rect 21196 18398 21198 18450
rect 21250 18398 21252 18450
rect 21196 18340 21252 18398
rect 21196 18274 21252 18284
rect 21084 17826 21140 17836
rect 20412 17556 20468 17566
rect 20412 17332 20468 17500
rect 20412 17106 20468 17276
rect 20412 17054 20414 17106
rect 20466 17054 20468 17106
rect 20412 17042 20468 17054
rect 20188 16718 20190 16770
rect 20242 16718 20244 16770
rect 20188 16706 20244 16718
rect 20524 16660 20580 16670
rect 20524 16658 20916 16660
rect 20524 16606 20526 16658
rect 20578 16606 20916 16658
rect 20524 16604 20916 16606
rect 20524 16594 20580 16604
rect 19292 16100 19348 16110
rect 19180 16098 19348 16100
rect 19180 16046 19294 16098
rect 19346 16046 19348 16098
rect 19180 16044 19348 16046
rect 19180 15428 19236 16044
rect 19292 16034 19348 16044
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 19852 15428 19908 15438
rect 19180 15426 19908 15428
rect 19180 15374 19854 15426
rect 19906 15374 19908 15426
rect 19180 15372 19908 15374
rect 19068 14644 19124 14654
rect 19180 14644 19236 15372
rect 19852 15362 19908 15372
rect 19964 15428 20020 15438
rect 19964 15334 20020 15372
rect 20860 15426 20916 16604
rect 21308 16324 21364 18620
rect 21532 18674 21588 18956
rect 21532 18622 21534 18674
rect 21586 18622 21588 18674
rect 21532 18610 21588 18622
rect 21644 18452 21700 19180
rect 21868 19170 21924 19180
rect 22092 20524 22204 20580
rect 21756 19012 21812 19022
rect 21756 19010 21924 19012
rect 21756 18958 21758 19010
rect 21810 18958 21924 19010
rect 21756 18956 21924 18958
rect 21756 18946 21812 18956
rect 20860 15374 20862 15426
rect 20914 15374 20916 15426
rect 20860 15362 20916 15374
rect 20972 16322 21364 16324
rect 20972 16270 21310 16322
rect 21362 16270 21364 16322
rect 20972 16268 21364 16270
rect 19068 14642 19236 14644
rect 19068 14590 19070 14642
rect 19122 14590 19236 14642
rect 19068 14588 19236 14590
rect 19516 15204 19572 15214
rect 19516 14642 19572 15148
rect 20636 15204 20692 15214
rect 20972 15204 21028 16268
rect 21308 16258 21364 16268
rect 21532 18396 21700 18452
rect 21308 16100 21364 16110
rect 21196 16098 21364 16100
rect 21196 16046 21310 16098
rect 21362 16046 21364 16098
rect 21196 16044 21364 16046
rect 21196 15428 21252 16044
rect 21308 16034 21364 16044
rect 21196 15334 21252 15372
rect 21532 15426 21588 18396
rect 21868 18116 21924 18956
rect 21980 18562 22036 18574
rect 21980 18510 21982 18562
rect 22034 18510 22036 18562
rect 21980 18452 22036 18510
rect 21980 18386 22036 18396
rect 21868 18050 21924 18060
rect 22092 17892 22148 20524
rect 22204 20486 22260 20524
rect 22540 20020 22596 22094
rect 24668 21812 24724 23102
rect 24668 21746 24724 21756
rect 25340 22258 25396 22270
rect 25340 22206 25342 22258
rect 25394 22206 25396 22258
rect 25340 21810 25396 22206
rect 25340 21758 25342 21810
rect 25394 21758 25396 21810
rect 25340 21746 25396 21758
rect 25228 21586 25284 21598
rect 25228 21534 25230 21586
rect 25282 21534 25284 21586
rect 23100 21474 23156 21486
rect 23100 21422 23102 21474
rect 23154 21422 23156 21474
rect 23100 20804 23156 21422
rect 23100 20710 23156 20748
rect 23100 20130 23156 20142
rect 23100 20078 23102 20130
rect 23154 20078 23156 20130
rect 22540 19954 22596 19964
rect 22764 20018 22820 20030
rect 22764 19966 22766 20018
rect 22818 19966 22820 20018
rect 22092 17826 22148 17836
rect 22204 19234 22260 19246
rect 22204 19182 22206 19234
rect 22258 19182 22260 19234
rect 22204 18676 22260 19182
rect 22652 18676 22708 18686
rect 22764 18676 22820 19966
rect 23100 20020 23156 20078
rect 23100 19954 23156 19964
rect 24444 20132 24500 20142
rect 24444 20018 24500 20076
rect 24444 19966 24446 20018
rect 24498 19966 24500 20018
rect 24444 19954 24500 19966
rect 24668 20130 24724 20142
rect 24668 20078 24670 20130
rect 24722 20078 24724 20130
rect 22988 19908 23044 19918
rect 22988 19236 23044 19852
rect 24668 19908 24724 20078
rect 23212 19460 23268 19470
rect 23212 19236 23268 19404
rect 22988 19180 23156 19236
rect 22204 18674 22820 18676
rect 22204 18622 22654 18674
rect 22706 18622 22820 18674
rect 22204 18620 22820 18622
rect 22876 19122 22932 19134
rect 22876 19070 22878 19122
rect 22930 19070 22932 19122
rect 21980 17668 22036 17678
rect 22204 17668 22260 18620
rect 22652 18610 22708 18620
rect 21644 17666 22260 17668
rect 21644 17614 21982 17666
rect 22034 17614 22260 17666
rect 21644 17612 22260 17614
rect 22316 18452 22372 18462
rect 22876 18452 22932 19070
rect 22316 18450 22932 18452
rect 22316 18398 22318 18450
rect 22370 18398 22932 18450
rect 22316 18396 22932 18398
rect 22988 19012 23044 19022
rect 23100 19012 23156 19180
rect 23212 19234 23604 19236
rect 23212 19182 23214 19234
rect 23266 19182 23604 19234
rect 23212 19180 23604 19182
rect 23212 19170 23268 19180
rect 23100 18956 23380 19012
rect 22988 18674 23044 18956
rect 22988 18622 22990 18674
rect 23042 18622 23044 18674
rect 22988 18452 23044 18622
rect 21644 16322 21700 17612
rect 21980 17602 22036 17612
rect 22316 17556 22372 18396
rect 22988 18386 23044 18396
rect 23100 18564 23156 18574
rect 22428 18116 22484 18126
rect 23100 18116 23156 18508
rect 22484 18060 22596 18116
rect 22428 18050 22484 18060
rect 22204 17500 22372 17556
rect 21756 17442 21812 17454
rect 21756 17390 21758 17442
rect 21810 17390 21812 17442
rect 21756 17332 21812 17390
rect 21756 17266 21812 17276
rect 21868 17442 21924 17454
rect 21868 17390 21870 17442
rect 21922 17390 21924 17442
rect 21868 17108 21924 17390
rect 21868 17052 22036 17108
rect 21756 16996 21812 17006
rect 21756 16902 21812 16940
rect 21980 16882 22036 17052
rect 22204 16996 22260 17500
rect 22204 16930 22260 16940
rect 21980 16830 21982 16882
rect 22034 16830 22036 16882
rect 21980 16818 22036 16830
rect 22316 16882 22372 16894
rect 22316 16830 22318 16882
rect 22370 16830 22372 16882
rect 21644 16270 21646 16322
rect 21698 16270 21700 16322
rect 21644 16258 21700 16270
rect 21868 16770 21924 16782
rect 21868 16718 21870 16770
rect 21922 16718 21924 16770
rect 21868 16324 21924 16718
rect 21868 16258 21924 16268
rect 21532 15374 21534 15426
rect 21586 15374 21588 15426
rect 20636 15202 21028 15204
rect 20636 15150 20638 15202
rect 20690 15150 21028 15202
rect 20636 15148 21028 15150
rect 20636 15138 20692 15148
rect 19516 14590 19518 14642
rect 19570 14590 19572 14642
rect 19068 14578 19124 14588
rect 19516 14578 19572 14590
rect 20300 15090 20356 15102
rect 20300 15038 20302 15090
rect 20354 15038 20356 15090
rect 20188 14532 20244 14542
rect 20300 14532 20356 15038
rect 21532 14644 21588 15374
rect 21532 14578 21588 14588
rect 21868 14644 21924 14654
rect 20188 14530 20356 14532
rect 20188 14478 20190 14530
rect 20242 14478 20356 14530
rect 20188 14476 20356 14478
rect 20188 14466 20244 14476
rect 20412 14308 20468 14318
rect 20412 14306 20692 14308
rect 20412 14254 20414 14306
rect 20466 14254 20692 14306
rect 20412 14252 20692 14254
rect 20412 14242 20468 14252
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 20636 13858 20692 14252
rect 20636 13806 20638 13858
rect 20690 13806 20692 13858
rect 20636 13794 20692 13806
rect 21420 13748 21476 13758
rect 21868 13748 21924 14588
rect 21420 13746 21924 13748
rect 21420 13694 21422 13746
rect 21474 13694 21870 13746
rect 21922 13694 21924 13746
rect 21420 13692 21924 13694
rect 21420 13682 21476 13692
rect 18508 13634 18788 13636
rect 18508 13582 18510 13634
rect 18562 13582 18788 13634
rect 18508 13580 18788 13582
rect 18508 13570 18564 13580
rect 21756 13074 21812 13692
rect 21868 13682 21924 13692
rect 22316 13636 22372 16830
rect 22540 16324 22596 18060
rect 22764 18060 23156 18116
rect 22652 17892 22708 17902
rect 22652 17798 22708 17836
rect 22764 17332 22820 18060
rect 22988 17780 23044 17790
rect 22988 17778 23268 17780
rect 22988 17726 22990 17778
rect 23042 17726 23268 17778
rect 22988 17724 23268 17726
rect 22988 17714 23044 17724
rect 22876 17554 22932 17566
rect 22876 17502 22878 17554
rect 22930 17502 22932 17554
rect 22876 17444 22932 17502
rect 22988 17444 23044 17454
rect 22876 17388 22988 17444
rect 22988 17378 23044 17388
rect 22764 17276 22932 17332
rect 22652 16884 22708 16894
rect 22708 16828 22820 16884
rect 22652 16790 22708 16828
rect 22764 16436 22820 16828
rect 22876 16882 22932 17276
rect 22876 16830 22878 16882
rect 22930 16830 22932 16882
rect 22876 16818 22932 16830
rect 23100 16770 23156 16782
rect 23100 16718 23102 16770
rect 23154 16718 23156 16770
rect 22876 16660 22932 16670
rect 23100 16660 23156 16718
rect 22932 16604 23156 16660
rect 23212 16660 23268 17724
rect 23324 17106 23380 18956
rect 23436 18676 23492 18686
rect 23436 18582 23492 18620
rect 23548 18562 23604 19180
rect 24668 18676 24724 19852
rect 25228 19460 25284 21534
rect 25452 21586 25508 21598
rect 25452 21534 25454 21586
rect 25506 21534 25508 21586
rect 25452 20916 25508 21534
rect 25228 19394 25284 19404
rect 25340 19794 25396 19806
rect 25340 19742 25342 19794
rect 25394 19742 25396 19794
rect 25004 19348 25060 19358
rect 25004 19254 25060 19292
rect 25340 19348 25396 19742
rect 25452 19796 25508 20860
rect 25564 20020 25620 23660
rect 37884 23268 37940 23278
rect 37660 23156 37716 23166
rect 37660 23062 37716 23100
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 26124 22372 26180 22382
rect 25676 21812 25732 21822
rect 25676 21718 25732 21756
rect 26124 21588 26180 22316
rect 37884 22370 37940 23212
rect 40012 22932 40068 22942
rect 40012 22838 40068 22876
rect 37884 22318 37886 22370
rect 37938 22318 37940 22370
rect 37884 22306 37940 22318
rect 40012 22482 40068 22494
rect 40012 22430 40014 22482
rect 40066 22430 40068 22482
rect 28140 22258 28196 22270
rect 28140 22206 28142 22258
rect 28194 22206 28196 22258
rect 26572 22146 26628 22158
rect 26572 22094 26574 22146
rect 26626 22094 26628 22146
rect 26236 21588 26292 21598
rect 26124 21586 26292 21588
rect 26124 21534 26238 21586
rect 26290 21534 26292 21586
rect 26124 21532 26292 21534
rect 25564 19926 25620 19964
rect 25900 20804 25956 20814
rect 25788 19906 25844 19918
rect 25788 19854 25790 19906
rect 25842 19854 25844 19906
rect 25452 19740 25620 19796
rect 25340 19282 25396 19292
rect 24668 18610 24724 18620
rect 23548 18510 23550 18562
rect 23602 18510 23604 18562
rect 23548 18498 23604 18510
rect 23660 18452 23716 18462
rect 23884 18452 23940 18462
rect 23716 18450 23940 18452
rect 23716 18398 23886 18450
rect 23938 18398 23940 18450
rect 23716 18396 23940 18398
rect 23660 18386 23716 18396
rect 23884 18386 23940 18396
rect 25228 18452 25284 18462
rect 25228 18358 25284 18396
rect 25452 18450 25508 18462
rect 25452 18398 25454 18450
rect 25506 18398 25508 18450
rect 24220 18340 24276 18350
rect 23436 18228 23492 18238
rect 23436 18226 23940 18228
rect 23436 18174 23438 18226
rect 23490 18174 23940 18226
rect 23436 18172 23940 18174
rect 23436 18162 23492 18172
rect 23548 17892 23604 17902
rect 23548 17666 23604 17836
rect 23548 17614 23550 17666
rect 23602 17614 23604 17666
rect 23548 17602 23604 17614
rect 23884 17666 23940 18172
rect 23996 18226 24052 18238
rect 23996 18174 23998 18226
rect 24050 18174 24052 18226
rect 23996 18004 24052 18174
rect 23996 17938 24052 17948
rect 24220 17890 24276 18284
rect 25340 18340 25396 18350
rect 25340 18246 25396 18284
rect 25452 18004 25508 18398
rect 25564 18228 25620 19740
rect 25788 19572 25844 19854
rect 25788 19506 25844 19516
rect 25900 19348 25956 20748
rect 26124 20692 26180 20702
rect 26236 20692 26292 21532
rect 26572 20692 26628 22094
rect 28028 22146 28084 22158
rect 28028 22094 28030 22146
rect 28082 22094 28084 22146
rect 26236 20690 26628 20692
rect 26236 20638 26574 20690
rect 26626 20638 26628 20690
rect 26236 20636 26628 20638
rect 26124 20242 26180 20636
rect 26124 20190 26126 20242
rect 26178 20190 26180 20242
rect 26124 20178 26180 20190
rect 26236 20468 26292 20478
rect 26012 20132 26068 20142
rect 26012 20038 26068 20076
rect 26236 20130 26292 20412
rect 26236 20078 26238 20130
rect 26290 20078 26292 20130
rect 26236 20066 26292 20078
rect 26572 20020 26628 20636
rect 26908 21474 26964 21486
rect 26908 21422 26910 21474
rect 26962 21422 26964 21474
rect 26908 20692 26964 21422
rect 26908 20626 26964 20636
rect 27468 20580 27524 20590
rect 27468 20130 27524 20524
rect 28028 20468 28084 22094
rect 28140 21476 28196 22206
rect 40012 22260 40068 22430
rect 40012 22194 40068 22204
rect 37660 21588 37716 21598
rect 37660 21494 37716 21532
rect 40012 21588 40068 21598
rect 28140 21410 28196 21420
rect 29036 21476 29092 21486
rect 29036 21382 29092 21420
rect 29484 21474 29540 21486
rect 29484 21422 29486 21474
rect 29538 21422 29540 21474
rect 29372 21364 29428 21374
rect 29260 21362 29428 21364
rect 29260 21310 29374 21362
rect 29426 21310 29428 21362
rect 29260 21308 29428 21310
rect 29260 20802 29316 21308
rect 29372 21298 29428 21308
rect 29484 21364 29540 21422
rect 29932 21476 29988 21486
rect 29932 21474 30100 21476
rect 29932 21422 29934 21474
rect 29986 21422 30100 21474
rect 29932 21420 30100 21422
rect 29932 21410 29988 21420
rect 29540 21308 29652 21364
rect 29484 21298 29540 21308
rect 29260 20750 29262 20802
rect 29314 20750 29316 20802
rect 29260 20738 29316 20750
rect 29372 20580 29428 20590
rect 29372 20486 29428 20524
rect 29484 20578 29540 20590
rect 29484 20526 29486 20578
rect 29538 20526 29540 20578
rect 28028 20402 28084 20412
rect 27468 20078 27470 20130
rect 27522 20078 27524 20130
rect 27468 20066 27524 20078
rect 26684 20020 26740 20030
rect 26572 20018 26740 20020
rect 26572 19966 26686 20018
rect 26738 19966 26740 20018
rect 26572 19964 26740 19966
rect 25956 19292 26292 19348
rect 25900 19254 25956 19292
rect 25564 18162 25620 18172
rect 25788 18450 25844 18462
rect 25788 18398 25790 18450
rect 25842 18398 25844 18450
rect 25452 17938 25508 17948
rect 24220 17838 24222 17890
rect 24274 17838 24276 17890
rect 24220 17826 24276 17838
rect 25788 17780 25844 18398
rect 26236 18450 26292 19292
rect 26236 18398 26238 18450
rect 26290 18398 26292 18450
rect 26236 18386 26292 18398
rect 26572 18452 26628 19964
rect 26684 19954 26740 19964
rect 26908 18676 26964 18686
rect 26908 18582 26964 18620
rect 29484 18676 29540 20526
rect 29596 19906 29652 21308
rect 29708 20916 29764 20926
rect 29708 20822 29764 20860
rect 29932 20802 29988 20814
rect 29932 20750 29934 20802
rect 29986 20750 29988 20802
rect 29932 20132 29988 20750
rect 29932 20066 29988 20076
rect 30044 20130 30100 21420
rect 40012 21474 40068 21532
rect 40012 21422 40014 21474
rect 40066 21422 40068 21474
rect 40012 21410 40068 21422
rect 37660 21364 37716 21374
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 30156 20804 30212 20814
rect 30604 20804 30660 20814
rect 30212 20802 30660 20804
rect 30212 20750 30606 20802
rect 30658 20750 30660 20802
rect 30212 20748 30660 20750
rect 30156 20710 30212 20748
rect 30604 20738 30660 20748
rect 37660 20802 37716 21308
rect 40012 20916 40068 20926
rect 40012 20822 40068 20860
rect 37660 20750 37662 20802
rect 37714 20750 37716 20802
rect 37660 20738 37716 20750
rect 30044 20078 30046 20130
rect 30098 20078 30100 20130
rect 29596 19854 29598 19906
rect 29650 19854 29652 19906
rect 29596 19842 29652 19854
rect 29484 18610 29540 18620
rect 26460 18226 26516 18238
rect 26460 18174 26462 18226
rect 26514 18174 26516 18226
rect 26460 18004 26516 18174
rect 26460 17938 26516 17948
rect 25788 17714 25844 17724
rect 23884 17614 23886 17666
rect 23938 17614 23940 17666
rect 23660 17556 23716 17566
rect 23660 17462 23716 17500
rect 23772 17444 23828 17454
rect 23772 17350 23828 17388
rect 23324 17054 23326 17106
rect 23378 17054 23380 17106
rect 23324 17042 23380 17054
rect 23548 16882 23604 16894
rect 23548 16830 23550 16882
rect 23602 16830 23604 16882
rect 23436 16770 23492 16782
rect 23436 16718 23438 16770
rect 23490 16718 23492 16770
rect 23212 16604 23380 16660
rect 22876 16594 22932 16604
rect 22764 16380 23044 16436
rect 22540 16268 22820 16324
rect 22764 16210 22820 16268
rect 22988 16322 23044 16380
rect 22988 16270 22990 16322
rect 23042 16270 23044 16322
rect 22988 16258 23044 16270
rect 23100 16324 23156 16334
rect 23156 16268 23268 16324
rect 23100 16258 23156 16268
rect 22764 16158 22766 16210
rect 22818 16158 22820 16210
rect 22764 16146 22820 16158
rect 23212 16210 23268 16268
rect 23324 16322 23380 16604
rect 23324 16270 23326 16322
rect 23378 16270 23380 16322
rect 23324 16258 23380 16270
rect 23212 16158 23214 16210
rect 23266 16158 23268 16210
rect 23212 16146 23268 16158
rect 22876 15874 22932 15886
rect 22876 15822 22878 15874
rect 22930 15822 22932 15874
rect 22764 15426 22820 15438
rect 22764 15374 22766 15426
rect 22818 15374 22820 15426
rect 22764 15148 22820 15374
rect 22876 15316 22932 15822
rect 22988 15316 23044 15326
rect 22876 15314 23044 15316
rect 22876 15262 22990 15314
rect 23042 15262 23044 15314
rect 22876 15260 23044 15262
rect 22988 15250 23044 15260
rect 22540 15092 22820 15148
rect 22540 13858 22596 15092
rect 22876 14644 22932 14654
rect 23436 14644 23492 16718
rect 23548 15540 23604 16830
rect 23884 16884 23940 17614
rect 23884 16818 23940 16828
rect 24668 17666 24724 17678
rect 24668 17614 24670 17666
rect 24722 17614 24724 17666
rect 24668 16884 24724 17614
rect 25340 17556 25396 17566
rect 25340 17462 25396 17500
rect 24668 16818 24724 16828
rect 26460 16884 26516 16894
rect 26572 16884 26628 18396
rect 27132 18452 27188 18462
rect 27916 18452 27972 18462
rect 30044 18452 30100 20078
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 27132 18450 27748 18452
rect 27132 18398 27134 18450
rect 27186 18398 27748 18450
rect 27132 18396 27748 18398
rect 27132 18386 27188 18396
rect 26684 18338 26740 18350
rect 26684 18286 26686 18338
rect 26738 18286 26740 18338
rect 26684 18228 26740 18286
rect 26684 18162 26740 18172
rect 27020 18338 27076 18350
rect 27020 18286 27022 18338
rect 27074 18286 27076 18338
rect 27020 16996 27076 18286
rect 27692 17890 27748 18396
rect 27692 17838 27694 17890
rect 27746 17838 27748 17890
rect 27692 17826 27748 17838
rect 27468 17780 27524 17790
rect 27468 17686 27524 17724
rect 27916 17778 27972 18396
rect 29820 18396 30044 18452
rect 28140 17892 28196 17902
rect 28364 17892 28420 17902
rect 28140 17890 28420 17892
rect 28140 17838 28142 17890
rect 28194 17838 28366 17890
rect 28418 17838 28420 17890
rect 28140 17836 28420 17838
rect 28140 17826 28196 17836
rect 28364 17826 28420 17836
rect 27916 17726 27918 17778
rect 27970 17726 27972 17778
rect 27916 17714 27972 17726
rect 28476 17668 28532 17678
rect 28476 17574 28532 17612
rect 29372 17668 29428 17678
rect 27244 16996 27300 17006
rect 27020 16994 27300 16996
rect 27020 16942 27246 16994
rect 27298 16942 27300 16994
rect 27020 16940 27300 16942
rect 27244 16930 27300 16940
rect 26516 16828 26628 16884
rect 23548 15474 23604 15484
rect 25228 15540 25284 15550
rect 25228 15446 25284 15484
rect 25340 15202 25396 15214
rect 25340 15150 25342 15202
rect 25394 15150 25396 15202
rect 25340 15148 25396 15150
rect 26460 15148 26516 16828
rect 29372 16770 29428 17612
rect 29820 17106 29876 18396
rect 30044 18386 30100 18396
rect 37660 18450 37716 18462
rect 37660 18398 37662 18450
rect 37714 18398 37716 18450
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 37660 17892 37716 18398
rect 40012 18228 40068 18238
rect 40012 18134 40068 18172
rect 37660 17826 37716 17836
rect 40012 17778 40068 17790
rect 40012 17726 40014 17778
rect 40066 17726 40068 17778
rect 37660 17668 37716 17678
rect 37660 17574 37716 17612
rect 40012 17556 40068 17726
rect 40012 17490 40068 17500
rect 29820 17054 29822 17106
rect 29874 17054 29876 17106
rect 29820 17042 29876 17054
rect 29372 16718 29374 16770
rect 29426 16718 29428 16770
rect 29372 16706 29428 16718
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 25340 15092 25508 15148
rect 23548 14644 23604 14654
rect 23436 14642 23604 14644
rect 23436 14590 23550 14642
rect 23602 14590 23604 14642
rect 23436 14588 23604 14590
rect 22876 14530 22932 14588
rect 23548 14578 23604 14588
rect 25340 14644 25396 14654
rect 25452 14644 25508 15092
rect 26124 15092 26516 15148
rect 25676 14644 25732 14654
rect 25452 14642 25732 14644
rect 25452 14590 25678 14642
rect 25730 14590 25732 14642
rect 25452 14588 25732 14590
rect 22876 14478 22878 14530
rect 22930 14478 22932 14530
rect 22876 14466 22932 14478
rect 25340 13970 25396 14588
rect 25340 13918 25342 13970
rect 25394 13918 25396 13970
rect 25340 13906 25396 13918
rect 22540 13806 22542 13858
rect 22594 13806 22596 13858
rect 22540 13794 22596 13806
rect 22316 13570 22372 13580
rect 24668 13636 24724 13646
rect 21756 13022 21758 13074
rect 21810 13022 21812 13074
rect 21756 13010 21812 13022
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 24668 8428 24724 13580
rect 25676 8428 25732 14588
rect 26124 14644 26180 15092
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 26124 14550 26180 14588
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 16828 8372 17108 8428
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 17052 3554 17108 8372
rect 24556 8372 24724 8428
rect 25228 8372 25732 8428
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 17052 3502 17054 3554
rect 17106 3502 17108 3554
rect 17052 3490 17108 3502
rect 23548 3668 23604 3678
rect 16828 3444 16884 3454
rect 16828 800 16884 3388
rect 18060 3444 18116 3454
rect 18060 3330 18116 3388
rect 18060 3278 18062 3330
rect 18114 3278 18116 3330
rect 18060 3266 18116 3278
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 23548 800 23604 3612
rect 24556 3554 24612 8372
rect 25228 4338 25284 8372
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 25228 4286 25230 4338
rect 25282 4286 25284 4338
rect 25228 4274 25284 4286
rect 24556 3502 24558 3554
rect 24610 3502 24612 3554
rect 24556 3490 24612 3502
rect 24892 4116 24948 4126
rect 24892 800 24948 4060
rect 26236 4116 26292 4126
rect 26236 4022 26292 4060
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 25564 3668 25620 3678
rect 25564 3574 25620 3612
rect 16800 0 16912 800
rect 23520 0 23632 800
rect 24864 0 24976 800
<< via2 >>
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 16828 37436 16884 37492
rect 16156 36652 16212 36708
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 1708 30268 1764 30324
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 4172 26908 4228 26964
rect 1932 24498 1988 24500
rect 1932 24446 1934 24498
rect 1934 24446 1986 24498
rect 1986 24446 1988 24498
rect 1932 24444 1988 24446
rect 1932 23548 1988 23604
rect 1932 22930 1988 22932
rect 1932 22878 1934 22930
rect 1934 22878 1986 22930
rect 1986 22878 1988 22930
rect 1932 22876 1988 22878
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 15596 26236 15652 26292
rect 14476 26178 14532 26180
rect 14476 26126 14478 26178
rect 14478 26126 14530 26178
rect 14530 26126 14532 26178
rect 14476 26124 14532 26126
rect 13804 25228 13860 25284
rect 15036 25228 15092 25284
rect 4284 24722 4340 24724
rect 4284 24670 4286 24722
rect 4286 24670 4338 24722
rect 4338 24670 4340 24722
rect 4284 24668 4340 24670
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 4284 23938 4340 23940
rect 4284 23886 4286 23938
rect 4286 23886 4338 23938
rect 4338 23886 4340 23938
rect 4284 23884 4340 23886
rect 11116 23884 11172 23940
rect 4284 23154 4340 23156
rect 4284 23102 4286 23154
rect 4286 23102 4338 23154
rect 4338 23102 4340 23154
rect 4284 23100 4340 23102
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 4172 21420 4228 21476
rect 11788 23100 11844 23156
rect 16268 26348 16324 26404
rect 15932 26124 15988 26180
rect 15708 25228 15764 25284
rect 16604 28082 16660 28084
rect 16604 28030 16606 28082
rect 16606 28030 16658 28082
rect 16658 28030 16660 28082
rect 16604 28028 16660 28030
rect 17388 36706 17444 36708
rect 17388 36654 17390 36706
rect 17390 36654 17442 36706
rect 17442 36654 17444 36706
rect 17388 36652 17444 36654
rect 17276 28028 17332 28084
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 18396 37490 18452 37492
rect 18396 37438 18398 37490
rect 18398 37438 18450 37490
rect 18450 37438 18452 37490
rect 18396 37436 18452 37438
rect 22876 38220 22932 38276
rect 21756 38050 21812 38052
rect 21756 37998 21758 38050
rect 21758 37998 21810 38050
rect 21810 37998 21812 38050
rect 21756 37996 21812 37998
rect 22428 37996 22484 38052
rect 20860 37436 20916 37492
rect 22092 37490 22148 37492
rect 22092 37438 22094 37490
rect 22094 37438 22146 37490
rect 22146 37438 22148 37490
rect 22092 37436 22148 37438
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 17612 27132 17668 27188
rect 16380 26124 16436 26180
rect 18508 27186 18564 27188
rect 18508 27134 18510 27186
rect 18510 27134 18562 27186
rect 18562 27134 18564 27186
rect 18508 27132 18564 27134
rect 20524 27746 20580 27748
rect 20524 27694 20526 27746
rect 20526 27694 20578 27746
rect 20578 27694 20580 27746
rect 20524 27692 20580 27694
rect 19628 27020 19684 27076
rect 17836 26402 17892 26404
rect 17836 26350 17838 26402
rect 17838 26350 17890 26402
rect 17890 26350 17892 26402
rect 17836 26348 17892 26350
rect 17388 26290 17444 26292
rect 17388 26238 17390 26290
rect 17390 26238 17442 26290
rect 17442 26238 17444 26290
rect 17388 26236 17444 26238
rect 18508 26178 18564 26180
rect 18508 26126 18510 26178
rect 18510 26126 18562 26178
rect 18562 26126 18564 26178
rect 18508 26124 18564 26126
rect 17164 25900 17220 25956
rect 11116 22316 11172 22372
rect 14588 23324 14644 23380
rect 14028 22594 14084 22596
rect 14028 22542 14030 22594
rect 14030 22542 14082 22594
rect 14082 22542 14084 22594
rect 14028 22540 14084 22542
rect 15036 23378 15092 23380
rect 15036 23326 15038 23378
rect 15038 23326 15090 23378
rect 15090 23326 15092 23378
rect 15036 23324 15092 23326
rect 14588 22540 14644 22596
rect 14700 22876 14756 22932
rect 13692 22370 13748 22372
rect 13692 22318 13694 22370
rect 13694 22318 13746 22370
rect 13746 22318 13748 22370
rect 13692 22316 13748 22318
rect 14476 22146 14532 22148
rect 14476 22094 14478 22146
rect 14478 22094 14530 22146
rect 14530 22094 14532 22146
rect 14476 22092 14532 22094
rect 15260 23154 15316 23156
rect 15260 23102 15262 23154
rect 15262 23102 15314 23154
rect 15314 23102 15316 23154
rect 15260 23100 15316 23102
rect 15148 23042 15204 23044
rect 15148 22990 15150 23042
rect 15150 22990 15202 23042
rect 15202 22990 15204 23042
rect 15148 22988 15204 22990
rect 15484 22092 15540 22148
rect 13580 21308 13636 21364
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 11228 20018 11284 20020
rect 11228 19966 11230 20018
rect 11230 19966 11282 20018
rect 11282 19966 11284 20018
rect 11228 19964 11284 19966
rect 11676 19964 11732 20020
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 12684 19740 12740 19796
rect 14140 19292 14196 19348
rect 14700 21308 14756 21364
rect 14476 20076 14532 20132
rect 14252 19964 14308 20020
rect 14700 19906 14756 19908
rect 14700 19854 14702 19906
rect 14702 19854 14754 19906
rect 14754 19854 14756 19906
rect 14700 19852 14756 19854
rect 15148 20130 15204 20132
rect 15148 20078 15150 20130
rect 15150 20078 15202 20130
rect 15202 20078 15204 20130
rect 15148 20076 15204 20078
rect 14364 19794 14420 19796
rect 14364 19742 14366 19794
rect 14366 19742 14418 19794
rect 14418 19742 14420 19794
rect 14364 19740 14420 19742
rect 14028 19068 14084 19124
rect 14924 19122 14980 19124
rect 14924 19070 14926 19122
rect 14926 19070 14978 19122
rect 14978 19070 14980 19122
rect 14924 19068 14980 19070
rect 13020 18508 13076 18564
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 4284 17666 4340 17668
rect 4284 17614 4286 17666
rect 4286 17614 4338 17666
rect 4338 17614 4340 17666
rect 4284 17612 4340 17614
rect 1932 16828 1988 16884
rect 14924 18284 14980 18340
rect 13468 17612 13524 17668
rect 12236 16716 12292 16772
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 14588 17612 14644 17668
rect 13916 17442 13972 17444
rect 13916 17390 13918 17442
rect 13918 17390 13970 17442
rect 13970 17390 13972 17442
rect 13916 17388 13972 17390
rect 14140 17276 14196 17332
rect 14028 16716 14084 16772
rect 14924 17388 14980 17444
rect 15148 19292 15204 19348
rect 15708 21756 15764 21812
rect 16828 25282 16884 25284
rect 16828 25230 16830 25282
rect 16830 25230 16882 25282
rect 16882 25230 16884 25282
rect 16828 25228 16884 25230
rect 16604 23660 16660 23716
rect 16828 23100 16884 23156
rect 16940 23324 16996 23380
rect 16380 22316 16436 22372
rect 16156 20076 16212 20132
rect 15260 19180 15316 19236
rect 15932 19740 15988 19796
rect 16604 20018 16660 20020
rect 16604 19966 16606 20018
rect 16606 19966 16658 20018
rect 16658 19966 16660 20018
rect 16604 19964 16660 19966
rect 15596 18620 15652 18676
rect 15708 18562 15764 18564
rect 15708 18510 15710 18562
rect 15710 18510 15762 18562
rect 15762 18510 15764 18562
rect 15708 18508 15764 18510
rect 15932 18284 15988 18340
rect 15260 17276 15316 17332
rect 15148 17164 15204 17220
rect 16156 18226 16212 18228
rect 16156 18174 16158 18226
rect 16158 18174 16210 18226
rect 16210 18174 16212 18226
rect 16156 18172 16212 18174
rect 16268 17948 16324 18004
rect 16044 17612 16100 17668
rect 18508 25900 18564 25956
rect 17836 24668 17892 24724
rect 17836 23548 17892 23604
rect 18060 23714 18116 23716
rect 18060 23662 18062 23714
rect 18062 23662 18114 23714
rect 18114 23662 18116 23714
rect 18060 23660 18116 23662
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 20300 24780 20356 24836
rect 18284 23548 18340 23604
rect 17948 23324 18004 23380
rect 17836 23154 17892 23156
rect 17836 23102 17838 23154
rect 17838 23102 17890 23154
rect 17890 23102 17892 23154
rect 17836 23100 17892 23102
rect 17276 22146 17332 22148
rect 17276 22094 17278 22146
rect 17278 22094 17330 22146
rect 17330 22094 17332 22146
rect 17276 22092 17332 22094
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 18396 23100 18452 23156
rect 18620 22428 18676 22484
rect 19852 22988 19908 23044
rect 18284 22316 18340 22372
rect 17948 22258 18004 22260
rect 17948 22206 17950 22258
rect 17950 22206 18002 22258
rect 18002 22206 18004 22258
rect 17948 22204 18004 22206
rect 19740 22370 19796 22372
rect 19740 22318 19742 22370
rect 19742 22318 19794 22370
rect 19794 22318 19796 22370
rect 19740 22316 19796 22318
rect 18396 22204 18452 22260
rect 17612 22092 17668 22148
rect 17836 21810 17892 21812
rect 17836 21758 17838 21810
rect 17838 21758 17890 21810
rect 17890 21758 17892 21810
rect 17836 21756 17892 21758
rect 18172 21756 18228 21812
rect 17724 20636 17780 20692
rect 18956 22258 19012 22260
rect 18956 22206 18958 22258
rect 18958 22206 19010 22258
rect 19010 22206 19012 22258
rect 18956 22204 19012 22206
rect 21644 27692 21700 27748
rect 22316 27074 22372 27076
rect 22316 27022 22318 27074
rect 22318 27022 22370 27074
rect 22370 27022 22372 27074
rect 22316 27020 22372 27022
rect 21308 25900 21364 25956
rect 21644 26348 21700 26404
rect 21756 26124 21812 26180
rect 20748 23042 20804 23044
rect 20748 22990 20750 23042
rect 20750 22990 20802 23042
rect 20802 22990 20804 23042
rect 20748 22988 20804 22990
rect 20076 22258 20132 22260
rect 20076 22206 20078 22258
rect 20078 22206 20130 22258
rect 20130 22206 20132 22258
rect 20076 22204 20132 22206
rect 17276 20188 17332 20244
rect 18060 20242 18116 20244
rect 18060 20190 18062 20242
rect 18062 20190 18114 20242
rect 18114 20190 18116 20242
rect 18060 20188 18116 20190
rect 17388 20130 17444 20132
rect 17388 20078 17390 20130
rect 17390 20078 17442 20130
rect 17442 20078 17444 20130
rect 17388 20076 17444 20078
rect 17276 19516 17332 19572
rect 18172 20130 18228 20132
rect 18172 20078 18174 20130
rect 18174 20078 18226 20130
rect 18226 20078 18228 20130
rect 18172 20076 18228 20078
rect 16940 19180 16996 19236
rect 16604 18060 16660 18116
rect 17276 18172 17332 18228
rect 18284 19964 18340 20020
rect 18172 19740 18228 19796
rect 18060 19516 18116 19572
rect 18060 19234 18116 19236
rect 18060 19182 18062 19234
rect 18062 19182 18114 19234
rect 18114 19182 18116 19234
rect 18060 19180 18116 19182
rect 17612 19068 17668 19124
rect 16940 17612 16996 17668
rect 17052 18060 17108 18116
rect 16380 17500 16436 17556
rect 16156 17442 16212 17444
rect 16156 17390 16158 17442
rect 16158 17390 16210 17442
rect 16210 17390 16212 17442
rect 16156 17388 16212 17390
rect 16604 17164 16660 17220
rect 18396 18508 18452 18564
rect 17724 18226 17780 18228
rect 17724 18174 17726 18226
rect 17726 18174 17778 18226
rect 17778 18174 17780 18226
rect 17724 18172 17780 18174
rect 18508 18450 18564 18452
rect 18508 18398 18510 18450
rect 18510 18398 18562 18450
rect 18562 18398 18564 18450
rect 18508 18396 18564 18398
rect 18284 18284 18340 18340
rect 18844 21420 18900 21476
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20044 21924 20100 21926
rect 20076 20802 20132 20804
rect 20076 20750 20078 20802
rect 20078 20750 20130 20802
rect 20130 20750 20132 20802
rect 20076 20748 20132 20750
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 19404 20130 19460 20132
rect 19404 20078 19406 20130
rect 19406 20078 19458 20130
rect 19458 20078 19460 20130
rect 19404 20076 19460 20078
rect 19964 19964 20020 20020
rect 19628 19794 19684 19796
rect 19628 19742 19630 19794
rect 19630 19742 19682 19794
rect 19682 19742 19684 19794
rect 19628 19740 19684 19742
rect 20860 22370 20916 22372
rect 20860 22318 20862 22370
rect 20862 22318 20914 22370
rect 20914 22318 20916 22370
rect 20860 22316 20916 22318
rect 20524 21756 20580 21812
rect 20412 20130 20468 20132
rect 20412 20078 20414 20130
rect 20414 20078 20466 20130
rect 20466 20078 20468 20130
rect 20412 20076 20468 20078
rect 20300 19740 20356 19796
rect 20636 20130 20692 20132
rect 20636 20078 20638 20130
rect 20638 20078 20690 20130
rect 20690 20078 20692 20130
rect 20636 20076 20692 20078
rect 20748 19010 20804 19012
rect 20748 18958 20750 19010
rect 20750 18958 20802 19010
rect 20802 18958 20804 19010
rect 20748 18956 20804 18958
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19068 18620 19124 18676
rect 20076 18508 20132 18564
rect 19404 18450 19460 18452
rect 19404 18398 19406 18450
rect 19406 18398 19458 18450
rect 19458 18398 19460 18450
rect 19404 18396 19460 18398
rect 18620 18060 18676 18116
rect 17612 17612 17668 17668
rect 15932 16828 15988 16884
rect 15596 16770 15652 16772
rect 15596 16718 15598 16770
rect 15598 16718 15650 16770
rect 15650 16718 15652 16770
rect 15596 16716 15652 16718
rect 16268 16716 16324 16772
rect 14252 16156 14308 16212
rect 15596 16210 15652 16212
rect 15596 16158 15598 16210
rect 15598 16158 15650 16210
rect 15650 16158 15652 16210
rect 15596 16156 15652 16158
rect 14700 16044 14756 16100
rect 18732 17836 18788 17892
rect 18284 17612 18340 17668
rect 17388 17164 17444 17220
rect 17836 17388 17892 17444
rect 17948 17276 18004 17332
rect 17612 16882 17668 16884
rect 17612 16830 17614 16882
rect 17614 16830 17666 16882
rect 17666 16830 17668 16882
rect 17612 16828 17668 16830
rect 18060 17164 18116 17220
rect 18620 17276 18676 17332
rect 18732 17612 18788 17668
rect 18956 17388 19012 17444
rect 18172 16940 18228 16996
rect 18732 16828 18788 16884
rect 17612 16604 17668 16660
rect 17500 16044 17556 16100
rect 16268 15148 16324 15204
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 17500 15202 17556 15204
rect 17500 15150 17502 15202
rect 17502 15150 17554 15202
rect 17554 15150 17556 15202
rect 17500 15148 17556 15150
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 16940 14642 16996 14644
rect 16940 14590 16942 14642
rect 16942 14590 16994 14642
rect 16994 14590 16996 14642
rect 16940 14588 16996 14590
rect 19516 18284 19572 18340
rect 20524 18450 20580 18452
rect 20524 18398 20526 18450
rect 20526 18398 20578 18450
rect 20578 18398 20580 18450
rect 20524 18396 20580 18398
rect 20748 18396 20804 18452
rect 20860 18172 20916 18228
rect 22092 25506 22148 25508
rect 22092 25454 22094 25506
rect 22094 25454 22146 25506
rect 22146 25454 22148 25506
rect 22092 25452 22148 25454
rect 22652 27746 22708 27748
rect 22652 27694 22654 27746
rect 22654 27694 22706 27746
rect 22706 27694 22708 27746
rect 22652 27692 22708 27694
rect 22428 25788 22484 25844
rect 25564 38274 25620 38276
rect 25564 38222 25566 38274
rect 25566 38222 25618 38274
rect 25618 38222 25620 38274
rect 25564 38220 25620 38222
rect 26236 38220 26292 38276
rect 27468 38274 27524 38276
rect 27468 38222 27470 38274
rect 27470 38222 27522 38274
rect 27522 38222 27524 38274
rect 27468 38220 27524 38222
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 24892 37436 24948 37492
rect 26236 37490 26292 37492
rect 26236 37438 26238 37490
rect 26238 37438 26290 37490
rect 26290 37438 26292 37490
rect 26236 37436 26292 37438
rect 24556 27692 24612 27748
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 23212 27020 23268 27076
rect 23548 26514 23604 26516
rect 23548 26462 23550 26514
rect 23550 26462 23602 26514
rect 23602 26462 23604 26514
rect 23548 26460 23604 26462
rect 24108 26572 24164 26628
rect 25228 26572 25284 26628
rect 24556 26460 24612 26516
rect 22988 26402 23044 26404
rect 22988 26350 22990 26402
rect 22990 26350 23042 26402
rect 23042 26350 23044 26402
rect 22988 26348 23044 26350
rect 23100 26290 23156 26292
rect 23100 26238 23102 26290
rect 23102 26238 23154 26290
rect 23154 26238 23156 26290
rect 23100 26236 23156 26238
rect 23884 26290 23940 26292
rect 23884 26238 23886 26290
rect 23886 26238 23938 26290
rect 23938 26238 23940 26290
rect 23884 26236 23940 26238
rect 23660 25452 23716 25508
rect 24220 25452 24276 25508
rect 40236 26850 40292 26852
rect 40236 26798 40238 26850
rect 40238 26798 40290 26850
rect 40290 26798 40292 26850
rect 40236 26796 40292 26798
rect 25676 26460 25732 26516
rect 27916 26460 27972 26516
rect 27468 25618 27524 25620
rect 27468 25566 27470 25618
rect 27470 25566 27522 25618
rect 27522 25566 27524 25618
rect 27468 25564 27524 25566
rect 21420 24834 21476 24836
rect 21420 24782 21422 24834
rect 21422 24782 21474 24834
rect 21474 24782 21476 24834
rect 21420 24780 21476 24782
rect 21196 23154 21252 23156
rect 21196 23102 21198 23154
rect 21198 23102 21250 23154
rect 21250 23102 21252 23154
rect 21196 23100 21252 23102
rect 23884 23324 23940 23380
rect 25116 25452 25172 25508
rect 25676 24834 25732 24836
rect 25676 24782 25678 24834
rect 25678 24782 25730 24834
rect 25730 24782 25732 24834
rect 25676 24780 25732 24782
rect 26460 24834 26516 24836
rect 26460 24782 26462 24834
rect 26462 24782 26514 24834
rect 26514 24782 26516 24834
rect 26460 24780 26516 24782
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 37660 25506 37716 25508
rect 37660 25454 37662 25506
rect 37662 25454 37714 25506
rect 37714 25454 37716 25506
rect 37660 25452 37716 25454
rect 40012 24892 40068 24948
rect 27468 24780 27524 24836
rect 25340 24668 25396 24724
rect 25788 24722 25844 24724
rect 25788 24670 25790 24722
rect 25790 24670 25842 24722
rect 25842 24670 25844 24722
rect 25788 24668 25844 24670
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 23212 23212 23268 23268
rect 21084 18620 21140 18676
rect 21644 22482 21700 22484
rect 21644 22430 21646 22482
rect 21646 22430 21698 22482
rect 21698 22430 21700 22482
rect 21644 22428 21700 22430
rect 21420 22316 21476 22372
rect 21308 22258 21364 22260
rect 21308 22206 21310 22258
rect 21310 22206 21362 22258
rect 21362 22206 21364 22258
rect 21308 22204 21364 22206
rect 21868 22146 21924 22148
rect 21868 22094 21870 22146
rect 21870 22094 21922 22146
rect 21922 22094 21924 22146
rect 21868 22092 21924 22094
rect 21308 19852 21364 19908
rect 22988 22988 23044 23044
rect 24332 23324 24388 23380
rect 24444 23266 24500 23268
rect 24444 23214 24446 23266
rect 24446 23214 24498 23266
rect 24498 23214 24500 23266
rect 24444 23212 24500 23214
rect 24220 23100 24276 23156
rect 23996 23042 24052 23044
rect 23996 22990 23998 23042
rect 23998 22990 24050 23042
rect 24050 22990 24052 23042
rect 23996 22988 24052 22990
rect 24220 22316 24276 22372
rect 22316 22146 22372 22148
rect 22316 22094 22318 22146
rect 22318 22094 22370 22146
rect 22370 22094 22372 22146
rect 22316 22092 22372 22094
rect 22092 21644 22148 21700
rect 21868 20636 21924 20692
rect 21756 20578 21812 20580
rect 21756 20526 21758 20578
rect 21758 20526 21810 20578
rect 21810 20526 21812 20578
rect 21756 20524 21812 20526
rect 21532 20076 21588 20132
rect 21420 19964 21476 20020
rect 21868 19516 21924 19572
rect 21532 18956 21588 19012
rect 20188 17948 20244 18004
rect 19740 17554 19796 17556
rect 19740 17502 19742 17554
rect 19742 17502 19794 17554
rect 19794 17502 19796 17554
rect 19740 17500 19796 17502
rect 19628 17388 19684 17444
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 19404 16882 19460 16884
rect 19404 16830 19406 16882
rect 19406 16830 19458 16882
rect 19458 16830 19460 16882
rect 19404 16828 19460 16830
rect 21196 18284 21252 18340
rect 21084 17836 21140 17892
rect 20412 17500 20468 17556
rect 20412 17276 20468 17332
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 19964 15426 20020 15428
rect 19964 15374 19966 15426
rect 19966 15374 20018 15426
rect 20018 15374 20020 15426
rect 19964 15372 20020 15374
rect 22204 20578 22260 20580
rect 22204 20526 22206 20578
rect 22206 20526 22258 20578
rect 22258 20526 22260 20578
rect 22204 20524 22260 20526
rect 19516 15148 19572 15204
rect 21196 15426 21252 15428
rect 21196 15374 21198 15426
rect 21198 15374 21250 15426
rect 21250 15374 21252 15426
rect 21196 15372 21252 15374
rect 21980 18396 22036 18452
rect 21868 18060 21924 18116
rect 24668 21756 24724 21812
rect 23100 20802 23156 20804
rect 23100 20750 23102 20802
rect 23102 20750 23154 20802
rect 23154 20750 23156 20802
rect 23100 20748 23156 20750
rect 22540 19964 22596 20020
rect 22092 17836 22148 17892
rect 23100 19964 23156 20020
rect 24444 20076 24500 20132
rect 22988 19852 23044 19908
rect 24668 19852 24724 19908
rect 23212 19404 23268 19460
rect 22988 19010 23044 19012
rect 22988 18958 22990 19010
rect 22990 18958 23042 19010
rect 23042 18958 23044 19010
rect 22988 18956 23044 18958
rect 22988 18396 23044 18452
rect 23100 18508 23156 18564
rect 22428 18060 22484 18116
rect 21756 17276 21812 17332
rect 21756 16994 21812 16996
rect 21756 16942 21758 16994
rect 21758 16942 21810 16994
rect 21810 16942 21812 16994
rect 21756 16940 21812 16942
rect 22204 16940 22260 16996
rect 21868 16268 21924 16324
rect 21532 14588 21588 14644
rect 21868 14588 21924 14644
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 22652 17890 22708 17892
rect 22652 17838 22654 17890
rect 22654 17838 22706 17890
rect 22706 17838 22708 17890
rect 22652 17836 22708 17838
rect 22988 17388 23044 17444
rect 22652 16882 22708 16884
rect 22652 16830 22654 16882
rect 22654 16830 22706 16882
rect 22706 16830 22708 16882
rect 22652 16828 22708 16830
rect 22876 16604 22932 16660
rect 23436 18674 23492 18676
rect 23436 18622 23438 18674
rect 23438 18622 23490 18674
rect 23490 18622 23492 18674
rect 23436 18620 23492 18622
rect 25452 20860 25508 20916
rect 25228 19404 25284 19460
rect 25004 19346 25060 19348
rect 25004 19294 25006 19346
rect 25006 19294 25058 19346
rect 25058 19294 25060 19346
rect 25004 19292 25060 19294
rect 37884 23212 37940 23268
rect 37660 23154 37716 23156
rect 37660 23102 37662 23154
rect 37662 23102 37714 23154
rect 37714 23102 37716 23154
rect 37660 23100 37716 23102
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 26124 22370 26180 22372
rect 26124 22318 26126 22370
rect 26126 22318 26178 22370
rect 26178 22318 26180 22370
rect 26124 22316 26180 22318
rect 25676 21810 25732 21812
rect 25676 21758 25678 21810
rect 25678 21758 25730 21810
rect 25730 21758 25732 21810
rect 25676 21756 25732 21758
rect 40012 22930 40068 22932
rect 40012 22878 40014 22930
rect 40014 22878 40066 22930
rect 40066 22878 40068 22930
rect 40012 22876 40068 22878
rect 25564 20018 25620 20020
rect 25564 19966 25566 20018
rect 25566 19966 25618 20018
rect 25618 19966 25620 20018
rect 25564 19964 25620 19966
rect 25900 20748 25956 20804
rect 25340 19292 25396 19348
rect 24668 18620 24724 18676
rect 23660 18396 23716 18452
rect 25228 18450 25284 18452
rect 25228 18398 25230 18450
rect 25230 18398 25282 18450
rect 25282 18398 25284 18450
rect 25228 18396 25284 18398
rect 24220 18284 24276 18340
rect 23548 17836 23604 17892
rect 23996 17948 24052 18004
rect 25340 18338 25396 18340
rect 25340 18286 25342 18338
rect 25342 18286 25394 18338
rect 25394 18286 25396 18338
rect 25340 18284 25396 18286
rect 25788 19516 25844 19572
rect 26124 20636 26180 20692
rect 26236 20412 26292 20468
rect 26012 20130 26068 20132
rect 26012 20078 26014 20130
rect 26014 20078 26066 20130
rect 26066 20078 26068 20130
rect 26012 20076 26068 20078
rect 26908 20636 26964 20692
rect 27468 20524 27524 20580
rect 40012 22204 40068 22260
rect 37660 21586 37716 21588
rect 37660 21534 37662 21586
rect 37662 21534 37714 21586
rect 37714 21534 37716 21586
rect 37660 21532 37716 21534
rect 40012 21532 40068 21588
rect 28140 21420 28196 21476
rect 29036 21474 29092 21476
rect 29036 21422 29038 21474
rect 29038 21422 29090 21474
rect 29090 21422 29092 21474
rect 29036 21420 29092 21422
rect 29484 21308 29540 21364
rect 29372 20578 29428 20580
rect 29372 20526 29374 20578
rect 29374 20526 29426 20578
rect 29426 20526 29428 20578
rect 29372 20524 29428 20526
rect 28028 20412 28084 20468
rect 25900 19346 25956 19348
rect 25900 19294 25902 19346
rect 25902 19294 25954 19346
rect 25954 19294 25956 19346
rect 25900 19292 25956 19294
rect 25564 18172 25620 18228
rect 25452 17948 25508 18004
rect 26908 18674 26964 18676
rect 26908 18622 26910 18674
rect 26910 18622 26962 18674
rect 26962 18622 26964 18674
rect 26908 18620 26964 18622
rect 29708 20914 29764 20916
rect 29708 20862 29710 20914
rect 29710 20862 29762 20914
rect 29762 20862 29764 20914
rect 29708 20860 29764 20862
rect 29932 20076 29988 20132
rect 37660 21308 37716 21364
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 30156 20802 30212 20804
rect 30156 20750 30158 20802
rect 30158 20750 30210 20802
rect 30210 20750 30212 20802
rect 30156 20748 30212 20750
rect 40012 20914 40068 20916
rect 40012 20862 40014 20914
rect 40014 20862 40066 20914
rect 40066 20862 40068 20914
rect 40012 20860 40068 20862
rect 29484 18620 29540 18676
rect 26572 18396 26628 18452
rect 26460 17948 26516 18004
rect 25788 17724 25844 17780
rect 23660 17554 23716 17556
rect 23660 17502 23662 17554
rect 23662 17502 23714 17554
rect 23714 17502 23716 17554
rect 23660 17500 23716 17502
rect 23772 17442 23828 17444
rect 23772 17390 23774 17442
rect 23774 17390 23826 17442
rect 23826 17390 23828 17442
rect 23772 17388 23828 17390
rect 23100 16268 23156 16324
rect 22876 14588 22932 14644
rect 23884 16828 23940 16884
rect 25340 17554 25396 17556
rect 25340 17502 25342 17554
rect 25342 17502 25394 17554
rect 25394 17502 25396 17554
rect 25340 17500 25396 17502
rect 24668 16828 24724 16884
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 26684 18172 26740 18228
rect 27916 18396 27972 18452
rect 27468 17778 27524 17780
rect 27468 17726 27470 17778
rect 27470 17726 27522 17778
rect 27522 17726 27524 17778
rect 27468 17724 27524 17726
rect 30044 18396 30100 18452
rect 28476 17666 28532 17668
rect 28476 17614 28478 17666
rect 28478 17614 28530 17666
rect 28530 17614 28532 17666
rect 28476 17612 28532 17614
rect 29372 17612 29428 17668
rect 26460 16882 26516 16884
rect 26460 16830 26462 16882
rect 26462 16830 26514 16882
rect 26514 16830 26516 16882
rect 26460 16828 26516 16830
rect 23548 15484 23604 15540
rect 25228 15538 25284 15540
rect 25228 15486 25230 15538
rect 25230 15486 25282 15538
rect 25282 15486 25284 15538
rect 25228 15484 25284 15486
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 40012 18226 40068 18228
rect 40012 18174 40014 18226
rect 40014 18174 40066 18226
rect 40066 18174 40068 18226
rect 40012 18172 40068 18174
rect 37660 17836 37716 17892
rect 37660 17666 37716 17668
rect 37660 17614 37662 17666
rect 37662 17614 37714 17666
rect 37714 17614 37716 17666
rect 37660 17612 37716 17614
rect 40012 17500 40068 17556
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 25340 14588 25396 14644
rect 22316 13580 22372 13636
rect 24668 13634 24724 13636
rect 24668 13582 24670 13634
rect 24670 13582 24722 13634
rect 24722 13582 24724 13634
rect 24668 13580 24724 13582
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 26124 14642 26180 14644
rect 26124 14590 26126 14642
rect 26126 14590 26178 14642
rect 26178 14590 26180 14642
rect 26124 14588 26180 14590
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 23548 3612 23604 3668
rect 16828 3388 16884 3444
rect 18060 3388 18116 3444
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 24892 4060 24948 4116
rect 26236 4114 26292 4116
rect 26236 4062 26238 4114
rect 26238 4062 26290 4114
rect 26290 4062 26292 4114
rect 26236 4060 26292 4062
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 25564 3666 25620 3668
rect 25564 3614 25566 3666
rect 25566 3614 25618 3666
rect 25618 3614 25620 3666
rect 25564 3612 25620 3614
<< metal3 >>
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 22866 38220 22876 38276
rect 22932 38220 25564 38276
rect 25620 38220 25630 38276
rect 26226 38220 26236 38276
rect 26292 38220 27468 38276
rect 27524 38220 27534 38276
rect 21746 37996 21756 38052
rect 21812 37996 22428 38052
rect 22484 37996 22494 38052
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 16818 37436 16828 37492
rect 16884 37436 18396 37492
rect 18452 37436 18462 37492
rect 20850 37436 20860 37492
rect 20916 37436 22092 37492
rect 22148 37436 22158 37492
rect 24882 37436 24892 37492
rect 24948 37436 26236 37492
rect 26292 37436 26302 37492
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 16146 36652 16156 36708
rect 16212 36652 17388 36708
rect 17444 36652 17454 36708
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 0 30324 800 30352
rect 0 30268 1708 30324
rect 1764 30268 1774 30324
rect 0 30240 800 30268
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 16594 28028 16604 28084
rect 16660 28028 17276 28084
rect 17332 28028 17342 28084
rect 20514 27692 20524 27748
rect 20580 27692 21644 27748
rect 21700 27692 21710 27748
rect 22642 27692 22652 27748
rect 22708 27692 24556 27748
rect 24612 27692 24622 27748
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 17602 27132 17612 27188
rect 17668 27132 18508 27188
rect 18564 27132 18574 27188
rect 19618 27020 19628 27076
rect 19684 27020 22316 27076
rect 22372 27020 23212 27076
rect 23268 27020 23278 27076
rect 0 26964 800 26992
rect 41200 26964 42000 26992
rect 0 26908 4172 26964
rect 4228 26908 4238 26964
rect 40236 26908 42000 26964
rect 0 26880 800 26908
rect 40236 26852 40292 26908
rect 41200 26880 42000 26908
rect 40226 26796 40236 26852
rect 40292 26796 40302 26852
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 24098 26572 24108 26628
rect 24164 26572 25228 26628
rect 25284 26572 25294 26628
rect 23538 26460 23548 26516
rect 23604 26460 24556 26516
rect 24612 26460 25676 26516
rect 25732 26460 27916 26516
rect 27972 26460 27982 26516
rect 16258 26348 16268 26404
rect 16324 26348 17836 26404
rect 17892 26348 17902 26404
rect 21634 26348 21644 26404
rect 21700 26348 22988 26404
rect 23044 26348 23054 26404
rect 15586 26236 15596 26292
rect 15652 26236 17388 26292
rect 17444 26236 17454 26292
rect 23090 26236 23100 26292
rect 23156 26236 23884 26292
rect 23940 26236 23950 26292
rect 14466 26124 14476 26180
rect 14532 26124 15932 26180
rect 15988 26124 15998 26180
rect 16370 26124 16380 26180
rect 16436 26124 18508 26180
rect 18564 26124 18574 26180
rect 21746 26124 21756 26180
rect 21812 26124 22484 26180
rect 17154 25900 17164 25956
rect 17220 25900 18508 25956
rect 18564 25900 21308 25956
rect 21364 25900 21374 25956
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 22428 25844 22484 26124
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 22418 25788 22428 25844
rect 22484 25788 22494 25844
rect 27458 25564 27468 25620
rect 27524 25564 31948 25620
rect 31892 25508 31948 25564
rect 22082 25452 22092 25508
rect 22148 25452 23660 25508
rect 23716 25452 24220 25508
rect 24276 25452 25116 25508
rect 25172 25452 25182 25508
rect 31892 25452 37660 25508
rect 37716 25452 37726 25508
rect 13794 25228 13804 25284
rect 13860 25228 15036 25284
rect 15092 25228 15708 25284
rect 15764 25228 16828 25284
rect 16884 25228 16894 25284
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 41200 24948 42000 24976
rect 40002 24892 40012 24948
rect 40068 24892 42000 24948
rect 41200 24864 42000 24892
rect 20290 24780 20300 24836
rect 20356 24780 21420 24836
rect 21476 24780 25676 24836
rect 25732 24780 25742 24836
rect 26450 24780 26460 24836
rect 26516 24780 27468 24836
rect 27524 24780 27534 24836
rect 4274 24668 4284 24724
rect 4340 24668 17836 24724
rect 17892 24668 17902 24724
rect 25330 24668 25340 24724
rect 25396 24668 25788 24724
rect 25844 24668 25854 24724
rect 1922 24444 1932 24500
rect 1988 24444 1998 24500
rect 0 24276 800 24304
rect 1932 24276 1988 24444
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 0 24220 1988 24276
rect 0 24192 800 24220
rect 4274 23884 4284 23940
rect 4340 23884 11116 23940
rect 11172 23884 11182 23940
rect 16594 23660 16604 23716
rect 16660 23660 18060 23716
rect 18116 23660 18126 23716
rect 0 23604 800 23632
rect 0 23548 1932 23604
rect 1988 23548 1998 23604
rect 17826 23548 17836 23604
rect 17892 23548 18284 23604
rect 18340 23548 18350 23604
rect 0 23520 800 23548
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 14578 23324 14588 23380
rect 14644 23324 15036 23380
rect 15092 23324 16940 23380
rect 16996 23324 17006 23380
rect 17938 23324 17948 23380
rect 18004 23324 23884 23380
rect 23940 23324 24332 23380
rect 24388 23324 24398 23380
rect 23202 23212 23212 23268
rect 23268 23212 24444 23268
rect 24500 23212 37884 23268
rect 37940 23212 37950 23268
rect 4274 23100 4284 23156
rect 4340 23100 11788 23156
rect 11844 23100 15260 23156
rect 15316 23100 15326 23156
rect 16818 23100 16828 23156
rect 16884 23100 17836 23156
rect 17892 23100 18396 23156
rect 18452 23100 18462 23156
rect 21186 23100 21196 23156
rect 21252 23100 24220 23156
rect 24276 23100 24286 23156
rect 31892 23100 37660 23156
rect 37716 23100 37726 23156
rect 31892 23044 31948 23100
rect 14700 22988 15148 23044
rect 15204 22988 15214 23044
rect 19842 22988 19852 23044
rect 19908 22988 20748 23044
rect 20804 22988 20814 23044
rect 22978 22988 22988 23044
rect 23044 22988 23996 23044
rect 24052 22988 31948 23044
rect 0 22932 800 22960
rect 14700 22932 14756 22988
rect 41200 22932 42000 22960
rect 0 22876 1932 22932
rect 1988 22876 1998 22932
rect 14690 22876 14700 22932
rect 14756 22876 14766 22932
rect 40002 22876 40012 22932
rect 40068 22876 42000 22932
rect 0 22848 800 22876
rect 41200 22848 42000 22876
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 14018 22540 14028 22596
rect 14084 22540 14588 22596
rect 14644 22540 14654 22596
rect 18610 22428 18620 22484
rect 18676 22428 21644 22484
rect 21700 22428 21710 22484
rect 11106 22316 11116 22372
rect 11172 22316 13692 22372
rect 13748 22316 13758 22372
rect 16370 22316 16380 22372
rect 16436 22316 18284 22372
rect 18340 22316 19740 22372
rect 19796 22316 19806 22372
rect 20850 22316 20860 22372
rect 20916 22316 21420 22372
rect 21476 22316 21486 22372
rect 24210 22316 24220 22372
rect 24276 22316 26124 22372
rect 26180 22316 26190 22372
rect 41200 22260 42000 22288
rect 17938 22204 17948 22260
rect 18004 22204 18396 22260
rect 18452 22204 18956 22260
rect 19012 22204 19022 22260
rect 20066 22204 20076 22260
rect 20132 22204 21308 22260
rect 21364 22204 21374 22260
rect 40002 22204 40012 22260
rect 40068 22204 42000 22260
rect 41200 22176 42000 22204
rect 14466 22092 14476 22148
rect 14532 22092 15484 22148
rect 15540 22092 15550 22148
rect 17266 22092 17276 22148
rect 17332 22092 17612 22148
rect 17668 22092 17678 22148
rect 21858 22092 21868 22148
rect 21924 22092 22316 22148
rect 22372 22092 22382 22148
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 15698 21756 15708 21812
rect 15764 21756 17836 21812
rect 17892 21756 18004 21812
rect 18162 21756 18172 21812
rect 18228 21756 20524 21812
rect 20580 21756 20590 21812
rect 24658 21756 24668 21812
rect 24724 21756 25676 21812
rect 25732 21756 25742 21812
rect 17948 21700 18004 21756
rect 17948 21644 22092 21700
rect 22148 21644 22158 21700
rect 41200 21588 42000 21616
rect 31892 21532 37660 21588
rect 37716 21532 37726 21588
rect 40002 21532 40012 21588
rect 40068 21532 42000 21588
rect 31892 21476 31948 21532
rect 41200 21504 42000 21532
rect 4162 21420 4172 21476
rect 4228 21420 18844 21476
rect 18900 21420 18910 21476
rect 28130 21420 28140 21476
rect 28196 21420 29036 21476
rect 29092 21420 31948 21476
rect 13570 21308 13580 21364
rect 13636 21308 14700 21364
rect 14756 21308 14766 21364
rect 29474 21308 29484 21364
rect 29540 21308 37660 21364
rect 37716 21308 37726 21364
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 41200 20916 42000 20944
rect 25442 20860 25452 20916
rect 25508 20860 29708 20916
rect 29764 20860 29774 20916
rect 40002 20860 40012 20916
rect 40068 20860 42000 20916
rect 41200 20832 42000 20860
rect 20066 20748 20076 20804
rect 20132 20748 23100 20804
rect 23156 20748 23166 20804
rect 25890 20748 25900 20804
rect 25956 20748 30156 20804
rect 30212 20748 30222 20804
rect 17714 20636 17724 20692
rect 17780 20636 21868 20692
rect 21924 20636 21934 20692
rect 26114 20636 26124 20692
rect 26180 20636 26908 20692
rect 26964 20636 26974 20692
rect 21746 20524 21756 20580
rect 21812 20524 22204 20580
rect 22260 20524 22270 20580
rect 27458 20524 27468 20580
rect 27524 20524 29372 20580
rect 29428 20524 29438 20580
rect 26226 20412 26236 20468
rect 26292 20412 28028 20468
rect 28084 20412 28094 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 17266 20188 17276 20244
rect 17332 20188 18060 20244
rect 18116 20188 18126 20244
rect 14466 20076 14476 20132
rect 14532 20076 15148 20132
rect 15204 20076 15214 20132
rect 16146 20076 16156 20132
rect 16212 20076 16222 20132
rect 17378 20076 17388 20132
rect 17444 20076 18172 20132
rect 18228 20076 19404 20132
rect 19460 20076 20412 20132
rect 20468 20076 20478 20132
rect 20626 20076 20636 20132
rect 20692 20076 21532 20132
rect 21588 20076 24444 20132
rect 24500 20076 26012 20132
rect 26068 20076 26078 20132
rect 26852 20076 29932 20132
rect 29988 20076 29998 20132
rect 11218 19964 11228 20020
rect 11284 19964 11676 20020
rect 11732 19964 14252 20020
rect 14308 19964 14318 20020
rect 16156 19908 16212 20076
rect 26852 20020 26908 20076
rect 16594 19964 16604 20020
rect 16660 19964 18284 20020
rect 18340 19964 18350 20020
rect 19954 19964 19964 20020
rect 20020 19964 21420 20020
rect 21476 19964 21486 20020
rect 22530 19964 22540 20020
rect 22596 19964 23100 20020
rect 23156 19964 25564 20020
rect 25620 19964 26908 20020
rect 14690 19852 14700 19908
rect 14756 19852 16212 19908
rect 16604 19796 16660 19964
rect 21298 19852 21308 19908
rect 21364 19852 22988 19908
rect 23044 19852 24668 19908
rect 24724 19852 24734 19908
rect 12674 19740 12684 19796
rect 12740 19740 14364 19796
rect 14420 19740 14430 19796
rect 15922 19740 15932 19796
rect 15988 19740 16660 19796
rect 18162 19740 18172 19796
rect 18228 19740 19628 19796
rect 19684 19740 20300 19796
rect 20356 19740 20366 19796
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 17266 19516 17276 19572
rect 17332 19516 18060 19572
rect 18116 19516 18126 19572
rect 21858 19516 21868 19572
rect 21924 19516 25788 19572
rect 25844 19516 25854 19572
rect 23202 19404 23212 19460
rect 23268 19404 25228 19460
rect 25284 19404 25294 19460
rect 14130 19292 14140 19348
rect 14196 19292 15148 19348
rect 15204 19292 25004 19348
rect 25060 19292 25340 19348
rect 25396 19292 25900 19348
rect 25956 19292 25966 19348
rect 15250 19180 15260 19236
rect 15316 19180 16940 19236
rect 16996 19180 18060 19236
rect 18116 19180 18126 19236
rect 14018 19068 14028 19124
rect 14084 19068 14924 19124
rect 14980 19068 17612 19124
rect 17668 19068 17678 19124
rect 20738 18956 20748 19012
rect 20804 18956 21532 19012
rect 21588 18956 22988 19012
rect 23044 18956 23054 19012
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 15586 18620 15596 18676
rect 15652 18620 19068 18676
rect 19124 18620 19134 18676
rect 21074 18620 21084 18676
rect 21140 18620 23436 18676
rect 23492 18620 23502 18676
rect 24658 18620 24668 18676
rect 24724 18620 26908 18676
rect 26964 18620 29484 18676
rect 29540 18620 29550 18676
rect 13010 18508 13020 18564
rect 13076 18508 15708 18564
rect 15764 18508 15774 18564
rect 18386 18508 18396 18564
rect 18452 18508 20076 18564
rect 20132 18508 23100 18564
rect 23156 18508 23166 18564
rect 18498 18396 18508 18452
rect 18564 18396 19404 18452
rect 19460 18396 20524 18452
rect 20580 18396 20590 18452
rect 20738 18396 20748 18452
rect 20804 18396 21980 18452
rect 22036 18396 22046 18452
rect 22978 18396 22988 18452
rect 23044 18396 23660 18452
rect 23716 18396 23726 18452
rect 23996 18396 25228 18452
rect 25284 18396 25294 18452
rect 26562 18396 26572 18452
rect 26628 18396 27916 18452
rect 27972 18396 30044 18452
rect 30100 18396 30110 18452
rect 21980 18340 22036 18396
rect 23996 18340 24052 18396
rect 14914 18284 14924 18340
rect 14980 18284 15932 18340
rect 15988 18284 15998 18340
rect 18274 18284 18284 18340
rect 18340 18284 19516 18340
rect 19572 18284 21196 18340
rect 21252 18284 21262 18340
rect 21980 18284 24052 18340
rect 24210 18284 24220 18340
rect 24276 18284 25340 18340
rect 25396 18284 25406 18340
rect 41200 18228 42000 18256
rect 16146 18172 16156 18228
rect 16212 18172 17276 18228
rect 17332 18172 17724 18228
rect 17780 18172 17790 18228
rect 20850 18172 20860 18228
rect 20916 18172 25564 18228
rect 25620 18172 26684 18228
rect 26740 18172 26750 18228
rect 40002 18172 40012 18228
rect 40068 18172 42000 18228
rect 41200 18144 42000 18172
rect 16594 18060 16604 18116
rect 16660 18060 17052 18116
rect 17108 18060 18620 18116
rect 18676 18060 18686 18116
rect 18844 18060 21868 18116
rect 21924 18060 22428 18116
rect 22484 18060 22494 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 18844 18004 18900 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 16258 17948 16268 18004
rect 16324 17948 18900 18004
rect 20178 17948 20188 18004
rect 20244 17948 23996 18004
rect 24052 17948 25452 18004
rect 25508 17948 26460 18004
rect 26516 17948 26526 18004
rect 18722 17836 18732 17892
rect 18788 17836 21084 17892
rect 21140 17836 21150 17892
rect 22082 17836 22092 17892
rect 22148 17836 22652 17892
rect 22708 17836 23548 17892
rect 23604 17836 23614 17892
rect 31892 17836 37660 17892
rect 37716 17836 37726 17892
rect 31892 17780 31948 17836
rect 25778 17724 25788 17780
rect 25844 17724 27468 17780
rect 27524 17724 31948 17780
rect 4274 17612 4284 17668
rect 4340 17612 13468 17668
rect 13524 17612 14588 17668
rect 14644 17612 14654 17668
rect 15092 17612 16044 17668
rect 16100 17612 16940 17668
rect 16996 17612 17006 17668
rect 17602 17612 17612 17668
rect 17668 17612 18284 17668
rect 18340 17612 18732 17668
rect 18788 17612 18798 17668
rect 28466 17612 28476 17668
rect 28532 17612 29372 17668
rect 29428 17612 37660 17668
rect 37716 17612 37726 17668
rect 15092 17444 15148 17612
rect 41200 17556 42000 17584
rect 16370 17500 16380 17556
rect 16436 17500 19740 17556
rect 19796 17500 20412 17556
rect 20468 17500 20478 17556
rect 23650 17500 23660 17556
rect 23716 17500 25340 17556
rect 25396 17500 25406 17556
rect 40002 17500 40012 17556
rect 40068 17500 42000 17556
rect 41200 17472 42000 17500
rect 13906 17388 13916 17444
rect 13972 17388 14924 17444
rect 14980 17388 15148 17444
rect 16146 17388 16156 17444
rect 16212 17388 17836 17444
rect 17892 17388 17902 17444
rect 18946 17388 18956 17444
rect 19012 17388 19628 17444
rect 19684 17388 22988 17444
rect 23044 17388 23772 17444
rect 23828 17388 23838 17444
rect 14130 17276 14140 17332
rect 14196 17276 15260 17332
rect 15316 17276 15326 17332
rect 17938 17276 17948 17332
rect 18004 17276 18620 17332
rect 18676 17276 18686 17332
rect 20402 17276 20412 17332
rect 20468 17276 21756 17332
rect 21812 17276 21822 17332
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 15138 17164 15148 17220
rect 15204 17164 16604 17220
rect 16660 17164 17388 17220
rect 17444 17164 18060 17220
rect 18116 17164 18126 17220
rect 18162 16940 18172 16996
rect 18228 16940 21756 16996
rect 21812 16940 22204 16996
rect 22260 16940 22270 16996
rect 0 16884 800 16912
rect 0 16828 1932 16884
rect 1988 16828 1998 16884
rect 15922 16828 15932 16884
rect 15988 16828 17612 16884
rect 17668 16828 17678 16884
rect 18722 16828 18732 16884
rect 18788 16828 19404 16884
rect 19460 16828 19470 16884
rect 22642 16828 22652 16884
rect 22708 16828 23884 16884
rect 23940 16828 23950 16884
rect 24658 16828 24668 16884
rect 24724 16828 26460 16884
rect 26516 16828 26526 16884
rect 0 16800 800 16828
rect 12226 16716 12236 16772
rect 12292 16716 14028 16772
rect 14084 16716 15596 16772
rect 15652 16716 16268 16772
rect 16324 16716 16334 16772
rect 17602 16604 17612 16660
rect 17668 16604 22876 16660
rect 22932 16604 22942 16660
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 21858 16268 21868 16324
rect 21924 16268 23100 16324
rect 23156 16268 23166 16324
rect 14242 16156 14252 16212
rect 14308 16156 15596 16212
rect 15652 16156 15662 16212
rect 14690 16044 14700 16100
rect 14756 16044 17500 16100
rect 17556 16044 17566 16100
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 23538 15484 23548 15540
rect 23604 15484 25228 15540
rect 25284 15484 25294 15540
rect 19954 15372 19964 15428
rect 20020 15372 21196 15428
rect 21252 15372 21262 15428
rect 16258 15148 16268 15204
rect 16324 15148 17500 15204
rect 17556 15148 19516 15204
rect 19572 15148 19582 15204
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 16930 14588 16940 14644
rect 16996 14588 21532 14644
rect 21588 14588 21598 14644
rect 21858 14588 21868 14644
rect 21924 14588 22876 14644
rect 22932 14588 25340 14644
rect 25396 14588 26124 14644
rect 26180 14588 26190 14644
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 22306 13580 22316 13636
rect 22372 13580 24668 13636
rect 24724 13580 24734 13636
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 24882 4060 24892 4116
rect 24948 4060 26236 4116
rect 26292 4060 26302 4116
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 23538 3612 23548 3668
rect 23604 3612 25564 3668
rect 25620 3612 25630 3668
rect 16818 3388 16828 3444
rect 16884 3388 18060 3444
rect 18116 3388 18126 3444
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
<< via3 >>
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 38444 4768 38476
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 37660 20128 38476
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 19808 17276 20128 18788
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 38444 35488 38476
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _096_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18368 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _097_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 17472 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _098_
timestamp 1698175906
transform 1 0 16464 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _099_
timestamp 1698175906
transform -1 0 18816 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _100_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _101_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18144 0 -1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _102_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 15680 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__and3_1  _103_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18704 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _104_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 17696 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _105_
timestamp 1698175906
transform -1 0 15232 0 -1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _106_
timestamp 1698175906
transform -1 0 14224 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _107_
timestamp 1698175906
transform -1 0 14000 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _108_
timestamp 1698175906
transform 1 0 19712 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _109_
timestamp 1698175906
transform 1 0 21056 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _110_
timestamp 1698175906
transform -1 0 20944 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _111_
timestamp 1698175906
transform -1 0 18144 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _112_
timestamp 1698175906
transform 1 0 14896 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _113_
timestamp 1698175906
transform -1 0 14896 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _114_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18368 0 -1 17248
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _115_
timestamp 1698175906
transform -1 0 19152 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _116_
timestamp 1698175906
transform -1 0 18144 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _117_
timestamp 1698175906
transform -1 0 24192 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _118_
timestamp 1698175906
transform -1 0 22288 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _119_
timestamp 1698175906
transform -1 0 21728 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _120_
timestamp 1698175906
transform 1 0 19264 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _121_
timestamp 1698175906
transform 1 0 20048 0 -1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _122_
timestamp 1698175906
transform -1 0 23184 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _123_
timestamp 1698175906
transform -1 0 21840 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _124_
timestamp 1698175906
transform -1 0 21056 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _125_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19936 0 1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _126_
timestamp 1698175906
transform -1 0 15456 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _127_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15904 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _128_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15456 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _129_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 17024 0 -1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _130_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 15120 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _131_
timestamp 1698175906
transform -1 0 12880 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _132_
timestamp 1698175906
transform 1 0 20160 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _133_
timestamp 1698175906
transform 1 0 24192 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _134_
timestamp 1698175906
transform 1 0 19264 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _135_
timestamp 1698175906
transform 1 0 20384 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _136_
timestamp 1698175906
transform 1 0 17920 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _137_
timestamp 1698175906
transform -1 0 22512 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _138_
timestamp 1698175906
transform 1 0 20160 0 1 21952
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _139_
timestamp 1698175906
transform 1 0 19600 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _140_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21168 0 1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _141_
timestamp 1698175906
transform 1 0 22624 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _142_
timestamp 1698175906
transform -1 0 14672 0 1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _143_
timestamp 1698175906
transform -1 0 29680 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _144_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 30352 0 1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _145_
timestamp 1698175906
transform 1 0 22736 0 1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _146_
timestamp 1698175906
transform 1 0 24192 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _147_
timestamp 1698175906
transform 1 0 25088 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _148_
timestamp 1698175906
transform 1 0 21280 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _149_
timestamp 1698175906
transform -1 0 24416 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _150_
timestamp 1698175906
transform -1 0 23296 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _151_
timestamp 1698175906
transform -1 0 22736 0 1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _152_
timestamp 1698175906
transform -1 0 23744 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _153_
timestamp 1698175906
transform -1 0 22176 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _154_
timestamp 1698175906
transform 1 0 21616 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _155_
timestamp 1698175906
transform 1 0 21280 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _156_
timestamp 1698175906
transform 1 0 22512 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _157_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 23632 0 1 15680
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _158_
timestamp 1698175906
transform -1 0 23296 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _159_
timestamp 1698175906
transform 1 0 25088 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _160_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 24416 0 1 17248
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _161_
timestamp 1698175906
transform -1 0 26656 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _162_
timestamp 1698175906
transform -1 0 26096 0 -1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _163_
timestamp 1698175906
transform 1 0 22176 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _164_
timestamp 1698175906
transform -1 0 22624 0 1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _165_
timestamp 1698175906
transform -1 0 28672 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _166_
timestamp 1698175906
transform 1 0 26096 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _167_
timestamp 1698175906
transform -1 0 18592 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _168_
timestamp 1698175906
transform 1 0 16016 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _169_
timestamp 1698175906
transform -1 0 16128 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _170_
timestamp 1698175906
transform -1 0 16352 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _171_
timestamp 1698175906
transform -1 0 25536 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _172_
timestamp 1698175906
transform 1 0 22512 0 -1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _173_
timestamp 1698175906
transform 1 0 16800 0 1 15680
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _174_
timestamp 1698175906
transform -1 0 16464 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _175_
timestamp 1698175906
transform -1 0 18256 0 -1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _176_
timestamp 1698175906
transform -1 0 14896 0 1 17248
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _177_
timestamp 1698175906
transform 1 0 13552 0 1 17248
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _178_
timestamp 1698175906
transform -1 0 22736 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _179_
timestamp 1698175906
transform 1 0 21168 0 1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _180_
timestamp 1698175906
transform -1 0 28336 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _181_
timestamp 1698175906
transform 1 0 25200 0 -1 20384
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _182_
timestamp 1698175906
transform 1 0 14784 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _183_
timestamp 1698175906
transform -1 0 19600 0 1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _184_
timestamp 1698175906
transform 1 0 21056 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _185_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 23744 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _186_
timestamp 1698175906
transform 1 0 17248 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _187_
timestamp 1698175906
transform -1 0 18592 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _188_
timestamp 1698175906
transform 1 0 18816 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _189_
timestamp 1698175906
transform 1 0 18704 0 -1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _190_
timestamp 1698175906
transform -1 0 18592 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _191_
timestamp 1698175906
transform -1 0 17920 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _192_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15456 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _193_
timestamp 1698175906
transform -1 0 14224 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _194_
timestamp 1698175906
transform -1 0 14896 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _195_
timestamp 1698175906
transform 1 0 19376 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _196_
timestamp 1698175906
transform 1 0 16016 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _197_
timestamp 1698175906
transform -1 0 21616 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _198_
timestamp 1698175906
transform 1 0 12096 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _199_
timestamp 1698175906
transform 1 0 10976 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _200_
timestamp 1698175906
transform 1 0 17696 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _201_
timestamp 1698175906
transform 1 0 26544 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _202_
timestamp 1698175906
transform -1 0 26320 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _203_
timestamp 1698175906
transform 1 0 22176 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _204_
timestamp 1698175906
transform 1 0 21616 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _205_
timestamp 1698175906
transform 1 0 24416 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _206_
timestamp 1698175906
transform 1 0 24416 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _207_
timestamp 1698175906
transform 1 0 20944 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _208_
timestamp 1698175906
transform 1 0 26320 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _209_
timestamp 1698175906
transform 1 0 14784 0 1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _210_
timestamp 1698175906
transform 1 0 13552 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _211_
timestamp 1698175906
transform 1 0 22624 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _212_
timestamp 1698175906
transform 1 0 13776 0 -1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _213_
timestamp 1698175906
transform -1 0 16576 0 1 15680
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _214_
timestamp 1698175906
transform 1 0 19600 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _215_
timestamp 1698175906
transform 1 0 25984 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _221_
timestamp 1698175906
transform 1 0 16128 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__144__A3 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 30576 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__166__A3
timestamp 1698175906
transform 1 0 25872 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__177__A1
timestamp 1698175906
transform 1 0 15120 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__181__A3
timestamp 1698175906
transform 1 0 24976 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__192__CLK
timestamp 1698175906
transform 1 0 18928 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__193__CLK
timestamp 1698175906
transform 1 0 14448 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__194__CLK
timestamp 1698175906
transform 1 0 15120 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__195__CLK
timestamp 1698175906
transform 1 0 23520 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__196__CLK
timestamp 1698175906
transform 1 0 19488 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__197__CLK
timestamp 1698175906
transform -1 0 21840 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__198__CLK
timestamp 1698175906
transform 1 0 15568 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__199__CLK
timestamp 1698175906
transform 1 0 14224 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__200__CLK
timestamp 1698175906
transform 1 0 17472 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__201__CLK
timestamp 1698175906
transform 1 0 30016 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__202__CLK
timestamp 1698175906
transform 1 0 26544 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__203__CLK
timestamp 1698175906
transform 1 0 25648 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__204__CLK
timestamp 1698175906
transform 1 0 25312 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__205__CLK
timestamp 1698175906
transform 1 0 27888 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__206__CLK
timestamp 1698175906
transform 1 0 27888 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__207__CLK
timestamp 1698175906
transform 1 0 24192 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__208__CLK
timestamp 1698175906
transform 1 0 29792 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__209__CLK
timestamp 1698175906
transform 1 0 18816 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__210__CLK
timestamp 1698175906
transform 1 0 16800 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__211__CLK
timestamp 1698175906
transform 1 0 26096 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__212__CLK
timestamp 1698175906
transform 1 0 17472 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__213__CLK
timestamp 1698175906
transform 1 0 17584 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__214__CLK
timestamp 1698175906
transform -1 0 23296 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__215__CLK
timestamp 1698175906
transform 1 0 29904 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform 1 0 18816 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19040 0 -1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 20720 0 1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 22960 0 1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16800 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_165 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19824 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_169
timestamp 1698175906
transform 1 0 20272 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_172
timestamp 1698175906
transform 1 0 20608 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_232
timestamp 1698175906
transform 1 0 27328 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_236 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 27776 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 28224 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 32032 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 35840 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 39648 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 40096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348
timestamp 1698175906
transform 1 0 40320 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_142
timestamp 1698175906
transform 1 0 17248 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_206
timestamp 1698175906
transform 1 0 24416 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_238
timestamp 1698175906
transform 1 0 28000 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_270 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 31584 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_278
timestamp 1698175906
transform 1 0 32480 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 32928 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 40096 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 40320 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 13328 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698175906
transform 1 0 21168 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 28336 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 36848 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 17248 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 25088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 32928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 40096 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 40320 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 21168 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 36848 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 32928 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 40096 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 40320 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 13328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 21168 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 36848 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 17248 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 25088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 32256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 32928 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 40096 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 40320 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 13328 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 21168 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 28336 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 29008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 36176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 36848 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 9408 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 17248 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 25088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 32256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 32928 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 40096 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 40320 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 13328 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 21168 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 29008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 36176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 36848 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 9408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 17248 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 24416 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 25088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 32928 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 40096 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 40320 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_107
timestamp 1698175906
transform 1 0 13328 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_171
timestamp 1698175906
transform 1 0 20496 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_177
timestamp 1698175906
transform 1 0 21168 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_183
timestamp 1698175906
transform 1 0 21840 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_215 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 25424 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_231
timestamp 1698175906
transform 1 0 27216 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_239
timestamp 1698175906
transform 1 0 28112 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_243
timestamp 1698175906
transform 1 0 28560 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 29008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 36848 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698175906
transform 1 0 9408 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698175906
transform 1 0 16576 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_142
timestamp 1698175906
transform 1 0 17248 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_150
timestamp 1698175906
transform 1 0 18144 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_212
timestamp 1698175906
transform 1 0 25088 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_216
timestamp 1698175906
transform 1 0 25536 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 32928 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 40096 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 40320 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_107
timestamp 1698175906
transform 1 0 13328 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_123
timestamp 1698175906
transform 1 0 15120 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_160
timestamp 1698175906
transform 1 0 19264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_164
timestamp 1698175906
transform 1 0 19712 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_172
timestamp 1698175906
transform 1 0 20608 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_174
timestamp 1698175906
transform 1 0 20832 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_177
timestamp 1698175906
transform 1 0 21168 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_185
timestamp 1698175906
transform 1 0 22064 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_189
timestamp 1698175906
transform 1 0 22512 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_219
timestamp 1698175906
transform 1 0 25872 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_223
timestamp 1698175906
transform 1 0 26320 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_239
timestamp 1698175906
transform 1 0 28112 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_243
timestamp 1698175906
transform 1 0 28560 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 29008 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 36176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 36848 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_72
timestamp 1698175906
transform 1 0 9408 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_104
timestamp 1698175906
transform 1 0 12992 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_108
timestamp 1698175906
transform 1 0 13440 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_110
timestamp 1698175906
transform 1 0 13664 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_142
timestamp 1698175906
transform 1 0 17248 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_146
timestamp 1698175906
transform 1 0 17696 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_162
timestamp 1698175906
transform 1 0 19488 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_182
timestamp 1698175906
transform 1 0 21728 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_196
timestamp 1698175906
transform 1 0 23296 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_204
timestamp 1698175906
transform 1 0 24192 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_208
timestamp 1698175906
transform 1 0 24640 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_216
timestamp 1698175906
transform 1 0 25536 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 32928 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698175906
transform 1 0 40096 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698175906
transform 1 0 40320 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_136
timestamp 1698175906
transform 1 0 16576 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_143
timestamp 1698175906
transform 1 0 17360 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_147
timestamp 1698175906
transform 1 0 17808 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_155
timestamp 1698175906
transform 1 0 18704 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_163
timestamp 1698175906
transform 1 0 19600 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_171
timestamp 1698175906
transform 1 0 20496 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_183
timestamp 1698175906
transform 1 0 21840 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_187
timestamp 1698175906
transform 1 0 22288 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_199
timestamp 1698175906
transform 1 0 23632 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_231
timestamp 1698175906
transform 1 0 27216 0 1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_239
timestamp 1698175906
transform 1 0 28112 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_243
timestamp 1698175906
transform 1 0 28560 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 29008 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 36176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_317
timestamp 1698175906
transform 1 0 36848 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698175906
transform 1 0 1568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698175906
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_72
timestamp 1698175906
transform 1 0 9408 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_88
timestamp 1698175906
transform 1 0 11200 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_125
timestamp 1698175906
transform 1 0 15344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_129
timestamp 1698175906
transform 1 0 15792 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_137
timestamp 1698175906
transform 1 0 16688 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_139
timestamp 1698175906
transform 1 0 16912 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_151
timestamp 1698175906
transform 1 0 18256 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_166
timestamp 1698175906
transform 1 0 19936 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_173
timestamp 1698175906
transform 1 0 20720 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_201
timestamp 1698175906
transform 1 0 23856 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1698175906
transform 1 0 24752 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_212
timestamp 1698175906
transform 1 0 25088 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_220
timestamp 1698175906
transform 1 0 25984 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_222
timestamp 1698175906
transform 1 0 26208 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_252
timestamp 1698175906
transform 1 0 29568 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_256
timestamp 1698175906
transform 1 0 30016 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_272
timestamp 1698175906
transform 1 0 31808 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_282
timestamp 1698175906
transform 1 0 32928 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_346
timestamp 1698175906
transform 1 0 40096 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_348
timestamp 1698175906
transform 1 0 40320 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_28
timestamp 1698175906
transform 1 0 4480 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_32
timestamp 1698175906
transform 1 0 4928 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698175906
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698175906
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_107
timestamp 1698175906
transform 1 0 13328 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_121
timestamp 1698175906
transform 1 0 14896 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_125
timestamp 1698175906
transform 1 0 15344 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_141
timestamp 1698175906
transform 1 0 17136 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_159
timestamp 1698175906
transform 1 0 19152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_166
timestamp 1698175906
transform 1 0 19936 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_174
timestamp 1698175906
transform 1 0 20832 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_177
timestamp 1698175906
transform 1 0 21168 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_179
timestamp 1698175906
transform 1 0 21392 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_186
timestamp 1698175906
transform 1 0 22176 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_188
timestamp 1698175906
transform 1 0 22400 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_195
timestamp 1698175906
transform 1 0 23184 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_235
timestamp 1698175906
transform 1 0 27664 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_239
timestamp 1698175906
transform 1 0 28112 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_244
timestamp 1698175906
transform 1 0 28672 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698175906
transform 1 0 29008 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698175906
transform 1 0 36176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_317
timestamp 1698175906
transform 1 0 36848 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_321
timestamp 1698175906
transform 1 0 37296 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698175906
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698175906
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_72
timestamp 1698175906
transform 1 0 9408 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_104
timestamp 1698175906
transform 1 0 12992 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_136
timestamp 1698175906
transform 1 0 16576 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_142
timestamp 1698175906
transform 1 0 17248 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_144
timestamp 1698175906
transform 1 0 17472 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_169
timestamp 1698175906
transform 1 0 20272 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_182
timestamp 1698175906
transform 1 0 21728 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_204
timestamp 1698175906
transform 1 0 24192 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_208
timestamp 1698175906
transform 1 0 24640 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_220
timestamp 1698175906
transform 1 0 25984 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_233
timestamp 1698175906
transform 1 0 27440 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_265
timestamp 1698175906
transform 1 0 31024 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_273
timestamp 1698175906
transform 1 0 31920 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_277
timestamp 1698175906
transform 1 0 32368 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_279
timestamp 1698175906
transform 1 0 32592 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_282
timestamp 1698175906
transform 1 0 32928 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_314
timestamp 1698175906
transform 1 0 36512 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_322
timestamp 1698175906
transform 1 0 37408 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_37
timestamp 1698175906
transform 1 0 5488 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_69
timestamp 1698175906
transform 1 0 9072 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_85
timestamp 1698175906
transform 1 0 10864 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_93
timestamp 1698175906
transform 1 0 11760 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_103
timestamp 1698175906
transform 1 0 12880 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_107
timestamp 1698175906
transform 1 0 13328 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_117
timestamp 1698175906
transform 1 0 14448 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_119
timestamp 1698175906
transform 1 0 14672 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_126
timestamp 1698175906
transform 1 0 15456 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_146
timestamp 1698175906
transform 1 0 17696 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_154
timestamp 1698175906
transform 1 0 18592 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_162
timestamp 1698175906
transform 1 0 19488 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_166
timestamp 1698175906
transform 1 0 19936 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_168
timestamp 1698175906
transform 1 0 20160 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_196
timestamp 1698175906
transform 1 0 23296 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_204
timestamp 1698175906
transform 1 0 24192 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_208
timestamp 1698175906
transform 1 0 24640 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_210
timestamp 1698175906
transform 1 0 24864 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_213
timestamp 1698175906
transform 1 0 25200 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_217
timestamp 1698175906
transform 1 0 25648 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_221
timestamp 1698175906
transform 1 0 26096 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_237
timestamp 1698175906
transform 1 0 27888 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698175906
transform 1 0 29008 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698175906
transform 1 0 36176 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_317
timestamp 1698175906
transform 1 0 36848 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698175906
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698175906
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_72
timestamp 1698175906
transform 1 0 9408 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_80
timestamp 1698175906
transform 1 0 10304 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_84
timestamp 1698175906
transform 1 0 10752 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_128
timestamp 1698175906
transform 1 0 15680 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_132
timestamp 1698175906
transform 1 0 16128 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_152
timestamp 1698175906
transform 1 0 18368 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_173
timestamp 1698175906
transform 1 0 20720 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_189
timestamp 1698175906
transform 1 0 22512 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_196
timestamp 1698175906
transform 1 0 23296 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_212
timestamp 1698175906
transform 1 0 25088 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_254
timestamp 1698175906
transform 1 0 29792 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_258
timestamp 1698175906
transform 1 0 30240 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_274
timestamp 1698175906
transform 1 0 32032 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_278
timestamp 1698175906
transform 1 0 32480 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_282
timestamp 1698175906
transform 1 0 32928 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_346
timestamp 1698175906
transform 1 0 40096 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_348
timestamp 1698175906
transform 1 0 40320 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698175906
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698175906
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_107
timestamp 1698175906
transform 1 0 13328 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_111
timestamp 1698175906
transform 1 0 13776 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_119
timestamp 1698175906
transform 1 0 14672 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_173
timestamp 1698175906
transform 1 0 20720 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_177
timestamp 1698175906
transform 1 0 21168 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_190
timestamp 1698175906
transform 1 0 22624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_192
timestamp 1698175906
transform 1 0 22848 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_243
timestamp 1698175906
transform 1 0 28560 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_259
timestamp 1698175906
transform 1 0 30352 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_263
timestamp 1698175906
transform 1 0 30800 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_295
timestamp 1698175906
transform 1 0 34384 0 1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698175906
transform 1 0 36176 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_317
timestamp 1698175906
transform 1 0 36848 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_321
timestamp 1698175906
transform 1 0 37296 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698175906
transform 1 0 1568 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698175906
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_72
timestamp 1698175906
transform 1 0 9408 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_80
timestamp 1698175906
transform 1 0 10304 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_84
timestamp 1698175906
transform 1 0 10752 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_115
timestamp 1698175906
transform 1 0 14224 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_124
timestamp 1698175906
transform 1 0 15232 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_154
timestamp 1698175906
transform 1 0 18592 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_208
timestamp 1698175906
transform 1 0 24640 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_253
timestamp 1698175906
transform 1 0 29680 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_257
timestamp 1698175906
transform 1 0 30128 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_273
timestamp 1698175906
transform 1 0 31920 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_277
timestamp 1698175906
transform 1 0 32368 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_279
timestamp 1698175906
transform 1 0 32592 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698175906
transform 1 0 32928 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_314
timestamp 1698175906
transform 1 0 36512 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_322
timestamp 1698175906
transform 1 0 37408 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698175906
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698175906
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698175906
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_107
timestamp 1698175906
transform 1 0 13328 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_121
timestamp 1698175906
transform 1 0 14896 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_125
timestamp 1698175906
transform 1 0 15344 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_133
timestamp 1698175906
transform 1 0 16240 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_137
timestamp 1698175906
transform 1 0 16688 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_162
timestamp 1698175906
transform 1 0 19488 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_223
timestamp 1698175906
transform 1 0 26320 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_227
timestamp 1698175906
transform 1 0 26768 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_235
timestamp 1698175906
transform 1 0 27664 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_241
timestamp 1698175906
transform 1 0 28336 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698175906
transform 1 0 29008 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 36176 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_317
timestamp 1698175906
transform 1 0 36848 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698175906
transform 1 0 37296 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_28
timestamp 1698175906
transform 1 0 4480 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_60
timestamp 1698175906
transform 1 0 8064 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_68
timestamp 1698175906
transform 1 0 8960 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_72
timestamp 1698175906
transform 1 0 9408 0 -1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_88
timestamp 1698175906
transform 1 0 11200 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_129
timestamp 1698175906
transform 1 0 15792 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_139
timestamp 1698175906
transform 1 0 16912 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_142
timestamp 1698175906
transform 1 0 17248 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_209
timestamp 1698175906
transform 1 0 24752 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_212
timestamp 1698175906
transform 1 0 25088 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_276
timestamp 1698175906
transform 1 0 32256 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_282
timestamp 1698175906
transform 1 0 32928 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_314
timestamp 1698175906
transform 1 0 36512 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_322
timestamp 1698175906
transform 1 0 37408 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_28
timestamp 1698175906
transform 1 0 4480 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_32
timestamp 1698175906
transform 1 0 4928 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698175906
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698175906
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_113
timestamp 1698175906
transform 1 0 14000 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_117
timestamp 1698175906
transform 1 0 14448 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_119
timestamp 1698175906
transform 1 0 14672 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_154
timestamp 1698175906
transform 1 0 18592 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_158
timestamp 1698175906
transform 1 0 19040 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_174
timestamp 1698175906
transform 1 0 20832 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_177
timestamp 1698175906
transform 1 0 21168 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_193
timestamp 1698175906
transform 1 0 22960 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_201
timestamp 1698175906
transform 1 0 23856 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_203
timestamp 1698175906
transform 1 0 24080 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_206
timestamp 1698175906
transform 1 0 24416 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_238
timestamp 1698175906
transform 1 0 28000 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_242
timestamp 1698175906
transform 1 0 28448 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_244
timestamp 1698175906
transform 1 0 28672 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 29008 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 36176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_317
timestamp 1698175906
transform 1 0 36848 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_28
timestamp 1698175906
transform 1 0 4480 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_60
timestamp 1698175906
transform 1 0 8064 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_68
timestamp 1698175906
transform 1 0 8960 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_72
timestamp 1698175906
transform 1 0 9408 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_136
timestamp 1698175906
transform 1 0 16576 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_142
timestamp 1698175906
transform 1 0 17248 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_174
timestamp 1698175906
transform 1 0 20832 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_183
timestamp 1698175906
transform 1 0 21840 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_191
timestamp 1698175906
transform 1 0 22736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_195
timestamp 1698175906
transform 1 0 23184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_197
timestamp 1698175906
transform 1 0 23408 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_204
timestamp 1698175906
transform 1 0 24192 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_208
timestamp 1698175906
transform 1 0 24640 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_221
timestamp 1698175906
transform 1 0 26096 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_226
timestamp 1698175906
transform 1 0 26656 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_258
timestamp 1698175906
transform 1 0 30240 0 -1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_274
timestamp 1698175906
transform 1 0 32032 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_278
timestamp 1698175906
transform 1 0 32480 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_282
timestamp 1698175906
transform 1 0 32928 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_346
timestamp 1698175906
transform 1 0 40096 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_348
timestamp 1698175906
transform 1 0 40320 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698175906
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_107
timestamp 1698175906
transform 1 0 13328 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_123
timestamp 1698175906
transform 1 0 15120 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_125
timestamp 1698175906
transform 1 0 15344 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_134
timestamp 1698175906
transform 1 0 16352 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_140
timestamp 1698175906
transform 1 0 17024 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_172
timestamp 1698175906
transform 1 0 20608 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_174
timestamp 1698175906
transform 1 0 20832 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_191
timestamp 1698175906
transform 1 0 22736 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_199
timestamp 1698175906
transform 1 0 23632 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_203
timestamp 1698175906
transform 1 0 24080 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_205
timestamp 1698175906
transform 1 0 24304 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_235
timestamp 1698175906
transform 1 0 27664 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_239
timestamp 1698175906
transform 1 0 28112 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_243
timestamp 1698175906
transform 1 0 28560 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 29008 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 36176 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_317
timestamp 1698175906
transform 1 0 36848 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_321
timestamp 1698175906
transform 1 0 37296 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2
timestamp 1698175906
transform 1 0 1568 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_66
timestamp 1698175906
transform 1 0 8736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_72
timestamp 1698175906
transform 1 0 9408 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_104
timestamp 1698175906
transform 1 0 12992 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_108
timestamp 1698175906
transform 1 0 13440 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_138
timestamp 1698175906
transform 1 0 16800 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_156
timestamp 1698175906
transform 1 0 18816 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_160
timestamp 1698175906
transform 1 0 19264 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_190
timestamp 1698175906
transform 1 0 22624 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_196
timestamp 1698175906
transform 1 0 23296 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_200
timestamp 1698175906
transform 1 0 23744 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_206
timestamp 1698175906
transform 1 0 24416 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_212
timestamp 1698175906
transform 1 0 25088 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_276
timestamp 1698175906
transform 1 0 32256 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_282
timestamp 1698175906
transform 1 0 32928 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_346
timestamp 1698175906
transform 1 0 40096 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_348
timestamp 1698175906
transform 1 0 40320 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698175906
transform 1 0 1568 0 1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_107
timestamp 1698175906
transform 1 0 13328 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_123
timestamp 1698175906
transform 1 0 15120 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_125
timestamp 1698175906
transform 1 0 15344 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_155
timestamp 1698175906
transform 1 0 18704 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_159
timestamp 1698175906
transform 1 0 19152 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_215
timestamp 1698175906
transform 1 0 25424 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_219
timestamp 1698175906
transform 1 0 25872 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_235
timestamp 1698175906
transform 1 0 27664 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_243
timestamp 1698175906
transform 1 0 28560 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 29008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 36176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_317
timestamp 1698175906
transform 1 0 36848 0 1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_333
timestamp 1698175906
transform 1 0 38640 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_341
timestamp 1698175906
transform 1 0 39536 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_72
timestamp 1698175906
transform 1 0 9408 0 -1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_104
timestamp 1698175906
transform 1 0 12992 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_120
timestamp 1698175906
transform 1 0 14784 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_138
timestamp 1698175906
transform 1 0 16800 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_142
timestamp 1698175906
transform 1 0 17248 0 -1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_158
timestamp 1698175906
transform 1 0 19040 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_162
timestamp 1698175906
transform 1 0 19488 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_192
timestamp 1698175906
transform 1 0 22848 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_196
timestamp 1698175906
transform 1 0 23296 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_204
timestamp 1698175906
transform 1 0 24192 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_208
timestamp 1698175906
transform 1 0 24640 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698175906
transform 1 0 25088 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698175906
transform 1 0 32256 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 32928 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 40096 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 40320 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698175906
transform 1 0 13328 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698175906
transform 1 0 20496 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698175906
transform 1 0 21168 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698175906
transform 1 0 28336 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 29008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 36176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 36848 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 9408 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 16576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 17248 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 24416 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 25088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 32256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 32928 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 40096 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 40320 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 13328 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 20496 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 21168 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 28336 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 29008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 36176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 36848 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_6
timestamp 1698175906
transform 1 0 2016 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 9408 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 17248 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 25088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 32928 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 40096 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 40320 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 13328 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 20496 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 21168 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 29008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 36176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 36848 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 9408 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 17248 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 24416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 25088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 32256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 32928 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 40096 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 40320 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 13328 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 20496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 21168 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 28336 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 29008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 36176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 36848 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 9408 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 16576 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 17248 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 24416 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 25088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 32256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 32928 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 40096 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 40320 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 13328 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 20496 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 21168 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 28336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 29008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 36176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 36848 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 9408 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 16576 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 17248 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 24416 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 25088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 32256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 32928 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 40096 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 40320 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_107
timestamp 1698175906
transform 1 0 13328 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_123
timestamp 1698175906
transform 1 0 15120 0 1 36064
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_131
timestamp 1698175906
transform 1 0 16016 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_42_159
timestamp 1698175906
transform 1 0 19152 0 1 36064
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698175906
transform 1 0 21168 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 28336 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 29008 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 36176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 36848 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 1568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 9408 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 16576 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_168
timestamp 1698175906
transform 1 0 20160 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_172
timestamp 1698175906
transform 1 0 20608 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_174
timestamp 1698175906
transform 1 0 20832 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_201
timestamp 1698175906
transform 1 0 23856 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 24752 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_238
timestamp 1698175906
transform 1 0 28000 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_270
timestamp 1698175906
transform 1 0 31584 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_278
timestamp 1698175906
transform 1 0 32480 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 32928 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 40096 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 40320 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_36
timestamp 1698175906
transform 1 0 5376 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_41
timestamp 1698175906
transform 1 0 5936 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_44_57
timestamp 1698175906
transform 1 0 7728 0 1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_65
timestamp 1698175906
transform 1 0 8624 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_67
timestamp 1698175906
transform 1 0 8848 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 9184 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 12992 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_138
timestamp 1698175906
transform 1 0 16800 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_142
timestamp 1698175906
transform 1 0 17248 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_172
timestamp 1698175906
transform 1 0 20608 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_176
timestamp 1698175906
transform 1 0 21056 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 27776 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_240
timestamp 1698175906
transform 1 0 28224 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_44_274
timestamp 1698175906
transform 1 0 32032 0 1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_290
timestamp 1698175906
transform 1 0 33824 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_294
timestamp 1698175906
transform 1 0 34272 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_299
timestamp 1698175906
transform 1 0 34832 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_303
timestamp 1698175906
transform 1 0 35280 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_305
timestamp 1698175906
transform 1 0 35504 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 35840 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 39648 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 40096 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 40320 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita44_22 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 5936 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita44_23
timestamp 1698175906
transform -1 0 2016 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita44_24
timestamp 1698175906
transform -1 0 34832 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita44_25
timestamp 1698175906
transform 1 0 39984 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__tieh  ita44_26 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 27776 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform 1 0 37520 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform 1 0 37520 0 -1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform 1 0 24416 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform 1 0 37520 0 1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform 1 0 16240 0 1 36064
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform 1 0 25088 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform 1 0 16912 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform -1 0 4480 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform 1 0 24416 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform 1 0 37520 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform -1 0 4480 0 -1 25088
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform 1 0 25088 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform 1 0 37520 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform 1 0 20944 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform 1 0 21280 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform -1 0 4480 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform 1 0 17472 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform -1 0 4480 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform 1 0 37520 0 1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform 1 0 37520 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 40656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 40656 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 40656 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 40656 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 40656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 40656 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 40656 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 40656 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 40656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 40656 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 40656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 40656 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 40656 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 40656 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 40656 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 40656 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 40656 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 40656 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 40656 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 40656 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 40656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 40656 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 40656 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 40656 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 40656 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 40656 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 40656 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 40656 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 40656 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 40656 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 40656 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 40656 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 40656 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 40656 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 40656 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 40656 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 40656 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 40656 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 40656 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 40656 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 40656 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 40656 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 40656 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 40656 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 40656 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 5152 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 8960 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 12768 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 16576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 20384 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 24192 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 28000 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 31808 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 35616 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 39424 0 1 37632
box -86 -86 310 870
<< labels >>
flabel metal3 s 0 26880 800 26992 0 FreeSans 448 0 0 0 clk
port 0 nsew signal input
flabel metal2 s 16800 41200 16912 42000 0 FreeSans 448 90 0 0 segm[0]
port 1 nsew signal tristate
flabel metal3 s 41200 22848 42000 22960 0 FreeSans 448 0 0 0 segm[10]
port 2 nsew signal tristate
flabel metal3 s 41200 18144 42000 18256 0 FreeSans 448 0 0 0 segm[11]
port 3 nsew signal tristate
flabel metal2 s 22848 41200 22960 42000 0 FreeSans 448 90 0 0 segm[12]
port 4 nsew signal tristate
flabel metal3 s 41200 24864 42000 24976 0 FreeSans 448 0 0 0 segm[13]
port 5 nsew signal tristate
flabel metal2 s 5376 41200 5488 42000 0 FreeSans 448 90 0 0 segm[1]
port 6 nsew signal tristate
flabel metal3 s 0 30240 800 30352 0 FreeSans 448 0 0 0 segm[2]
port 7 nsew signal tristate
flabel metal2 s 16128 41200 16240 42000 0 FreeSans 448 90 0 0 segm[3]
port 8 nsew signal tristate
flabel metal2 s 34272 41200 34384 42000 0 FreeSans 448 90 0 0 segm[4]
port 9 nsew signal tristate
flabel metal3 s 41200 26880 42000 26992 0 FreeSans 448 0 0 0 segm[5]
port 10 nsew signal tristate
flabel metal2 s 24864 0 24976 800 0 FreeSans 448 90 0 0 segm[6]
port 11 nsew signal tristate
flabel metal2 s 16800 0 16912 800 0 FreeSans 448 90 0 0 segm[7]
port 12 nsew signal tristate
flabel metal2 s 26208 41200 26320 42000 0 FreeSans 448 90 0 0 segm[8]
port 13 nsew signal tristate
flabel metal3 s 0 16800 800 16912 0 FreeSans 448 0 0 0 segm[9]
port 14 nsew signal tristate
flabel metal2 s 23520 0 23632 800 0 FreeSans 448 90 0 0 sel[0]
port 15 nsew signal tristate
flabel metal3 s 41200 17472 42000 17584 0 FreeSans 448 0 0 0 sel[10]
port 16 nsew signal tristate
flabel metal3 s 0 24192 800 24304 0 FreeSans 448 0 0 0 sel[11]
port 17 nsew signal tristate
flabel metal2 s 24864 41200 24976 42000 0 FreeSans 448 90 0 0 sel[1]
port 18 nsew signal tristate
flabel metal3 s 41200 22176 42000 22288 0 FreeSans 448 0 0 0 sel[2]
port 19 nsew signal tristate
flabel metal2 s 20832 41200 20944 42000 0 FreeSans 448 90 0 0 sel[3]
port 20 nsew signal tristate
flabel metal2 s 22176 41200 22288 42000 0 FreeSans 448 90 0 0 sel[4]
port 21 nsew signal tristate
flabel metal3 s 0 22848 800 22960 0 FreeSans 448 0 0 0 sel[5]
port 22 nsew signal tristate
flabel metal2 s 18144 41200 18256 42000 0 FreeSans 448 90 0 0 sel[6]
port 23 nsew signal tristate
flabel metal3 s 0 23520 800 23632 0 FreeSans 448 0 0 0 sel[7]
port 24 nsew signal tristate
flabel metal3 s 41200 20832 42000 20944 0 FreeSans 448 0 0 0 sel[8]
port 25 nsew signal tristate
flabel metal3 s 41200 21504 42000 21616 0 FreeSans 448 0 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 4448 3076 4768 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 35168 3076 35488 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 19808 3076 20128 38476 0 FreeSans 1280 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 21000 38416 21000 38416 0 vdd
rlabel metal1 21000 37632 21000 37632 0 vss
rlabel metal3 17472 26152 17472 26152 0 _000_
rlabel metal2 13272 22120 13272 22120 0 _001_
rlabel metal2 14392 22792 14392 22792 0 _002_
rlabel metal2 21224 25592 21224 25592 0 _003_
rlabel metal2 25816 19712 25816 19712 0 _004_
rlabel metal2 20664 14056 20664 14056 0 _005_
rlabel metal2 13048 17752 13048 17752 0 _006_
rlabel metal2 12376 19488 12376 19488 0 _007_
rlabel metal3 20160 22456 20160 22456 0 _008_
rlabel metal3 28448 20552 28448 20552 0 _009_
rlabel metal2 25368 22008 25368 22008 0 _010_
rlabel metal2 22960 26936 22960 26936 0 _011_
rlabel metal2 22568 14476 22568 14476 0 _012_
rlabel metal3 24528 17528 24528 17528 0 _013_
rlabel metal2 25592 25144 25592 25144 0 _014_
rlabel metal2 22008 21952 22008 21952 0 _015_
rlabel metal2 27160 16968 27160 16968 0 _016_
rlabel metal2 16296 23576 16296 23576 0 _017_
rlabel metal2 15960 25704 15960 25704 0 _018_
rlabel metal2 23520 14616 23520 14616 0 _019_
rlabel metal2 14728 15736 14728 15736 0 _020_
rlabel metal2 14280 16800 14280 16800 0 _021_
rlabel metal2 21672 27440 21672 27440 0 _022_
rlabel metal2 26936 21056 26936 21056 0 _023_
rlabel metal3 23576 24808 23576 24808 0 _024_
rlabel metal2 21560 22288 21560 22288 0 _025_
rlabel metal3 20720 22232 20720 22232 0 _026_
rlabel metal2 29960 20440 29960 20440 0 _027_
rlabel metal2 30408 20776 30408 20776 0 _028_
rlabel metal2 29288 21056 29288 21056 0 _029_
rlabel metal2 23240 19320 23240 19320 0 _030_
rlabel metal3 25200 21784 25200 21784 0 _031_
rlabel metal2 21616 26936 21616 26936 0 _032_
rlabel metal3 23520 26264 23520 26264 0 _033_
rlabel metal2 22792 16240 22792 16240 0 _034_
rlabel metal2 23912 17920 23912 17920 0 _035_
rlabel metal2 22008 16968 22008 16968 0 _036_
rlabel metal2 23240 16240 23240 16240 0 _037_
rlabel metal3 22008 20552 22008 20552 0 _038_
rlabel metal2 23352 16464 23352 16464 0 _039_
rlabel metal2 22960 15288 22960 15288 0 _040_
rlabel metal2 24248 18088 24248 18088 0 _041_
rlabel metal2 25984 24472 25984 24472 0 _042_
rlabel metal2 22456 21448 22456 21448 0 _043_
rlabel metal2 28280 17864 28280 17864 0 _044_
rlabel metal2 16632 23520 16632 23520 0 _045_
rlabel metal2 15848 26544 15848 26544 0 _046_
rlabel metal3 24416 15512 24416 15512 0 _047_
rlabel metal2 17304 16464 17304 16464 0 _048_
rlabel metal2 17864 17248 17864 17248 0 _049_
rlabel metal2 14056 17640 14056 17640 0 _050_
rlabel metal2 22456 25760 22456 25760 0 _051_
rlabel metal2 28056 21280 28056 21280 0 _052_
rlabel metal2 16968 19600 16968 19600 0 _053_
rlabel metal2 19264 17416 19264 17416 0 _054_
rlabel metal2 21560 18816 21560 18816 0 _055_
rlabel metal2 20216 17360 20216 17360 0 _056_
rlabel metal2 18200 18200 18200 18200 0 _057_
rlabel metal3 18480 22232 18480 22232 0 _058_
rlabel metal2 15624 18592 15624 18592 0 _059_
rlabel metal2 20104 18592 20104 18592 0 _060_
rlabel metal2 18648 26096 18648 26096 0 _061_
rlabel metal3 19936 20104 19936 20104 0 _062_
rlabel metal2 17304 20888 17304 20888 0 _063_
rlabel metal2 15064 23632 15064 23632 0 _064_
rlabel metal2 16632 18592 16632 18592 0 _065_
rlabel metal2 18312 22288 18312 22288 0 _066_
rlabel metal2 18088 26040 18088 26040 0 _067_
rlabel metal2 14560 20776 14560 20776 0 _068_
rlabel metal3 16968 18200 16968 18200 0 _069_
rlabel metal2 15008 17416 15008 17416 0 _070_
rlabel metal2 14840 21336 14840 21336 0 _071_
rlabel metal2 13832 23128 13832 23128 0 _072_
rlabel metal3 20608 15400 20608 15400 0 _073_
rlabel metal2 18088 21784 18088 21784 0 _074_
rlabel metal3 17920 21784 17920 21784 0 _075_
rlabel metal2 14728 22736 14728 22736 0 _076_
rlabel metal2 22904 17472 22904 17472 0 _077_
rlabel metal3 22288 18648 22288 18648 0 _078_
rlabel metal2 18200 23912 18200 23912 0 _079_
rlabel metal2 22120 26152 22120 26152 0 _080_
rlabel metal2 21672 25368 21672 25368 0 _081_
rlabel metal2 16408 19656 16408 19656 0 _082_
rlabel metal2 20888 16016 20888 16016 0 _083_
rlabel metal2 21840 17640 21840 17640 0 _084_
rlabel metal2 21336 17472 21336 17472 0 _085_
rlabel metal2 20272 14504 20272 14504 0 _086_
rlabel metal2 14952 18424 14952 18424 0 _087_
rlabel metal2 16184 18704 16184 18704 0 _088_
rlabel metal2 16240 20104 16240 20104 0 _089_
rlabel metal2 12712 19488 12712 19488 0 _090_
rlabel metal2 24472 20048 24472 20048 0 _091_
rlabel metal3 28224 18648 28224 18648 0 _092_
rlabel metal3 22120 22120 22120 22120 0 _093_
rlabel metal2 20888 20384 20888 20384 0 _094_
rlabel metal3 19992 16968 19992 16968 0 _095_
rlabel metal3 2478 26936 2478 26936 0 clk
rlabel metal2 23128 21112 23128 21112 0 clknet_0_clk
rlabel metal2 14952 24584 14952 24584 0 clknet_1_0__leaf_clk
rlabel metal2 23240 27384 23240 27384 0 clknet_1_1__leaf_clk
rlabel metal2 19152 14616 19152 14616 0 dut44.count\[0\]
rlabel metal2 18648 13608 18648 13608 0 dut44.count\[1\]
rlabel metal2 16632 17304 16632 17304 0 dut44.count\[2\]
rlabel metal2 14056 19488 14056 19488 0 dut44.count\[3\]
rlabel metal3 16968 28056 16968 28056 0 net1
rlabel metal2 24584 5964 24584 5964 0 net10
rlabel metal2 29400 17192 29400 17192 0 net11
rlabel metal2 17864 24360 17864 24360 0 net12
rlabel metal2 25256 32200 25256 32200 0 net13
rlabel metal2 37912 22792 37912 22792 0 net14
rlabel metal2 20944 31920 20944 31920 0 net15
rlabel metal3 22120 38024 22120 38024 0 net16
rlabel metal2 11816 23072 11816 23072 0 net17
rlabel metal3 18088 27160 18088 27160 0 net18
rlabel metal2 11144 22680 11144 22680 0 net19
rlabel metal3 31920 23072 31920 23072 0 net2
rlabel metal2 29512 21392 29512 21392 0 net20
rlabel metal2 28168 21840 28168 21840 0 net21
rlabel metal2 5544 37912 5544 37912 0 net22
rlabel metal3 1246 30296 1246 30296 0 net23
rlabel metal2 34440 37912 34440 37912 0 net24
rlabel metal3 40264 26880 40264 26880 0 net25
rlabel metal3 26880 38248 26880 38248 0 net26
rlabel metal3 29708 17752 29708 17752 0 net3
rlabel metal3 23632 27720 23632 27720 0 net4
rlabel metal2 27496 25200 27496 25200 0 net5
rlabel metal2 15960 28000 15960 28000 0 net6
rlabel metal2 25256 6356 25256 6356 0 net7
rlabel metal2 17080 5964 17080 5964 0 net8
rlabel metal2 14616 17584 14616 17584 0 net9
rlabel metal2 16856 39354 16856 39354 0 segm[0]
rlabel metal3 40642 22904 40642 22904 0 segm[10]
rlabel metal3 40642 18200 40642 18200 0 segm[11]
rlabel metal2 22904 39746 22904 39746 0 segm[12]
rlabel metal2 40040 25256 40040 25256 0 segm[13]
rlabel metal2 16184 38962 16184 38962 0 segm[3]
rlabel metal2 24920 2422 24920 2422 0 segm[6]
rlabel metal2 16856 2086 16856 2086 0 segm[7]
rlabel metal3 1358 16856 1358 16856 0 segm[9]
rlabel metal2 23576 2198 23576 2198 0 sel[0]
rlabel metal2 40040 17640 40040 17640 0 sel[10]
rlabel metal3 1358 24248 1358 24248 0 sel[11]
rlabel metal2 24920 39354 24920 39354 0 sel[1]
rlabel metal2 40040 22344 40040 22344 0 sel[2]
rlabel metal2 20888 39354 20888 39354 0 sel[3]
rlabel metal2 22232 39746 22232 39746 0 sel[4]
rlabel metal3 1358 22904 1358 22904 0 sel[5]
rlabel metal2 18200 39746 18200 39746 0 sel[6]
rlabel metal3 1358 23576 1358 23576 0 sel[7]
rlabel metal3 40642 20888 40642 20888 0 sel[8]
rlabel metal2 40040 21504 40040 21504 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 42000 42000
<< end >>
