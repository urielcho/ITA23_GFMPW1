magic
tech gf180mcuD
magscale 1 5
timestamp 1699642150
<< metal1 >>
rect 672 19221 20328 19238
rect 672 19195 2239 19221
rect 2265 19195 2291 19221
rect 2317 19195 2343 19221
rect 2369 19195 17599 19221
rect 17625 19195 17651 19221
rect 17677 19195 17703 19221
rect 17729 19195 20328 19221
rect 672 19178 20328 19195
rect 9591 19137 9617 19143
rect 9591 19105 9617 19111
rect 11215 19137 11241 19143
rect 11215 19105 11241 19111
rect 12783 19137 12809 19143
rect 12783 19105 12809 19111
rect 9865 18999 9871 19025
rect 9897 18999 9903 19025
rect 10705 18999 10711 19025
rect 10737 18999 10743 19025
rect 12273 18999 12279 19025
rect 12305 18999 12311 19025
rect 10543 18969 10569 18975
rect 10543 18937 10569 18943
rect 672 18829 20328 18846
rect 672 18803 9919 18829
rect 9945 18803 9971 18829
rect 9997 18803 10023 18829
rect 10049 18803 20328 18829
rect 672 18786 20328 18803
rect 9367 18745 9393 18751
rect 9367 18713 9393 18719
rect 11047 18745 11073 18751
rect 11047 18713 11073 18719
rect 8857 18607 8863 18633
rect 8889 18607 8895 18633
rect 10761 18607 10767 18633
rect 10793 18607 10799 18633
rect 672 18437 20328 18454
rect 672 18411 2239 18437
rect 2265 18411 2291 18437
rect 2317 18411 2343 18437
rect 2369 18411 17599 18437
rect 17625 18411 17651 18437
rect 17677 18411 17703 18437
rect 17729 18411 20328 18437
rect 672 18394 20328 18411
rect 672 18045 20328 18062
rect 672 18019 9919 18045
rect 9945 18019 9971 18045
rect 9997 18019 10023 18045
rect 10049 18019 20328 18045
rect 672 18002 20328 18019
rect 672 17653 20328 17670
rect 672 17627 2239 17653
rect 2265 17627 2291 17653
rect 2317 17627 2343 17653
rect 2369 17627 17599 17653
rect 17625 17627 17651 17653
rect 17677 17627 17703 17653
rect 17729 17627 20328 17653
rect 672 17610 20328 17627
rect 20119 17345 20145 17351
rect 20119 17313 20145 17319
rect 672 17261 20328 17278
rect 672 17235 9919 17261
rect 9945 17235 9971 17261
rect 9997 17235 10023 17261
rect 10049 17235 20328 17261
rect 672 17218 20328 17235
rect 672 16869 20328 16886
rect 672 16843 2239 16869
rect 2265 16843 2291 16869
rect 2317 16843 2343 16869
rect 2369 16843 17599 16869
rect 17625 16843 17651 16869
rect 17677 16843 17703 16869
rect 17729 16843 20328 16869
rect 672 16826 20328 16843
rect 672 16477 20328 16494
rect 672 16451 9919 16477
rect 9945 16451 9971 16477
rect 9997 16451 10023 16477
rect 10049 16451 20328 16477
rect 672 16434 20328 16451
rect 672 16085 20328 16102
rect 672 16059 2239 16085
rect 2265 16059 2291 16085
rect 2317 16059 2343 16085
rect 2369 16059 17599 16085
rect 17625 16059 17651 16085
rect 17677 16059 17703 16085
rect 17729 16059 20328 16085
rect 672 16042 20328 16059
rect 672 15693 20328 15710
rect 672 15667 9919 15693
rect 9945 15667 9971 15693
rect 9997 15667 10023 15693
rect 10049 15667 20328 15693
rect 672 15650 20328 15667
rect 672 15301 20328 15318
rect 672 15275 2239 15301
rect 2265 15275 2291 15301
rect 2317 15275 2343 15301
rect 2369 15275 17599 15301
rect 17625 15275 17651 15301
rect 17677 15275 17703 15301
rect 17729 15275 20328 15301
rect 672 15258 20328 15275
rect 672 14909 20328 14926
rect 672 14883 9919 14909
rect 9945 14883 9971 14909
rect 9997 14883 10023 14909
rect 10049 14883 20328 14909
rect 672 14866 20328 14883
rect 672 14517 20328 14534
rect 672 14491 2239 14517
rect 2265 14491 2291 14517
rect 2317 14491 2343 14517
rect 2369 14491 17599 14517
rect 17625 14491 17651 14517
rect 17677 14491 17703 14517
rect 17729 14491 20328 14517
rect 672 14474 20328 14491
rect 672 14125 20328 14142
rect 672 14099 9919 14125
rect 9945 14099 9971 14125
rect 9997 14099 10023 14125
rect 10049 14099 20328 14125
rect 672 14082 20328 14099
rect 11159 14041 11185 14047
rect 11159 14009 11185 14015
rect 10985 13959 10991 13985
rect 11017 13959 11023 13985
rect 9417 13903 9423 13929
rect 9449 13903 9455 13929
rect 11439 13873 11465 13879
rect 9753 13847 9759 13873
rect 9785 13847 9791 13873
rect 10817 13847 10823 13873
rect 10849 13847 10855 13873
rect 11439 13841 11465 13847
rect 672 13733 20328 13750
rect 672 13707 2239 13733
rect 2265 13707 2291 13733
rect 2317 13707 2343 13733
rect 2369 13707 17599 13733
rect 17625 13707 17651 13733
rect 17677 13707 17703 13733
rect 17729 13707 20328 13733
rect 672 13690 20328 13707
rect 9983 13649 10009 13655
rect 9983 13617 10009 13623
rect 10375 13593 10401 13599
rect 9809 13567 9815 13593
rect 9841 13567 9847 13593
rect 10375 13561 10401 13567
rect 20007 13593 20033 13599
rect 20007 13561 20033 13567
rect 13455 13537 13481 13543
rect 8409 13511 8415 13537
rect 8441 13511 8447 13537
rect 9977 13511 9983 13537
rect 10009 13511 10015 13537
rect 18825 13511 18831 13537
rect 18857 13511 18863 13537
rect 13455 13505 13481 13511
rect 10151 13481 10177 13487
rect 8745 13455 8751 13481
rect 8777 13455 8783 13481
rect 10151 13449 10177 13455
rect 10599 13481 10625 13487
rect 10599 13449 10625 13455
rect 10711 13481 10737 13487
rect 10711 13449 10737 13455
rect 10767 13481 10793 13487
rect 10767 13449 10793 13455
rect 13399 13481 13425 13487
rect 13399 13449 13425 13455
rect 12447 13425 12473 13431
rect 12447 13393 12473 13399
rect 672 13341 20328 13358
rect 672 13315 9919 13341
rect 9945 13315 9971 13341
rect 9997 13315 10023 13341
rect 10049 13315 20328 13341
rect 672 13298 20328 13315
rect 8751 13257 8777 13263
rect 8751 13225 8777 13231
rect 9535 13257 9561 13263
rect 9535 13225 9561 13231
rect 10207 13257 10233 13263
rect 10207 13225 10233 13231
rect 10263 13257 10289 13263
rect 10263 13225 10289 13231
rect 14239 13257 14265 13263
rect 14239 13225 14265 13231
rect 9479 13201 9505 13207
rect 14401 13175 14407 13201
rect 14433 13175 14439 13201
rect 9479 13169 9505 13175
rect 9647 13145 9673 13151
rect 2137 13119 2143 13145
rect 2169 13119 2175 13145
rect 6953 13119 6959 13145
rect 6985 13119 6991 13145
rect 9647 13113 9673 13119
rect 9759 13145 9785 13151
rect 9759 13113 9785 13119
rect 10151 13145 10177 13151
rect 10151 13113 10177 13119
rect 10319 13145 10345 13151
rect 10319 13113 10345 13119
rect 10375 13145 10401 13151
rect 10649 13119 10655 13145
rect 10681 13119 10687 13145
rect 12609 13119 12615 13145
rect 12641 13119 12647 13145
rect 18825 13119 18831 13145
rect 18857 13119 18863 13145
rect 10375 13113 10401 13119
rect 12335 13089 12361 13095
rect 7345 13063 7351 13089
rect 7377 13063 7383 13089
rect 8409 13063 8415 13089
rect 8441 13063 8447 13089
rect 11041 13063 11047 13089
rect 11073 13063 11079 13089
rect 12105 13063 12111 13089
rect 12137 13063 12143 13089
rect 13001 13063 13007 13089
rect 13033 13063 13039 13089
rect 14065 13063 14071 13089
rect 14097 13063 14103 13089
rect 19945 13063 19951 13089
rect 19977 13063 19983 13089
rect 12335 13057 12361 13063
rect 967 13033 993 13039
rect 967 13001 993 13007
rect 672 12949 20328 12966
rect 672 12923 2239 12949
rect 2265 12923 2291 12949
rect 2317 12923 2343 12949
rect 2369 12923 17599 12949
rect 17625 12923 17651 12949
rect 17677 12923 17703 12949
rect 17729 12923 20328 12949
rect 672 12906 20328 12923
rect 20007 12809 20033 12815
rect 1017 12783 1023 12809
rect 1049 12783 1055 12809
rect 12497 12783 12503 12809
rect 12529 12783 12535 12809
rect 14121 12783 14127 12809
rect 14153 12783 14159 12809
rect 20007 12777 20033 12783
rect 10823 12753 10849 12759
rect 2137 12727 2143 12753
rect 2169 12727 2175 12753
rect 10823 12721 10849 12727
rect 10935 12753 10961 12759
rect 11327 12753 11353 12759
rect 11041 12727 11047 12753
rect 11073 12727 11079 12753
rect 10935 12721 10961 12727
rect 11327 12721 11353 12727
rect 11495 12753 11521 12759
rect 12441 12727 12447 12753
rect 12473 12727 12479 12753
rect 12665 12727 12671 12753
rect 12697 12727 12703 12753
rect 18825 12727 18831 12753
rect 18857 12727 18863 12753
rect 11495 12721 11521 12727
rect 7071 12697 7097 12703
rect 7071 12665 7097 12671
rect 8135 12697 8161 12703
rect 8135 12665 8161 12671
rect 8303 12697 8329 12703
rect 8303 12665 8329 12671
rect 11215 12697 11241 12703
rect 11215 12665 11241 12671
rect 12223 12697 12249 12703
rect 12223 12665 12249 12671
rect 12279 12697 12305 12703
rect 13057 12671 13063 12697
rect 13089 12671 13095 12697
rect 12279 12665 12305 12671
rect 6959 12641 6985 12647
rect 6959 12609 6985 12615
rect 7015 12641 7041 12647
rect 7015 12609 7041 12615
rect 10991 12641 11017 12647
rect 10991 12609 11017 12615
rect 11271 12641 11297 12647
rect 11271 12609 11297 12615
rect 11943 12641 11969 12647
rect 11943 12609 11969 12615
rect 12111 12641 12137 12647
rect 12111 12609 12137 12615
rect 672 12557 20328 12574
rect 672 12531 9919 12557
rect 9945 12531 9971 12557
rect 9997 12531 10023 12557
rect 10049 12531 20328 12557
rect 672 12514 20328 12531
rect 7631 12473 7657 12479
rect 12727 12473 12753 12479
rect 9417 12447 9423 12473
rect 9449 12447 9455 12473
rect 7631 12441 7657 12447
rect 12727 12441 12753 12447
rect 7799 12417 7825 12423
rect 7009 12391 7015 12417
rect 7041 12391 7047 12417
rect 7799 12385 7825 12391
rect 8807 12417 8833 12423
rect 8807 12385 8833 12391
rect 8975 12417 9001 12423
rect 12839 12417 12865 12423
rect 9361 12391 9367 12417
rect 9393 12391 9399 12417
rect 10089 12391 10095 12417
rect 10121 12391 10127 12417
rect 10649 12391 10655 12417
rect 10681 12391 10687 12417
rect 8975 12385 9001 12391
rect 12839 12385 12865 12391
rect 12895 12417 12921 12423
rect 13623 12417 13649 12423
rect 12945 12391 12951 12417
rect 12977 12391 12983 12417
rect 12895 12385 12921 12391
rect 13623 12385 13649 12391
rect 13679 12417 13705 12423
rect 13679 12385 13705 12391
rect 8919 12361 8945 12367
rect 7401 12335 7407 12361
rect 7433 12335 7439 12361
rect 8919 12329 8945 12335
rect 9031 12361 9057 12367
rect 10823 12361 10849 12367
rect 9137 12335 9143 12361
rect 9169 12335 9175 12361
rect 9641 12335 9647 12361
rect 9673 12335 9679 12361
rect 9809 12335 9815 12361
rect 9841 12335 9847 12361
rect 9031 12329 9057 12335
rect 10823 12329 10849 12335
rect 5945 12279 5951 12305
rect 5977 12279 5983 12305
rect 13113 12279 13119 12305
rect 13145 12279 13151 12305
rect 7855 12249 7881 12255
rect 7855 12217 7881 12223
rect 672 12165 20328 12182
rect 672 12139 2239 12165
rect 2265 12139 2291 12165
rect 2317 12139 2343 12165
rect 2369 12139 17599 12165
rect 17625 12139 17651 12165
rect 17677 12139 17703 12165
rect 17729 12139 20328 12165
rect 672 12122 20328 12139
rect 7183 12081 7209 12087
rect 7183 12049 7209 12055
rect 10151 12081 10177 12087
rect 10151 12049 10177 12055
rect 10711 12081 10737 12087
rect 10711 12049 10737 12055
rect 12951 12081 12977 12087
rect 12951 12049 12977 12055
rect 6735 12025 6761 12031
rect 6735 11993 6761 11999
rect 6791 11969 6817 11975
rect 6791 11937 6817 11943
rect 6903 11969 6929 11975
rect 6903 11937 6929 11943
rect 7295 11969 7321 11975
rect 7295 11937 7321 11943
rect 7687 11969 7713 11975
rect 7687 11937 7713 11943
rect 7855 11969 7881 11975
rect 10145 11943 10151 11969
rect 10177 11943 10183 11969
rect 11657 11943 11663 11969
rect 11689 11943 11695 11969
rect 7855 11937 7881 11943
rect 7407 11913 7433 11919
rect 7065 11887 7071 11913
rect 7097 11887 7103 11913
rect 7407 11881 7433 11887
rect 7575 11913 7601 11919
rect 7575 11881 7601 11887
rect 9983 11913 10009 11919
rect 9983 11881 10009 11887
rect 10655 11913 10681 11919
rect 10655 11881 10681 11887
rect 11439 11913 11465 11919
rect 11439 11881 11465 11887
rect 13007 11913 13033 11919
rect 13007 11881 13033 11887
rect 7183 11857 7209 11863
rect 7183 11825 7209 11831
rect 7631 11857 7657 11863
rect 7631 11825 7657 11831
rect 10711 11857 10737 11863
rect 10711 11825 10737 11831
rect 11271 11857 11297 11863
rect 11271 11825 11297 11831
rect 11327 11857 11353 11863
rect 11327 11825 11353 11831
rect 11383 11857 11409 11863
rect 11383 11825 11409 11831
rect 12951 11857 12977 11863
rect 12951 11825 12977 11831
rect 672 11773 20328 11790
rect 672 11747 9919 11773
rect 9945 11747 9971 11773
rect 9997 11747 10023 11773
rect 10049 11747 20328 11773
rect 672 11730 20328 11747
rect 7127 11689 7153 11695
rect 7127 11657 7153 11663
rect 7407 11689 7433 11695
rect 7407 11657 7433 11663
rect 8247 11689 8273 11695
rect 8689 11663 8695 11689
rect 8721 11663 8727 11689
rect 8247 11657 8273 11663
rect 7631 11633 7657 11639
rect 6505 11607 6511 11633
rect 6537 11607 6543 11633
rect 7631 11601 7657 11607
rect 8359 11633 8385 11639
rect 13735 11633 13761 11639
rect 9193 11607 9199 11633
rect 9225 11607 9231 11633
rect 10425 11607 10431 11633
rect 10457 11607 10463 11633
rect 8359 11601 8385 11607
rect 13735 11601 13761 11607
rect 7351 11577 7377 11583
rect 6897 11551 6903 11577
rect 6929 11551 6935 11577
rect 7351 11545 7377 11551
rect 7519 11577 7545 11583
rect 7519 11545 7545 11551
rect 7855 11577 7881 11583
rect 7855 11545 7881 11551
rect 8415 11577 8441 11583
rect 8415 11545 8441 11551
rect 8863 11577 8889 11583
rect 8863 11545 8889 11551
rect 9031 11577 9057 11583
rect 13511 11577 13537 11583
rect 9529 11551 9535 11577
rect 9561 11551 9567 11577
rect 9031 11545 9057 11551
rect 13511 11545 13537 11551
rect 13623 11577 13649 11583
rect 18825 11551 18831 11577
rect 18857 11551 18863 11577
rect 13623 11545 13649 11551
rect 13567 11521 13593 11527
rect 5441 11495 5447 11521
rect 5473 11495 5479 11521
rect 13567 11489 13593 11495
rect 20007 11465 20033 11471
rect 20007 11433 20033 11439
rect 672 11381 20328 11398
rect 672 11355 2239 11381
rect 2265 11355 2291 11381
rect 2317 11355 2343 11381
rect 2369 11355 17599 11381
rect 17625 11355 17651 11381
rect 17677 11355 17703 11381
rect 17729 11355 20328 11381
rect 672 11338 20328 11355
rect 6791 11241 6817 11247
rect 5385 11215 5391 11241
rect 5417 11215 5423 11241
rect 6449 11215 6455 11241
rect 6481 11215 6487 11241
rect 6791 11209 6817 11215
rect 8807 11241 8833 11247
rect 8807 11209 8833 11215
rect 9759 11241 9785 11247
rect 9759 11209 9785 11215
rect 10095 11241 10121 11247
rect 12559 11241 12585 11247
rect 20007 11241 20033 11247
rect 11265 11215 11271 11241
rect 11297 11215 11303 11241
rect 12329 11215 12335 11241
rect 12361 11215 12367 11241
rect 14289 11215 14295 11241
rect 14321 11215 14327 11241
rect 10095 11209 10121 11215
rect 12559 11209 12585 11215
rect 20007 11209 20033 11215
rect 7295 11185 7321 11191
rect 5049 11159 5055 11185
rect 5081 11159 5087 11185
rect 7295 11153 7321 11159
rect 9087 11185 9113 11191
rect 9087 11153 9113 11159
rect 9479 11185 9505 11191
rect 10929 11159 10935 11185
rect 10961 11159 10967 11185
rect 12889 11159 12895 11185
rect 12921 11159 12927 11185
rect 13225 11159 13231 11185
rect 13257 11159 13263 11185
rect 18825 11159 18831 11185
rect 18857 11159 18863 11185
rect 9479 11153 9505 11159
rect 6959 11129 6985 11135
rect 6959 11097 6985 11103
rect 7127 11129 7153 11135
rect 7127 11097 7153 11103
rect 8975 11129 9001 11135
rect 8975 11097 9001 11103
rect 9703 11129 9729 11135
rect 9703 11097 9729 11103
rect 10263 11129 10289 11135
rect 10263 11097 10289 11103
rect 8527 11073 8553 11079
rect 9815 11073 9841 11079
rect 7457 11047 7463 11073
rect 7489 11047 7495 11073
rect 9249 11047 9255 11073
rect 9281 11047 9287 11073
rect 8527 11041 8553 11047
rect 9815 11041 9841 11047
rect 10039 11073 10065 11079
rect 10039 11041 10065 11047
rect 10151 11073 10177 11079
rect 10151 11041 10177 11047
rect 672 10989 20328 11006
rect 672 10963 9919 10989
rect 9945 10963 9971 10989
rect 9997 10963 10023 10989
rect 10049 10963 20328 10989
rect 672 10946 20328 10963
rect 7519 10905 7545 10911
rect 7519 10873 7545 10879
rect 8303 10905 8329 10911
rect 8303 10873 8329 10879
rect 8919 10905 8945 10911
rect 8919 10873 8945 10879
rect 9255 10905 9281 10911
rect 11999 10905 12025 10911
rect 9255 10873 9281 10879
rect 10711 10877 10737 10883
rect 7071 10849 7097 10855
rect 7071 10817 7097 10823
rect 8695 10849 8721 10855
rect 8695 10817 8721 10823
rect 8751 10849 8777 10855
rect 8751 10817 8777 10823
rect 9031 10849 9057 10855
rect 9871 10849 9897 10855
rect 11999 10873 12025 10879
rect 12671 10905 12697 10911
rect 12671 10873 12697 10879
rect 13343 10905 13369 10911
rect 13343 10873 13369 10879
rect 9417 10823 9423 10849
rect 9449 10823 9455 10849
rect 10369 10823 10375 10849
rect 10401 10823 10407 10849
rect 10711 10845 10737 10851
rect 12055 10849 12081 10855
rect 11713 10823 11719 10849
rect 11745 10823 11751 10849
rect 9031 10817 9057 10823
rect 9871 10817 9897 10823
rect 12055 10817 12081 10823
rect 12111 10849 12137 10855
rect 12111 10817 12137 10823
rect 13455 10849 13481 10855
rect 13455 10817 13481 10823
rect 13567 10849 13593 10855
rect 13567 10817 13593 10823
rect 8135 10793 8161 10799
rect 8017 10767 8023 10793
rect 8049 10767 8055 10793
rect 8135 10761 8161 10767
rect 9087 10793 9113 10799
rect 9087 10761 9113 10767
rect 9647 10793 9673 10799
rect 9647 10761 9673 10767
rect 9703 10793 9729 10799
rect 10655 10793 10681 10799
rect 10257 10767 10263 10793
rect 10289 10767 10295 10793
rect 9703 10761 9729 10767
rect 10655 10761 10681 10767
rect 10935 10793 10961 10799
rect 11943 10793 11969 10799
rect 13287 10793 13313 10799
rect 11209 10767 11215 10793
rect 11241 10767 11247 10793
rect 11545 10767 11551 10793
rect 11577 10767 11583 10793
rect 12329 10767 12335 10793
rect 12361 10767 12367 10793
rect 18825 10767 18831 10793
rect 18857 10767 18863 10793
rect 10935 10761 10961 10767
rect 11943 10761 11969 10767
rect 13287 10761 13313 10767
rect 6567 10737 6593 10743
rect 7631 10737 7657 10743
rect 7457 10711 7463 10737
rect 7489 10711 7495 10737
rect 11657 10711 11663 10737
rect 11689 10711 11695 10737
rect 19945 10711 19951 10737
rect 19977 10711 19983 10737
rect 6567 10705 6593 10711
rect 7631 10705 7657 10711
rect 7127 10681 7153 10687
rect 7127 10649 7153 10655
rect 8751 10681 8777 10687
rect 8751 10649 8777 10655
rect 9815 10681 9841 10687
rect 9815 10649 9841 10655
rect 10711 10681 10737 10687
rect 10711 10649 10737 10655
rect 672 10597 20328 10614
rect 672 10571 2239 10597
rect 2265 10571 2291 10597
rect 2317 10571 2343 10597
rect 2369 10571 17599 10597
rect 17625 10571 17651 10597
rect 17677 10571 17703 10597
rect 17729 10571 20328 10597
rect 672 10554 20328 10571
rect 10823 10513 10849 10519
rect 7737 10487 7743 10513
rect 7769 10487 7775 10513
rect 10823 10481 10849 10487
rect 6847 10457 6873 10463
rect 5385 10431 5391 10457
rect 5417 10431 5423 10457
rect 6449 10431 6455 10457
rect 6481 10431 6487 10457
rect 6847 10425 6873 10431
rect 8247 10457 8273 10463
rect 8247 10425 8273 10431
rect 10039 10457 10065 10463
rect 10039 10425 10065 10431
rect 12671 10457 12697 10463
rect 20007 10457 20033 10463
rect 14289 10431 14295 10457
rect 14321 10431 14327 10457
rect 12671 10425 12697 10431
rect 20007 10425 20033 10431
rect 6903 10401 6929 10407
rect 7407 10401 7433 10407
rect 10095 10401 10121 10407
rect 5049 10375 5055 10401
rect 5081 10375 5087 10401
rect 7121 10375 7127 10401
rect 7153 10375 7159 10401
rect 7513 10375 7519 10401
rect 7545 10375 7551 10401
rect 9025 10375 9031 10401
rect 9057 10375 9063 10401
rect 9585 10375 9591 10401
rect 9617 10375 9623 10401
rect 6903 10369 6929 10375
rect 7407 10369 7433 10375
rect 10095 10369 10121 10375
rect 10207 10401 10233 10407
rect 10207 10369 10233 10375
rect 11047 10401 11073 10407
rect 11047 10369 11073 10375
rect 11383 10401 11409 10407
rect 11383 10369 11409 10375
rect 11831 10401 11857 10407
rect 11993 10375 11999 10401
rect 12025 10375 12031 10401
rect 12833 10375 12839 10401
rect 12865 10375 12871 10401
rect 14625 10375 14631 10401
rect 14657 10375 14663 10401
rect 18825 10375 18831 10401
rect 18857 10375 18863 10401
rect 11831 10369 11857 10375
rect 7967 10345 7993 10351
rect 9983 10345 10009 10351
rect 7233 10319 7239 10345
rect 7265 10319 7271 10345
rect 9081 10319 9087 10345
rect 9113 10319 9119 10345
rect 7967 10313 7993 10319
rect 9983 10313 10009 10319
rect 10655 10345 10681 10351
rect 12111 10345 12137 10351
rect 11209 10319 11215 10345
rect 11241 10319 11247 10345
rect 11545 10319 11551 10345
rect 11577 10319 11583 10345
rect 13225 10319 13231 10345
rect 13257 10319 13263 10345
rect 10655 10313 10681 10319
rect 12111 10313 12137 10319
rect 8863 10289 8889 10295
rect 10767 10289 10793 10295
rect 9473 10263 9479 10289
rect 9505 10263 9511 10289
rect 8863 10257 8889 10263
rect 10767 10257 10793 10263
rect 12167 10289 12193 10295
rect 14737 10263 14743 10289
rect 14769 10263 14775 10289
rect 12167 10257 12193 10263
rect 672 10205 20328 10222
rect 672 10179 9919 10205
rect 9945 10179 9971 10205
rect 9997 10179 10023 10205
rect 10049 10179 20328 10205
rect 672 10162 20328 10179
rect 7463 10121 7489 10127
rect 7463 10089 7489 10095
rect 12951 10121 12977 10127
rect 12951 10089 12977 10095
rect 6735 10065 6761 10071
rect 6735 10033 6761 10039
rect 7911 10065 7937 10071
rect 13567 10065 13593 10071
rect 8857 10039 8863 10065
rect 8889 10039 8895 10065
rect 10145 10039 10151 10065
rect 10177 10039 10183 10065
rect 7911 10033 7937 10039
rect 13567 10033 13593 10039
rect 13791 10065 13817 10071
rect 13791 10033 13817 10039
rect 7743 10009 7769 10015
rect 7743 9977 7769 9983
rect 8079 10009 8105 10015
rect 8079 9977 8105 9983
rect 8695 10009 8721 10015
rect 12895 10009 12921 10015
rect 9025 9983 9031 10009
rect 9057 9983 9063 10009
rect 8695 9977 8721 9983
rect 12895 9977 12921 9983
rect 13007 10009 13033 10015
rect 13007 9977 13033 9983
rect 13231 10009 13257 10015
rect 13673 9983 13679 10009
rect 13705 9983 13711 10009
rect 13231 9977 13257 9983
rect 11943 9953 11969 9959
rect 8129 9927 8135 9953
rect 8161 9927 8167 9953
rect 11943 9921 11969 9927
rect 12783 9953 12809 9959
rect 12783 9921 12809 9927
rect 13623 9953 13649 9959
rect 13623 9921 13649 9927
rect 672 9813 20328 9830
rect 672 9787 2239 9813
rect 2265 9787 2291 9813
rect 2317 9787 2343 9813
rect 2369 9787 17599 9813
rect 17625 9787 17651 9813
rect 17677 9787 17703 9813
rect 17729 9787 20328 9813
rect 672 9770 20328 9787
rect 8135 9729 8161 9735
rect 8135 9697 8161 9703
rect 9143 9729 9169 9735
rect 9753 9703 9759 9729
rect 9785 9703 9791 9729
rect 9143 9697 9169 9703
rect 20007 9673 20033 9679
rect 9641 9647 9647 9673
rect 9673 9647 9679 9673
rect 10257 9647 10263 9673
rect 10289 9647 10295 9673
rect 11545 9647 11551 9673
rect 11577 9647 11583 9673
rect 20007 9641 20033 9647
rect 7799 9617 7825 9623
rect 7799 9585 7825 9591
rect 8303 9617 8329 9623
rect 10711 9617 10737 9623
rect 11943 9617 11969 9623
rect 8969 9591 8975 9617
rect 9001 9591 9007 9617
rect 9193 9591 9199 9617
rect 9225 9591 9231 9617
rect 9585 9591 9591 9617
rect 9617 9591 9623 9617
rect 10089 9591 10095 9617
rect 10121 9591 10127 9617
rect 10201 9591 10207 9617
rect 10233 9591 10239 9617
rect 11657 9591 11663 9617
rect 11689 9591 11695 9617
rect 8303 9585 8329 9591
rect 10711 9585 10737 9591
rect 11943 9585 11969 9591
rect 12111 9617 12137 9623
rect 12111 9585 12137 9591
rect 12895 9617 12921 9623
rect 12895 9585 12921 9591
rect 13231 9617 13257 9623
rect 18825 9591 18831 9617
rect 18857 9591 18863 9617
rect 13231 9585 13257 9591
rect 8415 9561 8441 9567
rect 7961 9535 7967 9561
rect 7993 9535 7999 9561
rect 8415 9529 8441 9535
rect 8863 9561 8889 9567
rect 12391 9561 12417 9567
rect 10929 9535 10935 9561
rect 10961 9535 10967 9561
rect 11097 9535 11103 9561
rect 11129 9535 11135 9561
rect 8863 9529 8889 9535
rect 12391 9529 12417 9535
rect 13119 9561 13145 9567
rect 13119 9529 13145 9535
rect 13567 9561 13593 9567
rect 13567 9529 13593 9535
rect 13679 9561 13705 9567
rect 13679 9529 13705 9535
rect 13735 9561 13761 9567
rect 13735 9529 13761 9535
rect 9087 9505 9113 9511
rect 9087 9473 9113 9479
rect 10319 9505 10345 9511
rect 11719 9505 11745 9511
rect 10705 9479 10711 9505
rect 10737 9479 10743 9505
rect 10319 9473 10345 9479
rect 11719 9473 11745 9479
rect 11999 9505 12025 9511
rect 13063 9505 13089 9511
rect 12553 9479 12559 9505
rect 12585 9479 12591 9505
rect 11999 9473 12025 9479
rect 13063 9473 13089 9479
rect 672 9421 20328 9438
rect 672 9395 9919 9421
rect 9945 9395 9971 9421
rect 9997 9395 10023 9421
rect 10049 9395 20328 9421
rect 672 9378 20328 9395
rect 9703 9337 9729 9343
rect 9703 9305 9729 9311
rect 10543 9337 10569 9343
rect 10543 9305 10569 9311
rect 10655 9337 10681 9343
rect 11383 9337 11409 9343
rect 11041 9311 11047 9337
rect 11073 9311 11079 9337
rect 10655 9305 10681 9311
rect 11383 9305 11409 9311
rect 11495 9337 11521 9343
rect 11495 9305 11521 9311
rect 7687 9281 7713 9287
rect 7687 9249 7713 9255
rect 9255 9281 9281 9287
rect 13225 9255 13231 9281
rect 13257 9255 13263 9281
rect 9255 9249 9281 9255
rect 7855 9225 7881 9231
rect 5889 9199 5895 9225
rect 5921 9199 5927 9225
rect 6225 9199 6231 9225
rect 6257 9199 6263 9225
rect 7855 9193 7881 9199
rect 7967 9225 7993 9231
rect 7967 9193 7993 9199
rect 8135 9225 8161 9231
rect 9871 9225 9897 9231
rect 8969 9199 8975 9225
rect 9001 9199 9007 9225
rect 8135 9193 8161 9199
rect 9871 9193 9897 9199
rect 10879 9225 10905 9231
rect 10879 9193 10905 9199
rect 11215 9225 11241 9231
rect 11215 9193 11241 9199
rect 11439 9225 11465 9231
rect 11439 9193 11465 9199
rect 11719 9225 11745 9231
rect 12833 9199 12839 9225
rect 12865 9199 12871 9225
rect 11719 9193 11745 9199
rect 7575 9169 7601 9175
rect 7289 9143 7295 9169
rect 7321 9143 7327 9169
rect 7575 9137 7601 9143
rect 7743 9169 7769 9175
rect 10599 9169 10625 9175
rect 8353 9143 8359 9169
rect 8385 9143 8391 9169
rect 7743 9137 7769 9143
rect 10599 9137 10625 9143
rect 12727 9169 12753 9175
rect 14289 9143 14295 9169
rect 14321 9143 14327 9169
rect 12727 9137 12753 9143
rect 672 9029 20328 9046
rect 672 9003 2239 9029
rect 2265 9003 2291 9029
rect 2317 9003 2343 9029
rect 2369 9003 17599 9029
rect 17625 9003 17651 9029
rect 17677 9003 17703 9029
rect 17729 9003 20328 9029
rect 672 8986 20328 9003
rect 10823 8945 10849 8951
rect 10823 8913 10849 8919
rect 9647 8889 9673 8895
rect 9647 8857 9673 8863
rect 10431 8889 10457 8895
rect 10431 8857 10457 8863
rect 20007 8889 20033 8895
rect 20007 8857 20033 8863
rect 10375 8833 10401 8839
rect 7513 8807 7519 8833
rect 7545 8807 7551 8833
rect 8409 8807 8415 8833
rect 8441 8807 8447 8833
rect 8745 8807 8751 8833
rect 8777 8807 8783 8833
rect 10375 8801 10401 8807
rect 11159 8833 11185 8839
rect 11159 8801 11185 8807
rect 11663 8833 11689 8839
rect 11663 8801 11689 8807
rect 13007 8833 13033 8839
rect 13007 8801 13033 8807
rect 13231 8833 13257 8839
rect 13231 8801 13257 8807
rect 13343 8833 13369 8839
rect 13343 8801 13369 8807
rect 13567 8833 13593 8839
rect 13567 8801 13593 8807
rect 13623 8833 13649 8839
rect 18825 8807 18831 8833
rect 18857 8807 18863 8833
rect 13623 8801 13649 8807
rect 7631 8777 7657 8783
rect 7631 8745 7657 8751
rect 7967 8777 7993 8783
rect 10711 8777 10737 8783
rect 8521 8751 8527 8777
rect 8553 8751 8559 8777
rect 8857 8751 8863 8777
rect 8889 8751 8895 8777
rect 9865 8751 9871 8777
rect 9897 8751 9903 8777
rect 10089 8751 10095 8777
rect 10121 8751 10127 8777
rect 11321 8751 11327 8777
rect 11353 8751 11359 8777
rect 7967 8745 7993 8751
rect 10711 8745 10737 8751
rect 8023 8721 8049 8727
rect 8023 8689 8049 8695
rect 8079 8721 8105 8727
rect 8079 8689 8105 8695
rect 9031 8721 9057 8727
rect 9367 8721 9393 8727
rect 13175 8721 13201 8727
rect 9193 8695 9199 8721
rect 9225 8695 9231 8721
rect 10985 8695 10991 8721
rect 11017 8695 11023 8721
rect 11825 8695 11831 8721
rect 11857 8695 11863 8721
rect 9031 8689 9057 8695
rect 9367 8689 9393 8695
rect 13175 8689 13201 8695
rect 13511 8721 13537 8727
rect 13511 8689 13537 8695
rect 13735 8721 13761 8727
rect 13735 8689 13761 8695
rect 672 8637 20328 8654
rect 672 8611 9919 8637
rect 9945 8611 9971 8637
rect 9997 8611 10023 8637
rect 10049 8611 20328 8637
rect 672 8594 20328 8611
rect 8359 8553 8385 8559
rect 8359 8521 8385 8527
rect 8751 8553 8777 8559
rect 8751 8521 8777 8527
rect 8303 8497 8329 8503
rect 6449 8471 6455 8497
rect 6481 8471 6487 8497
rect 8303 8465 8329 8471
rect 8695 8497 8721 8503
rect 8695 8465 8721 8471
rect 9199 8497 9225 8503
rect 9199 8465 9225 8471
rect 9255 8497 9281 8503
rect 10929 8471 10935 8497
rect 10961 8471 10967 8497
rect 13225 8471 13231 8497
rect 13257 8471 13263 8497
rect 9255 8465 9281 8471
rect 7743 8441 7769 8447
rect 6057 8415 6063 8441
rect 6089 8415 6095 8441
rect 7743 8409 7769 8415
rect 9367 8441 9393 8447
rect 9473 8415 9479 8441
rect 9505 8415 9511 8441
rect 12833 8415 12839 8441
rect 12865 8415 12871 8441
rect 9367 8409 9393 8415
rect 12671 8385 12697 8391
rect 7513 8359 7519 8385
rect 7545 8359 7551 8385
rect 14289 8359 14295 8385
rect 14321 8359 14327 8385
rect 12671 8353 12697 8359
rect 672 8245 20328 8262
rect 672 8219 2239 8245
rect 2265 8219 2291 8245
rect 2317 8219 2343 8245
rect 2369 8219 17599 8245
rect 17625 8219 17651 8245
rect 17677 8219 17703 8245
rect 17729 8219 20328 8245
rect 672 8202 20328 8219
rect 9479 8161 9505 8167
rect 8857 8135 8863 8161
rect 8889 8135 8895 8161
rect 9479 8129 9505 8135
rect 20007 8105 20033 8111
rect 20007 8073 20033 8079
rect 8975 8049 9001 8055
rect 8745 8023 8751 8049
rect 8777 8023 8783 8049
rect 8975 8017 9001 8023
rect 9143 8049 9169 8055
rect 9423 8049 9449 8055
rect 9305 8023 9311 8049
rect 9337 8023 9343 8049
rect 9143 8017 9169 8023
rect 9423 8017 9449 8023
rect 10039 8049 10065 8055
rect 10039 8017 10065 8023
rect 10263 8049 10289 8055
rect 10263 8017 10289 8023
rect 10375 8049 10401 8055
rect 10767 8049 10793 8055
rect 13063 8049 13089 8055
rect 10649 8023 10655 8049
rect 10681 8023 10687 8049
rect 10985 8023 10991 8049
rect 11017 8023 11023 8049
rect 10375 8017 10401 8023
rect 10767 8017 10793 8023
rect 13063 8017 13089 8023
rect 13287 8049 13313 8055
rect 13287 8017 13313 8023
rect 13455 8049 13481 8055
rect 13455 8017 13481 8023
rect 13623 8049 13649 8055
rect 18825 8023 18831 8049
rect 18857 8023 18863 8049
rect 13623 8017 13649 8023
rect 10151 7993 10177 7999
rect 10151 7961 10177 7967
rect 12951 7993 12977 7999
rect 12951 7961 12977 7967
rect 9087 7937 9113 7943
rect 9087 7905 9113 7911
rect 9983 7937 10009 7943
rect 9983 7905 10009 7911
rect 10823 7937 10849 7943
rect 10823 7905 10849 7911
rect 10879 7937 10905 7943
rect 10879 7905 10905 7911
rect 13175 7937 13201 7943
rect 13175 7905 13201 7911
rect 13567 7937 13593 7943
rect 13567 7905 13593 7911
rect 672 7853 20328 7870
rect 672 7827 9919 7853
rect 9945 7827 9971 7853
rect 9997 7827 10023 7853
rect 10049 7827 20328 7853
rect 672 7810 20328 7827
rect 8751 7769 8777 7775
rect 8751 7737 8777 7743
rect 10207 7769 10233 7775
rect 10207 7737 10233 7743
rect 10319 7769 10345 7775
rect 10319 7737 10345 7743
rect 11887 7769 11913 7775
rect 11887 7737 11913 7743
rect 10095 7713 10121 7719
rect 10095 7681 10121 7687
rect 11831 7713 11857 7719
rect 11831 7681 11857 7687
rect 11943 7713 11969 7719
rect 13169 7687 13175 7713
rect 13201 7687 13207 7713
rect 11943 7681 11969 7687
rect 8975 7657 9001 7663
rect 7009 7631 7015 7657
rect 7041 7631 7047 7657
rect 8975 7625 9001 7631
rect 9087 7657 9113 7663
rect 9087 7625 9113 7631
rect 9703 7657 9729 7663
rect 9703 7625 9729 7631
rect 9815 7657 9841 7663
rect 9815 7625 9841 7631
rect 12335 7657 12361 7663
rect 12777 7631 12783 7657
rect 12809 7631 12815 7657
rect 12335 7625 12361 7631
rect 8919 7601 8945 7607
rect 7345 7575 7351 7601
rect 7377 7575 7383 7601
rect 8409 7575 8415 7601
rect 8441 7575 8447 7601
rect 8919 7569 8945 7575
rect 9143 7601 9169 7607
rect 14233 7575 14239 7601
rect 14265 7575 14271 7601
rect 9143 7569 9169 7575
rect 10151 7545 10177 7551
rect 9529 7519 9535 7545
rect 9561 7519 9567 7545
rect 10151 7513 10177 7519
rect 672 7461 20328 7478
rect 672 7435 2239 7461
rect 2265 7435 2291 7461
rect 2317 7435 2343 7461
rect 2369 7435 17599 7461
rect 17625 7435 17651 7461
rect 17677 7435 17703 7461
rect 17729 7435 20328 7461
rect 672 7418 20328 7435
rect 10039 7377 10065 7383
rect 10039 7345 10065 7351
rect 10151 7377 10177 7383
rect 10151 7345 10177 7351
rect 12783 7377 12809 7383
rect 12783 7345 12809 7351
rect 9087 7321 9113 7327
rect 12447 7321 12473 7327
rect 8857 7295 8863 7321
rect 8889 7295 8895 7321
rect 11153 7295 11159 7321
rect 11185 7295 11191 7321
rect 12217 7295 12223 7321
rect 12249 7295 12255 7321
rect 9087 7289 9113 7295
rect 12447 7289 12473 7295
rect 10263 7265 10289 7271
rect 7401 7239 7407 7265
rect 7433 7239 7439 7265
rect 10369 7239 10375 7265
rect 10401 7239 10407 7265
rect 10817 7239 10823 7265
rect 10849 7239 10855 7265
rect 10263 7233 10289 7239
rect 7793 7183 7799 7209
rect 7825 7183 7831 7209
rect 10319 7153 10345 7159
rect 10319 7121 10345 7127
rect 12839 7153 12865 7159
rect 12839 7121 12865 7127
rect 12895 7153 12921 7159
rect 12895 7121 12921 7127
rect 672 7069 20328 7086
rect 672 7043 9919 7069
rect 9945 7043 9971 7069
rect 9997 7043 10023 7069
rect 10049 7043 20328 7069
rect 672 7026 20328 7043
rect 9143 6985 9169 6991
rect 9143 6953 9169 6959
rect 11271 6985 11297 6991
rect 11271 6953 11297 6959
rect 8303 6929 8329 6935
rect 8303 6897 8329 6903
rect 8975 6929 9001 6935
rect 8975 6897 9001 6903
rect 9927 6929 9953 6935
rect 9927 6897 9953 6903
rect 10151 6929 10177 6935
rect 10151 6897 10177 6903
rect 10207 6929 10233 6935
rect 10207 6897 10233 6903
rect 12783 6929 12809 6935
rect 12783 6897 12809 6903
rect 8415 6873 8441 6879
rect 8415 6841 8441 6847
rect 9087 6873 9113 6879
rect 9087 6841 9113 6847
rect 9311 6873 9337 6879
rect 9311 6841 9337 6847
rect 9647 6873 9673 6879
rect 9647 6841 9673 6847
rect 9759 6873 9785 6879
rect 9759 6841 9785 6847
rect 10039 6873 10065 6879
rect 10039 6841 10065 6847
rect 11215 6873 11241 6879
rect 11377 6847 11383 6873
rect 11409 6847 11415 6873
rect 12609 6847 12615 6873
rect 12641 6847 12647 6873
rect 11215 6841 11241 6847
rect 9871 6817 9897 6823
rect 8241 6791 8247 6817
rect 8273 6791 8279 6817
rect 9871 6785 9897 6791
rect 12615 6761 12641 6767
rect 12615 6729 12641 6735
rect 672 6677 20328 6694
rect 672 6651 2239 6677
rect 2265 6651 2291 6677
rect 2317 6651 2343 6677
rect 2369 6651 17599 6677
rect 17625 6651 17651 6677
rect 17677 6651 17703 6677
rect 17729 6651 20328 6677
rect 672 6634 20328 6651
rect 10319 6537 10345 6543
rect 9025 6511 9031 6537
rect 9057 6511 9063 6537
rect 10089 6511 10095 6537
rect 10121 6511 10127 6537
rect 10319 6505 10345 6511
rect 11831 6537 11857 6543
rect 12385 6511 12391 6537
rect 12417 6511 12423 6537
rect 13449 6511 13455 6537
rect 13481 6511 13487 6537
rect 11831 6505 11857 6511
rect 8689 6455 8695 6481
rect 8721 6455 8727 6481
rect 10761 6455 10767 6481
rect 10793 6455 10799 6481
rect 11993 6455 11999 6481
rect 12025 6455 12031 6481
rect 10655 6369 10681 6375
rect 10655 6337 10681 6343
rect 672 6285 20328 6302
rect 672 6259 9919 6285
rect 9945 6259 9971 6285
rect 9997 6259 10023 6285
rect 10049 6259 20328 6285
rect 672 6242 20328 6259
rect 11887 6201 11913 6207
rect 11887 6169 11913 6175
rect 10593 6119 10599 6145
rect 10625 6119 10631 6145
rect 10257 6063 10263 6089
rect 10289 6063 10295 6089
rect 11657 6007 11663 6033
rect 11689 6007 11695 6033
rect 672 5893 20328 5910
rect 672 5867 2239 5893
rect 2265 5867 2291 5893
rect 2317 5867 2343 5893
rect 2369 5867 17599 5893
rect 17625 5867 17651 5893
rect 17677 5867 17703 5893
rect 17729 5867 20328 5893
rect 672 5850 20328 5867
rect 672 5501 20328 5518
rect 672 5475 9919 5501
rect 9945 5475 9971 5501
rect 9997 5475 10023 5501
rect 10049 5475 20328 5501
rect 672 5458 20328 5475
rect 672 5109 20328 5126
rect 672 5083 2239 5109
rect 2265 5083 2291 5109
rect 2317 5083 2343 5109
rect 2369 5083 17599 5109
rect 17625 5083 17651 5109
rect 17677 5083 17703 5109
rect 17729 5083 20328 5109
rect 672 5066 20328 5083
rect 672 4717 20328 4734
rect 672 4691 9919 4717
rect 9945 4691 9971 4717
rect 9997 4691 10023 4717
rect 10049 4691 20328 4717
rect 672 4674 20328 4691
rect 672 4325 20328 4342
rect 672 4299 2239 4325
rect 2265 4299 2291 4325
rect 2317 4299 2343 4325
rect 2369 4299 17599 4325
rect 17625 4299 17651 4325
rect 17677 4299 17703 4325
rect 17729 4299 20328 4325
rect 672 4282 20328 4299
rect 672 3933 20328 3950
rect 672 3907 9919 3933
rect 9945 3907 9971 3933
rect 9997 3907 10023 3933
rect 10049 3907 20328 3933
rect 672 3890 20328 3907
rect 672 3541 20328 3558
rect 672 3515 2239 3541
rect 2265 3515 2291 3541
rect 2317 3515 2343 3541
rect 2369 3515 17599 3541
rect 17625 3515 17651 3541
rect 17677 3515 17703 3541
rect 17729 3515 20328 3541
rect 672 3498 20328 3515
rect 672 3149 20328 3166
rect 672 3123 9919 3149
rect 9945 3123 9971 3149
rect 9997 3123 10023 3149
rect 10049 3123 20328 3149
rect 672 3106 20328 3123
rect 672 2757 20328 2774
rect 672 2731 2239 2757
rect 2265 2731 2291 2757
rect 2317 2731 2343 2757
rect 2369 2731 17599 2757
rect 17625 2731 17651 2757
rect 17677 2731 17703 2757
rect 17729 2731 20328 2757
rect 672 2714 20328 2731
rect 672 2365 20328 2382
rect 672 2339 9919 2365
rect 9945 2339 9971 2365
rect 9997 2339 10023 2365
rect 10049 2339 20328 2365
rect 672 2322 20328 2339
rect 8857 2143 8863 2169
rect 8889 2143 8895 2169
rect 12665 2143 12671 2169
rect 12697 2143 12703 2169
rect 9367 2057 9393 2063
rect 9367 2025 9393 2031
rect 13119 2057 13145 2063
rect 13119 2025 13145 2031
rect 672 1973 20328 1990
rect 672 1947 2239 1973
rect 2265 1947 2291 1973
rect 2317 1947 2343 1973
rect 2369 1947 17599 1973
rect 17625 1947 17651 1973
rect 17677 1947 17703 1973
rect 17729 1947 20328 1973
rect 672 1930 20328 1947
rect 9311 1833 9337 1839
rect 9311 1801 9337 1807
rect 12783 1833 12809 1839
rect 12783 1801 12809 1807
rect 14687 1833 14713 1839
rect 14687 1801 14713 1807
rect 9025 1751 9031 1777
rect 9057 1751 9063 1777
rect 10369 1751 10375 1777
rect 10401 1751 10407 1777
rect 12273 1751 12279 1777
rect 12305 1751 12311 1777
rect 14289 1751 14295 1777
rect 14321 1751 14327 1777
rect 3487 1665 3513 1671
rect 3487 1633 3513 1639
rect 10879 1665 10905 1671
rect 10879 1633 10905 1639
rect 672 1581 20328 1598
rect 672 1555 9919 1581
rect 9945 1555 9971 1581
rect 9997 1555 10023 1581
rect 10049 1555 20328 1581
rect 672 1538 20328 1555
<< via1 >>
rect 2239 19195 2265 19221
rect 2291 19195 2317 19221
rect 2343 19195 2369 19221
rect 17599 19195 17625 19221
rect 17651 19195 17677 19221
rect 17703 19195 17729 19221
rect 9591 19111 9617 19137
rect 11215 19111 11241 19137
rect 12783 19111 12809 19137
rect 9871 18999 9897 19025
rect 10711 18999 10737 19025
rect 12279 18999 12305 19025
rect 10543 18943 10569 18969
rect 9919 18803 9945 18829
rect 9971 18803 9997 18829
rect 10023 18803 10049 18829
rect 9367 18719 9393 18745
rect 11047 18719 11073 18745
rect 8863 18607 8889 18633
rect 10767 18607 10793 18633
rect 2239 18411 2265 18437
rect 2291 18411 2317 18437
rect 2343 18411 2369 18437
rect 17599 18411 17625 18437
rect 17651 18411 17677 18437
rect 17703 18411 17729 18437
rect 9919 18019 9945 18045
rect 9971 18019 9997 18045
rect 10023 18019 10049 18045
rect 2239 17627 2265 17653
rect 2291 17627 2317 17653
rect 2343 17627 2369 17653
rect 17599 17627 17625 17653
rect 17651 17627 17677 17653
rect 17703 17627 17729 17653
rect 20119 17319 20145 17345
rect 9919 17235 9945 17261
rect 9971 17235 9997 17261
rect 10023 17235 10049 17261
rect 2239 16843 2265 16869
rect 2291 16843 2317 16869
rect 2343 16843 2369 16869
rect 17599 16843 17625 16869
rect 17651 16843 17677 16869
rect 17703 16843 17729 16869
rect 9919 16451 9945 16477
rect 9971 16451 9997 16477
rect 10023 16451 10049 16477
rect 2239 16059 2265 16085
rect 2291 16059 2317 16085
rect 2343 16059 2369 16085
rect 17599 16059 17625 16085
rect 17651 16059 17677 16085
rect 17703 16059 17729 16085
rect 9919 15667 9945 15693
rect 9971 15667 9997 15693
rect 10023 15667 10049 15693
rect 2239 15275 2265 15301
rect 2291 15275 2317 15301
rect 2343 15275 2369 15301
rect 17599 15275 17625 15301
rect 17651 15275 17677 15301
rect 17703 15275 17729 15301
rect 9919 14883 9945 14909
rect 9971 14883 9997 14909
rect 10023 14883 10049 14909
rect 2239 14491 2265 14517
rect 2291 14491 2317 14517
rect 2343 14491 2369 14517
rect 17599 14491 17625 14517
rect 17651 14491 17677 14517
rect 17703 14491 17729 14517
rect 9919 14099 9945 14125
rect 9971 14099 9997 14125
rect 10023 14099 10049 14125
rect 11159 14015 11185 14041
rect 10991 13959 11017 13985
rect 9423 13903 9449 13929
rect 9759 13847 9785 13873
rect 10823 13847 10849 13873
rect 11439 13847 11465 13873
rect 2239 13707 2265 13733
rect 2291 13707 2317 13733
rect 2343 13707 2369 13733
rect 17599 13707 17625 13733
rect 17651 13707 17677 13733
rect 17703 13707 17729 13733
rect 9983 13623 10009 13649
rect 9815 13567 9841 13593
rect 10375 13567 10401 13593
rect 20007 13567 20033 13593
rect 8415 13511 8441 13537
rect 9983 13511 10009 13537
rect 13455 13511 13481 13537
rect 18831 13511 18857 13537
rect 8751 13455 8777 13481
rect 10151 13455 10177 13481
rect 10599 13455 10625 13481
rect 10711 13455 10737 13481
rect 10767 13455 10793 13481
rect 13399 13455 13425 13481
rect 12447 13399 12473 13425
rect 9919 13315 9945 13341
rect 9971 13315 9997 13341
rect 10023 13315 10049 13341
rect 8751 13231 8777 13257
rect 9535 13231 9561 13257
rect 10207 13231 10233 13257
rect 10263 13231 10289 13257
rect 14239 13231 14265 13257
rect 9479 13175 9505 13201
rect 14407 13175 14433 13201
rect 2143 13119 2169 13145
rect 6959 13119 6985 13145
rect 9647 13119 9673 13145
rect 9759 13119 9785 13145
rect 10151 13119 10177 13145
rect 10319 13119 10345 13145
rect 10375 13119 10401 13145
rect 10655 13119 10681 13145
rect 12615 13119 12641 13145
rect 18831 13119 18857 13145
rect 7351 13063 7377 13089
rect 8415 13063 8441 13089
rect 11047 13063 11073 13089
rect 12111 13063 12137 13089
rect 12335 13063 12361 13089
rect 13007 13063 13033 13089
rect 14071 13063 14097 13089
rect 19951 13063 19977 13089
rect 967 13007 993 13033
rect 2239 12923 2265 12949
rect 2291 12923 2317 12949
rect 2343 12923 2369 12949
rect 17599 12923 17625 12949
rect 17651 12923 17677 12949
rect 17703 12923 17729 12949
rect 1023 12783 1049 12809
rect 12503 12783 12529 12809
rect 14127 12783 14153 12809
rect 20007 12783 20033 12809
rect 2143 12727 2169 12753
rect 10823 12727 10849 12753
rect 10935 12727 10961 12753
rect 11047 12727 11073 12753
rect 11327 12727 11353 12753
rect 11495 12727 11521 12753
rect 12447 12727 12473 12753
rect 12671 12727 12697 12753
rect 18831 12727 18857 12753
rect 7071 12671 7097 12697
rect 8135 12671 8161 12697
rect 8303 12671 8329 12697
rect 11215 12671 11241 12697
rect 12223 12671 12249 12697
rect 12279 12671 12305 12697
rect 13063 12671 13089 12697
rect 6959 12615 6985 12641
rect 7015 12615 7041 12641
rect 10991 12615 11017 12641
rect 11271 12615 11297 12641
rect 11943 12615 11969 12641
rect 12111 12615 12137 12641
rect 9919 12531 9945 12557
rect 9971 12531 9997 12557
rect 10023 12531 10049 12557
rect 7631 12447 7657 12473
rect 9423 12447 9449 12473
rect 12727 12447 12753 12473
rect 7015 12391 7041 12417
rect 7799 12391 7825 12417
rect 8807 12391 8833 12417
rect 8975 12391 9001 12417
rect 9367 12391 9393 12417
rect 10095 12391 10121 12417
rect 10655 12391 10681 12417
rect 12839 12391 12865 12417
rect 12895 12391 12921 12417
rect 12951 12391 12977 12417
rect 13623 12391 13649 12417
rect 13679 12391 13705 12417
rect 7407 12335 7433 12361
rect 8919 12335 8945 12361
rect 9031 12335 9057 12361
rect 9143 12335 9169 12361
rect 9647 12335 9673 12361
rect 9815 12335 9841 12361
rect 10823 12335 10849 12361
rect 5951 12279 5977 12305
rect 13119 12279 13145 12305
rect 7855 12223 7881 12249
rect 2239 12139 2265 12165
rect 2291 12139 2317 12165
rect 2343 12139 2369 12165
rect 17599 12139 17625 12165
rect 17651 12139 17677 12165
rect 17703 12139 17729 12165
rect 7183 12055 7209 12081
rect 10151 12055 10177 12081
rect 10711 12055 10737 12081
rect 12951 12055 12977 12081
rect 6735 11999 6761 12025
rect 6791 11943 6817 11969
rect 6903 11943 6929 11969
rect 7295 11943 7321 11969
rect 7687 11943 7713 11969
rect 7855 11943 7881 11969
rect 10151 11943 10177 11969
rect 11663 11943 11689 11969
rect 7071 11887 7097 11913
rect 7407 11887 7433 11913
rect 7575 11887 7601 11913
rect 9983 11887 10009 11913
rect 10655 11887 10681 11913
rect 11439 11887 11465 11913
rect 13007 11887 13033 11913
rect 7183 11831 7209 11857
rect 7631 11831 7657 11857
rect 10711 11831 10737 11857
rect 11271 11831 11297 11857
rect 11327 11831 11353 11857
rect 11383 11831 11409 11857
rect 12951 11831 12977 11857
rect 9919 11747 9945 11773
rect 9971 11747 9997 11773
rect 10023 11747 10049 11773
rect 7127 11663 7153 11689
rect 7407 11663 7433 11689
rect 8247 11663 8273 11689
rect 8695 11663 8721 11689
rect 6511 11607 6537 11633
rect 7631 11607 7657 11633
rect 8359 11607 8385 11633
rect 9199 11607 9225 11633
rect 10431 11607 10457 11633
rect 13735 11607 13761 11633
rect 6903 11551 6929 11577
rect 7351 11551 7377 11577
rect 7519 11551 7545 11577
rect 7855 11551 7881 11577
rect 8415 11551 8441 11577
rect 8863 11551 8889 11577
rect 9031 11551 9057 11577
rect 9535 11551 9561 11577
rect 13511 11551 13537 11577
rect 13623 11551 13649 11577
rect 18831 11551 18857 11577
rect 5447 11495 5473 11521
rect 13567 11495 13593 11521
rect 20007 11439 20033 11465
rect 2239 11355 2265 11381
rect 2291 11355 2317 11381
rect 2343 11355 2369 11381
rect 17599 11355 17625 11381
rect 17651 11355 17677 11381
rect 17703 11355 17729 11381
rect 5391 11215 5417 11241
rect 6455 11215 6481 11241
rect 6791 11215 6817 11241
rect 8807 11215 8833 11241
rect 9759 11215 9785 11241
rect 10095 11215 10121 11241
rect 11271 11215 11297 11241
rect 12335 11215 12361 11241
rect 12559 11215 12585 11241
rect 14295 11215 14321 11241
rect 20007 11215 20033 11241
rect 5055 11159 5081 11185
rect 7295 11159 7321 11185
rect 9087 11159 9113 11185
rect 9479 11159 9505 11185
rect 10935 11159 10961 11185
rect 12895 11159 12921 11185
rect 13231 11159 13257 11185
rect 18831 11159 18857 11185
rect 6959 11103 6985 11129
rect 7127 11103 7153 11129
rect 8975 11103 9001 11129
rect 9703 11103 9729 11129
rect 10263 11103 10289 11129
rect 7463 11047 7489 11073
rect 8527 11047 8553 11073
rect 9255 11047 9281 11073
rect 9815 11047 9841 11073
rect 10039 11047 10065 11073
rect 10151 11047 10177 11073
rect 9919 10963 9945 10989
rect 9971 10963 9997 10989
rect 10023 10963 10049 10989
rect 7519 10879 7545 10905
rect 8303 10879 8329 10905
rect 8919 10879 8945 10905
rect 9255 10879 9281 10905
rect 7071 10823 7097 10849
rect 8695 10823 8721 10849
rect 8751 10823 8777 10849
rect 10711 10851 10737 10877
rect 11999 10879 12025 10905
rect 12671 10879 12697 10905
rect 13343 10879 13369 10905
rect 9031 10823 9057 10849
rect 9423 10823 9449 10849
rect 9871 10823 9897 10849
rect 10375 10823 10401 10849
rect 11719 10823 11745 10849
rect 12055 10823 12081 10849
rect 12111 10823 12137 10849
rect 13455 10823 13481 10849
rect 13567 10823 13593 10849
rect 8023 10767 8049 10793
rect 8135 10767 8161 10793
rect 9087 10767 9113 10793
rect 9647 10767 9673 10793
rect 9703 10767 9729 10793
rect 10263 10767 10289 10793
rect 10655 10767 10681 10793
rect 10935 10767 10961 10793
rect 11215 10767 11241 10793
rect 11551 10767 11577 10793
rect 11943 10767 11969 10793
rect 12335 10767 12361 10793
rect 13287 10767 13313 10793
rect 18831 10767 18857 10793
rect 6567 10711 6593 10737
rect 7463 10711 7489 10737
rect 7631 10711 7657 10737
rect 11663 10711 11689 10737
rect 19951 10711 19977 10737
rect 7127 10655 7153 10681
rect 8751 10655 8777 10681
rect 9815 10655 9841 10681
rect 10711 10655 10737 10681
rect 2239 10571 2265 10597
rect 2291 10571 2317 10597
rect 2343 10571 2369 10597
rect 17599 10571 17625 10597
rect 17651 10571 17677 10597
rect 17703 10571 17729 10597
rect 7743 10487 7769 10513
rect 10823 10487 10849 10513
rect 5391 10431 5417 10457
rect 6455 10431 6481 10457
rect 6847 10431 6873 10457
rect 8247 10431 8273 10457
rect 10039 10431 10065 10457
rect 12671 10431 12697 10457
rect 14295 10431 14321 10457
rect 20007 10431 20033 10457
rect 5055 10375 5081 10401
rect 6903 10375 6929 10401
rect 7127 10375 7153 10401
rect 7407 10375 7433 10401
rect 7519 10375 7545 10401
rect 9031 10375 9057 10401
rect 9591 10375 9617 10401
rect 10095 10375 10121 10401
rect 10207 10375 10233 10401
rect 11047 10375 11073 10401
rect 11383 10375 11409 10401
rect 11831 10375 11857 10401
rect 11999 10375 12025 10401
rect 12839 10375 12865 10401
rect 14631 10375 14657 10401
rect 18831 10375 18857 10401
rect 7239 10319 7265 10345
rect 7967 10319 7993 10345
rect 9087 10319 9113 10345
rect 9983 10319 10009 10345
rect 10655 10319 10681 10345
rect 11215 10319 11241 10345
rect 11551 10319 11577 10345
rect 12111 10319 12137 10345
rect 13231 10319 13257 10345
rect 8863 10263 8889 10289
rect 9479 10263 9505 10289
rect 10767 10263 10793 10289
rect 12167 10263 12193 10289
rect 14743 10263 14769 10289
rect 9919 10179 9945 10205
rect 9971 10179 9997 10205
rect 10023 10179 10049 10205
rect 7463 10095 7489 10121
rect 12951 10095 12977 10121
rect 6735 10039 6761 10065
rect 7911 10039 7937 10065
rect 8863 10039 8889 10065
rect 10151 10039 10177 10065
rect 13567 10039 13593 10065
rect 13791 10039 13817 10065
rect 7743 9983 7769 10009
rect 8079 9983 8105 10009
rect 8695 9983 8721 10009
rect 9031 9983 9057 10009
rect 12895 9983 12921 10009
rect 13007 9983 13033 10009
rect 13231 9983 13257 10009
rect 13679 9983 13705 10009
rect 8135 9927 8161 9953
rect 11943 9927 11969 9953
rect 12783 9927 12809 9953
rect 13623 9927 13649 9953
rect 2239 9787 2265 9813
rect 2291 9787 2317 9813
rect 2343 9787 2369 9813
rect 17599 9787 17625 9813
rect 17651 9787 17677 9813
rect 17703 9787 17729 9813
rect 8135 9703 8161 9729
rect 9143 9703 9169 9729
rect 9759 9703 9785 9729
rect 9647 9647 9673 9673
rect 10263 9647 10289 9673
rect 11551 9647 11577 9673
rect 20007 9647 20033 9673
rect 7799 9591 7825 9617
rect 8303 9591 8329 9617
rect 8975 9591 9001 9617
rect 9199 9591 9225 9617
rect 9591 9591 9617 9617
rect 10095 9591 10121 9617
rect 10207 9591 10233 9617
rect 10711 9591 10737 9617
rect 11663 9591 11689 9617
rect 11943 9591 11969 9617
rect 12111 9591 12137 9617
rect 12895 9591 12921 9617
rect 13231 9591 13257 9617
rect 18831 9591 18857 9617
rect 7967 9535 7993 9561
rect 8415 9535 8441 9561
rect 8863 9535 8889 9561
rect 10935 9535 10961 9561
rect 11103 9535 11129 9561
rect 12391 9535 12417 9561
rect 13119 9535 13145 9561
rect 13567 9535 13593 9561
rect 13679 9535 13705 9561
rect 13735 9535 13761 9561
rect 9087 9479 9113 9505
rect 10319 9479 10345 9505
rect 10711 9479 10737 9505
rect 11719 9479 11745 9505
rect 11999 9479 12025 9505
rect 12559 9479 12585 9505
rect 13063 9479 13089 9505
rect 9919 9395 9945 9421
rect 9971 9395 9997 9421
rect 10023 9395 10049 9421
rect 9703 9311 9729 9337
rect 10543 9311 10569 9337
rect 10655 9311 10681 9337
rect 11047 9311 11073 9337
rect 11383 9311 11409 9337
rect 11495 9311 11521 9337
rect 7687 9255 7713 9281
rect 9255 9255 9281 9281
rect 13231 9255 13257 9281
rect 5895 9199 5921 9225
rect 6231 9199 6257 9225
rect 7855 9199 7881 9225
rect 7967 9199 7993 9225
rect 8135 9199 8161 9225
rect 8975 9199 9001 9225
rect 9871 9199 9897 9225
rect 10879 9199 10905 9225
rect 11215 9199 11241 9225
rect 11439 9199 11465 9225
rect 11719 9199 11745 9225
rect 12839 9199 12865 9225
rect 7295 9143 7321 9169
rect 7575 9143 7601 9169
rect 7743 9143 7769 9169
rect 8359 9143 8385 9169
rect 10599 9143 10625 9169
rect 12727 9143 12753 9169
rect 14295 9143 14321 9169
rect 2239 9003 2265 9029
rect 2291 9003 2317 9029
rect 2343 9003 2369 9029
rect 17599 9003 17625 9029
rect 17651 9003 17677 9029
rect 17703 9003 17729 9029
rect 10823 8919 10849 8945
rect 9647 8863 9673 8889
rect 10431 8863 10457 8889
rect 20007 8863 20033 8889
rect 7519 8807 7545 8833
rect 8415 8807 8441 8833
rect 8751 8807 8777 8833
rect 10375 8807 10401 8833
rect 11159 8807 11185 8833
rect 11663 8807 11689 8833
rect 13007 8807 13033 8833
rect 13231 8807 13257 8833
rect 13343 8807 13369 8833
rect 13567 8807 13593 8833
rect 13623 8807 13649 8833
rect 18831 8807 18857 8833
rect 7631 8751 7657 8777
rect 7967 8751 7993 8777
rect 8527 8751 8553 8777
rect 8863 8751 8889 8777
rect 9871 8751 9897 8777
rect 10095 8751 10121 8777
rect 10711 8751 10737 8777
rect 11327 8751 11353 8777
rect 8023 8695 8049 8721
rect 8079 8695 8105 8721
rect 9031 8695 9057 8721
rect 9199 8695 9225 8721
rect 9367 8695 9393 8721
rect 10991 8695 11017 8721
rect 11831 8695 11857 8721
rect 13175 8695 13201 8721
rect 13511 8695 13537 8721
rect 13735 8695 13761 8721
rect 9919 8611 9945 8637
rect 9971 8611 9997 8637
rect 10023 8611 10049 8637
rect 8359 8527 8385 8553
rect 8751 8527 8777 8553
rect 6455 8471 6481 8497
rect 8303 8471 8329 8497
rect 8695 8471 8721 8497
rect 9199 8471 9225 8497
rect 9255 8471 9281 8497
rect 10935 8471 10961 8497
rect 13231 8471 13257 8497
rect 6063 8415 6089 8441
rect 7743 8415 7769 8441
rect 9367 8415 9393 8441
rect 9479 8415 9505 8441
rect 12839 8415 12865 8441
rect 7519 8359 7545 8385
rect 12671 8359 12697 8385
rect 14295 8359 14321 8385
rect 2239 8219 2265 8245
rect 2291 8219 2317 8245
rect 2343 8219 2369 8245
rect 17599 8219 17625 8245
rect 17651 8219 17677 8245
rect 17703 8219 17729 8245
rect 8863 8135 8889 8161
rect 9479 8135 9505 8161
rect 20007 8079 20033 8105
rect 8751 8023 8777 8049
rect 8975 8023 9001 8049
rect 9143 8023 9169 8049
rect 9311 8023 9337 8049
rect 9423 8023 9449 8049
rect 10039 8023 10065 8049
rect 10263 8023 10289 8049
rect 10375 8023 10401 8049
rect 10655 8023 10681 8049
rect 10767 8023 10793 8049
rect 10991 8023 11017 8049
rect 13063 8023 13089 8049
rect 13287 8023 13313 8049
rect 13455 8023 13481 8049
rect 13623 8023 13649 8049
rect 18831 8023 18857 8049
rect 10151 7967 10177 7993
rect 12951 7967 12977 7993
rect 9087 7911 9113 7937
rect 9983 7911 10009 7937
rect 10823 7911 10849 7937
rect 10879 7911 10905 7937
rect 13175 7911 13201 7937
rect 13567 7911 13593 7937
rect 9919 7827 9945 7853
rect 9971 7827 9997 7853
rect 10023 7827 10049 7853
rect 8751 7743 8777 7769
rect 10207 7743 10233 7769
rect 10319 7743 10345 7769
rect 11887 7743 11913 7769
rect 10095 7687 10121 7713
rect 11831 7687 11857 7713
rect 11943 7687 11969 7713
rect 13175 7687 13201 7713
rect 7015 7631 7041 7657
rect 8975 7631 9001 7657
rect 9087 7631 9113 7657
rect 9703 7631 9729 7657
rect 9815 7631 9841 7657
rect 12335 7631 12361 7657
rect 12783 7631 12809 7657
rect 7351 7575 7377 7601
rect 8415 7575 8441 7601
rect 8919 7575 8945 7601
rect 9143 7575 9169 7601
rect 14239 7575 14265 7601
rect 9535 7519 9561 7545
rect 10151 7519 10177 7545
rect 2239 7435 2265 7461
rect 2291 7435 2317 7461
rect 2343 7435 2369 7461
rect 17599 7435 17625 7461
rect 17651 7435 17677 7461
rect 17703 7435 17729 7461
rect 10039 7351 10065 7377
rect 10151 7351 10177 7377
rect 12783 7351 12809 7377
rect 8863 7295 8889 7321
rect 9087 7295 9113 7321
rect 11159 7295 11185 7321
rect 12223 7295 12249 7321
rect 12447 7295 12473 7321
rect 7407 7239 7433 7265
rect 10263 7239 10289 7265
rect 10375 7239 10401 7265
rect 10823 7239 10849 7265
rect 7799 7183 7825 7209
rect 10319 7127 10345 7153
rect 12839 7127 12865 7153
rect 12895 7127 12921 7153
rect 9919 7043 9945 7069
rect 9971 7043 9997 7069
rect 10023 7043 10049 7069
rect 9143 6959 9169 6985
rect 11271 6959 11297 6985
rect 8303 6903 8329 6929
rect 8975 6903 9001 6929
rect 9927 6903 9953 6929
rect 10151 6903 10177 6929
rect 10207 6903 10233 6929
rect 12783 6903 12809 6929
rect 8415 6847 8441 6873
rect 9087 6847 9113 6873
rect 9311 6847 9337 6873
rect 9647 6847 9673 6873
rect 9759 6847 9785 6873
rect 10039 6847 10065 6873
rect 11215 6847 11241 6873
rect 11383 6847 11409 6873
rect 12615 6847 12641 6873
rect 8247 6791 8273 6817
rect 9871 6791 9897 6817
rect 12615 6735 12641 6761
rect 2239 6651 2265 6677
rect 2291 6651 2317 6677
rect 2343 6651 2369 6677
rect 17599 6651 17625 6677
rect 17651 6651 17677 6677
rect 17703 6651 17729 6677
rect 9031 6511 9057 6537
rect 10095 6511 10121 6537
rect 10319 6511 10345 6537
rect 11831 6511 11857 6537
rect 12391 6511 12417 6537
rect 13455 6511 13481 6537
rect 8695 6455 8721 6481
rect 10767 6455 10793 6481
rect 11999 6455 12025 6481
rect 10655 6343 10681 6369
rect 9919 6259 9945 6285
rect 9971 6259 9997 6285
rect 10023 6259 10049 6285
rect 11887 6175 11913 6201
rect 10599 6119 10625 6145
rect 10263 6063 10289 6089
rect 11663 6007 11689 6033
rect 2239 5867 2265 5893
rect 2291 5867 2317 5893
rect 2343 5867 2369 5893
rect 17599 5867 17625 5893
rect 17651 5867 17677 5893
rect 17703 5867 17729 5893
rect 9919 5475 9945 5501
rect 9971 5475 9997 5501
rect 10023 5475 10049 5501
rect 2239 5083 2265 5109
rect 2291 5083 2317 5109
rect 2343 5083 2369 5109
rect 17599 5083 17625 5109
rect 17651 5083 17677 5109
rect 17703 5083 17729 5109
rect 9919 4691 9945 4717
rect 9971 4691 9997 4717
rect 10023 4691 10049 4717
rect 2239 4299 2265 4325
rect 2291 4299 2317 4325
rect 2343 4299 2369 4325
rect 17599 4299 17625 4325
rect 17651 4299 17677 4325
rect 17703 4299 17729 4325
rect 9919 3907 9945 3933
rect 9971 3907 9997 3933
rect 10023 3907 10049 3933
rect 2239 3515 2265 3541
rect 2291 3515 2317 3541
rect 2343 3515 2369 3541
rect 17599 3515 17625 3541
rect 17651 3515 17677 3541
rect 17703 3515 17729 3541
rect 9919 3123 9945 3149
rect 9971 3123 9997 3149
rect 10023 3123 10049 3149
rect 2239 2731 2265 2757
rect 2291 2731 2317 2757
rect 2343 2731 2369 2757
rect 17599 2731 17625 2757
rect 17651 2731 17677 2757
rect 17703 2731 17729 2757
rect 9919 2339 9945 2365
rect 9971 2339 9997 2365
rect 10023 2339 10049 2365
rect 8863 2143 8889 2169
rect 12671 2143 12697 2169
rect 9367 2031 9393 2057
rect 13119 2031 13145 2057
rect 2239 1947 2265 1973
rect 2291 1947 2317 1973
rect 2343 1947 2369 1973
rect 17599 1947 17625 1973
rect 17651 1947 17677 1973
rect 17703 1947 17729 1973
rect 9311 1807 9337 1833
rect 12783 1807 12809 1833
rect 14687 1807 14713 1833
rect 9031 1751 9057 1777
rect 10375 1751 10401 1777
rect 12279 1751 12305 1777
rect 14295 1751 14321 1777
rect 3487 1639 3513 1665
rect 10879 1639 10905 1665
rect 9919 1555 9945 1581
rect 9971 1555 9997 1581
rect 10023 1555 10049 1581
<< metal2 >>
rect 8736 20600 8792 21000
rect 9744 20600 9800 21000
rect 10416 20600 10472 21000
rect 10752 20600 10808 21000
rect 11088 20600 11144 21000
rect 12096 20600 12152 21000
rect 2238 19222 2370 19227
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2238 19189 2370 19194
rect 8750 18746 8778 20600
rect 9590 19138 9618 19143
rect 9758 19138 9786 20600
rect 9590 19137 9786 19138
rect 9590 19111 9591 19137
rect 9617 19111 9786 19137
rect 9590 19110 9786 19111
rect 9590 19105 9618 19110
rect 9870 19026 9898 19031
rect 9702 19025 9898 19026
rect 9702 18999 9871 19025
rect 9897 18999 9898 19025
rect 9702 18998 9898 18999
rect 8750 18713 8778 18718
rect 9366 18746 9394 18751
rect 9366 18699 9394 18718
rect 8862 18633 8890 18639
rect 8862 18607 8863 18633
rect 8889 18607 8890 18633
rect 2238 18438 2370 18443
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2238 18405 2370 18410
rect 2238 17654 2370 17659
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2238 17621 2370 17626
rect 2238 16870 2370 16875
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2238 16837 2370 16842
rect 2238 16086 2370 16091
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2238 16053 2370 16058
rect 8862 15974 8890 18607
rect 8414 15946 8890 15974
rect 2238 15302 2370 15307
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2238 15269 2370 15274
rect 2238 14518 2370 14523
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2238 14485 2370 14490
rect 2086 13818 2114 13823
rect 966 13033 994 13039
rect 966 13007 967 13033
rect 993 13007 994 13033
rect 966 12810 994 13007
rect 966 12777 994 12782
rect 1022 12809 1050 12815
rect 1022 12783 1023 12809
rect 1049 12783 1050 12809
rect 1022 12474 1050 12783
rect 1022 12441 1050 12446
rect 2086 10290 2114 13790
rect 2238 13734 2370 13739
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2238 13701 2370 13706
rect 8414 13650 8442 15946
rect 9422 13930 9450 13935
rect 9422 13883 9450 13902
rect 9702 13762 9730 18998
rect 9870 18993 9898 18998
rect 9918 18830 10050 18835
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 9918 18797 10050 18802
rect 10430 18746 10458 20600
rect 10766 19138 10794 20600
rect 10766 19105 10794 19110
rect 10710 19025 10738 19031
rect 10710 18999 10711 19025
rect 10737 18999 10738 19025
rect 10542 18970 10570 18975
rect 10542 18923 10570 18942
rect 10430 18713 10458 18718
rect 9918 18046 10050 18051
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 9918 18013 10050 18018
rect 9918 17262 10050 17267
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 9918 17229 10050 17234
rect 9918 16478 10050 16483
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 9918 16445 10050 16450
rect 9918 15694 10050 15699
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 9918 15661 10050 15666
rect 9918 14910 10050 14915
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 9918 14877 10050 14882
rect 9918 14126 10050 14131
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 9918 14093 10050 14098
rect 10318 14042 10346 14047
rect 9758 13874 9786 13879
rect 9758 13873 10010 13874
rect 9758 13847 9759 13873
rect 9785 13847 10010 13873
rect 9758 13846 10010 13847
rect 9758 13841 9786 13846
rect 9702 13734 9842 13762
rect 8358 13622 8442 13650
rect 8358 13454 8386 13622
rect 9814 13594 9842 13734
rect 9982 13649 10010 13846
rect 9982 13623 9983 13649
rect 10009 13623 10010 13649
rect 9982 13617 10010 13623
rect 9814 13547 9842 13566
rect 8414 13538 8442 13543
rect 8414 13537 8498 13538
rect 8414 13511 8415 13537
rect 8441 13511 8498 13537
rect 8414 13510 8498 13511
rect 8414 13505 8442 13510
rect 8470 13454 8498 13510
rect 9982 13537 10010 13543
rect 9982 13511 9983 13537
rect 10009 13511 10010 13537
rect 8750 13481 8778 13487
rect 8750 13455 8751 13481
rect 8777 13455 8778 13481
rect 8358 13426 8442 13454
rect 2142 13146 2170 13151
rect 2142 13099 2170 13118
rect 5950 13146 5978 13151
rect 6958 13146 6986 13151
rect 2238 12950 2370 12955
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2238 12917 2370 12922
rect 2142 12754 2170 12759
rect 2142 12707 2170 12726
rect 5446 12754 5474 12759
rect 2238 12166 2370 12171
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2238 12133 2370 12138
rect 5446 12026 5474 12726
rect 5950 12418 5978 13118
rect 5950 12305 5978 12390
rect 5950 12279 5951 12305
rect 5977 12279 5978 12305
rect 5950 12273 5978 12279
rect 6902 13145 6986 13146
rect 6902 13119 6959 13145
rect 6985 13119 6986 13145
rect 6902 13118 6986 13119
rect 6902 12306 6930 13118
rect 6958 13113 6986 13118
rect 7350 13090 7378 13095
rect 7350 13043 7378 13062
rect 8134 13090 8162 13095
rect 7070 12698 7098 12703
rect 7070 12697 7378 12698
rect 7070 12671 7071 12697
rect 7097 12671 7378 12697
rect 7070 12670 7378 12671
rect 7070 12665 7098 12670
rect 6902 12273 6930 12278
rect 6958 12641 6986 12647
rect 6958 12615 6959 12641
rect 6985 12615 6986 12641
rect 6958 12082 6986 12615
rect 7014 12641 7042 12647
rect 7014 12615 7015 12641
rect 7041 12615 7042 12641
rect 7014 12417 7042 12615
rect 7014 12391 7015 12417
rect 7041 12391 7042 12417
rect 7014 12385 7042 12391
rect 6958 12049 6986 12054
rect 7126 12306 7154 12311
rect 5446 11521 5474 11998
rect 6734 12026 6762 12031
rect 6734 11979 6762 11998
rect 6790 11970 6818 11975
rect 6902 11970 6930 11975
rect 6790 11969 6930 11970
rect 6790 11943 6791 11969
rect 6817 11943 6903 11969
rect 6929 11943 6930 11969
rect 6790 11942 6930 11943
rect 6790 11937 6818 11942
rect 6902 11937 6930 11942
rect 7070 11914 7098 11919
rect 7070 11867 7098 11886
rect 6510 11858 6538 11863
rect 6510 11633 6538 11830
rect 7126 11690 7154 12278
rect 7182 12082 7210 12087
rect 7182 12035 7210 12054
rect 7294 11969 7322 11975
rect 7294 11943 7295 11969
rect 7321 11943 7322 11969
rect 7182 11858 7210 11863
rect 7182 11811 7210 11830
rect 7294 11802 7322 11943
rect 7294 11769 7322 11774
rect 6510 11607 6511 11633
rect 6537 11607 6538 11633
rect 6510 11601 6538 11607
rect 6902 11689 7154 11690
rect 6902 11663 7127 11689
rect 7153 11663 7154 11689
rect 6902 11662 7154 11663
rect 7350 11690 7378 12670
rect 8134 12697 8162 13062
rect 8414 13089 8442 13426
rect 8414 13063 8415 13089
rect 8441 13063 8442 13089
rect 8134 12671 8135 12697
rect 8161 12671 8162 12697
rect 8134 12665 8162 12671
rect 8302 12697 8330 12703
rect 8302 12671 8303 12697
rect 8329 12671 8330 12697
rect 7630 12586 7658 12591
rect 7630 12473 7658 12558
rect 8302 12530 8330 12671
rect 8302 12497 8330 12502
rect 7630 12447 7631 12473
rect 7657 12447 7658 12473
rect 7406 12361 7434 12367
rect 7406 12335 7407 12361
rect 7433 12335 7434 12361
rect 7406 12306 7434 12335
rect 7406 12273 7434 12278
rect 7630 12306 7658 12447
rect 7798 12418 7826 12423
rect 8414 12418 8442 13063
rect 8470 13426 8722 13454
rect 8470 12586 8498 13426
rect 8694 13258 8722 13426
rect 8750 13370 8778 13455
rect 8750 13337 8778 13342
rect 9478 13482 9506 13487
rect 9982 13454 10010 13511
rect 8750 13258 8778 13263
rect 8694 13257 8778 13258
rect 8694 13231 8751 13257
rect 8777 13231 8778 13257
rect 8694 13230 8778 13231
rect 8750 13225 8778 13230
rect 9478 13201 9506 13454
rect 9758 13426 10010 13454
rect 10150 13482 10178 13487
rect 10318 13482 10346 14014
rect 10710 13986 10738 18999
rect 11102 18970 11130 20600
rect 11214 19138 11242 19143
rect 11214 19091 11242 19110
rect 12110 19138 12138 20600
rect 17598 19222 17730 19227
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17598 19189 17730 19194
rect 12110 19105 12138 19110
rect 12782 19138 12810 19143
rect 12782 19091 12810 19110
rect 11102 18937 11130 18942
rect 12278 19025 12306 19031
rect 12278 18999 12279 19025
rect 12305 18999 12306 19025
rect 11046 18746 11074 18751
rect 11046 18699 11074 18718
rect 10766 18634 10794 18639
rect 10766 18633 10850 18634
rect 10766 18607 10767 18633
rect 10793 18607 10850 18633
rect 10766 18606 10850 18607
rect 10766 18601 10794 18606
rect 10710 13953 10738 13958
rect 10822 14042 10850 18606
rect 12278 15974 12306 18999
rect 17598 18438 17730 18443
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17598 18405 17730 18410
rect 17598 17654 17730 17659
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17598 17621 17730 17626
rect 20118 17345 20146 17351
rect 20118 17319 20119 17345
rect 20145 17319 20146 17345
rect 20118 17178 20146 17319
rect 20118 17145 20146 17150
rect 17598 16870 17730 16875
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17598 16837 17730 16842
rect 17598 16086 17730 16091
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17598 16053 17730 16058
rect 12054 15946 12306 15974
rect 10374 13874 10402 13879
rect 10374 13594 10402 13846
rect 10822 13873 10850 14014
rect 11158 14042 11186 14047
rect 11158 13995 11186 14014
rect 10990 13986 11018 13991
rect 10990 13939 11018 13958
rect 10822 13847 10823 13873
rect 10849 13847 10850 13873
rect 10822 13841 10850 13847
rect 11438 13874 11466 13879
rect 11438 13827 11466 13846
rect 11942 13874 11970 13879
rect 10710 13594 10738 13599
rect 10374 13593 10682 13594
rect 10374 13567 10375 13593
rect 10401 13567 10682 13593
rect 10374 13566 10682 13567
rect 10374 13561 10402 13566
rect 10598 13482 10626 13487
rect 10150 13481 10290 13482
rect 10150 13455 10151 13481
rect 10177 13455 10290 13481
rect 10150 13454 10290 13455
rect 10318 13454 10402 13482
rect 10150 13449 10178 13454
rect 9534 13370 9562 13375
rect 9534 13257 9562 13342
rect 9534 13231 9535 13257
rect 9561 13231 9562 13257
rect 9534 13225 9562 13231
rect 9478 13175 9479 13201
rect 9505 13175 9506 13201
rect 9478 13169 9506 13175
rect 9646 13146 9674 13151
rect 9646 13145 9730 13146
rect 9646 13119 9647 13145
rect 9673 13119 9730 13145
rect 9646 13118 9730 13119
rect 9646 13113 9674 13118
rect 8470 12553 8498 12558
rect 9086 12586 9114 12591
rect 8806 12418 8834 12423
rect 8414 12417 8834 12418
rect 8414 12391 8807 12417
rect 8833 12391 8834 12417
rect 8414 12390 8834 12391
rect 7798 12371 7826 12390
rect 8806 12385 8834 12390
rect 8974 12418 9002 12423
rect 8974 12371 9002 12390
rect 7630 12273 7658 12278
rect 8246 12362 8274 12367
rect 7854 12249 7882 12255
rect 7854 12223 7855 12249
rect 7881 12223 7882 12249
rect 7686 11969 7714 11975
rect 7686 11943 7687 11969
rect 7713 11943 7714 11969
rect 7406 11914 7434 11919
rect 7406 11913 7490 11914
rect 7406 11887 7407 11913
rect 7433 11887 7490 11913
rect 7406 11886 7490 11887
rect 7406 11881 7434 11886
rect 7406 11690 7434 11695
rect 7350 11689 7434 11690
rect 7350 11663 7407 11689
rect 7433 11663 7434 11689
rect 7350 11662 7434 11663
rect 6902 11578 6930 11662
rect 7126 11657 7154 11662
rect 7406 11657 7434 11662
rect 5446 11495 5447 11521
rect 5473 11495 5474 11521
rect 5446 11489 5474 11495
rect 6790 11577 6930 11578
rect 6790 11551 6903 11577
rect 6929 11551 6930 11577
rect 6790 11550 6930 11551
rect 2238 11382 2370 11387
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2238 11349 2370 11354
rect 5390 11354 5418 11359
rect 5390 11241 5418 11326
rect 5390 11215 5391 11241
rect 5417 11215 5418 11241
rect 5390 11209 5418 11215
rect 6454 11242 6482 11247
rect 6454 11195 6482 11214
rect 6790 11241 6818 11550
rect 6902 11545 6930 11550
rect 7350 11577 7378 11583
rect 7350 11551 7351 11577
rect 7377 11551 7378 11577
rect 6790 11215 6791 11241
rect 6817 11215 6818 11241
rect 5054 11185 5082 11191
rect 5054 11159 5055 11185
rect 5081 11159 5082 11185
rect 5054 10962 5082 11159
rect 2238 10598 2370 10603
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2238 10565 2370 10570
rect 5054 10401 5082 10934
rect 6790 10962 6818 11215
rect 6958 11354 6986 11359
rect 6958 11129 6986 11326
rect 6958 11103 6959 11129
rect 6985 11103 6986 11129
rect 6958 11097 6986 11103
rect 7070 11242 7098 11247
rect 6566 10737 6594 10743
rect 6566 10711 6567 10737
rect 6593 10711 6594 10737
rect 5390 10626 5418 10631
rect 5390 10457 5418 10598
rect 6566 10626 6594 10711
rect 6566 10593 6594 10598
rect 5390 10431 5391 10457
rect 5417 10431 5418 10457
rect 5390 10425 5418 10431
rect 6454 10458 6482 10463
rect 6454 10411 6482 10430
rect 5054 10375 5055 10401
rect 5081 10375 5082 10401
rect 5054 10369 5082 10375
rect 2086 10257 2114 10262
rect 6734 10066 6762 10071
rect 6790 10066 6818 10934
rect 7070 10849 7098 11214
rect 7294 11242 7322 11247
rect 7294 11185 7322 11214
rect 7294 11159 7295 11185
rect 7321 11159 7322 11185
rect 7294 11153 7322 11159
rect 7126 11130 7154 11135
rect 7350 11130 7378 11551
rect 7462 11354 7490 11886
rect 7574 11913 7602 11919
rect 7574 11887 7575 11913
rect 7601 11887 7602 11913
rect 7574 11802 7602 11887
rect 7574 11769 7602 11774
rect 7630 11857 7658 11863
rect 7630 11831 7631 11857
rect 7657 11831 7658 11857
rect 7630 11633 7658 11831
rect 7630 11607 7631 11633
rect 7657 11607 7658 11633
rect 7630 11601 7658 11607
rect 7518 11578 7546 11583
rect 7518 11531 7546 11550
rect 7574 11578 7602 11583
rect 7462 11321 7490 11326
rect 7126 11129 7266 11130
rect 7126 11103 7127 11129
rect 7153 11103 7266 11129
rect 7126 11102 7266 11103
rect 7126 11097 7154 11102
rect 7238 10962 7266 11102
rect 7350 11097 7378 11102
rect 7462 11074 7490 11079
rect 7462 11027 7490 11046
rect 7238 10934 7490 10962
rect 7070 10823 7071 10849
rect 7097 10823 7098 10849
rect 7070 10817 7098 10823
rect 7462 10737 7490 10934
rect 7518 10906 7546 10911
rect 7518 10859 7546 10878
rect 7462 10711 7463 10737
rect 7489 10711 7490 10737
rect 7462 10705 7490 10711
rect 7126 10682 7154 10687
rect 7126 10681 7434 10682
rect 7126 10655 7127 10681
rect 7153 10655 7434 10681
rect 7126 10654 7434 10655
rect 7126 10649 7154 10654
rect 7238 10570 7266 10575
rect 6846 10458 6874 10463
rect 6846 10411 6874 10430
rect 7126 10458 7154 10463
rect 6902 10402 6930 10407
rect 6902 10355 6930 10374
rect 7126 10401 7154 10430
rect 7126 10375 7127 10401
rect 7153 10375 7154 10401
rect 7126 10369 7154 10375
rect 7238 10345 7266 10542
rect 7238 10319 7239 10345
rect 7265 10319 7266 10345
rect 7238 10313 7266 10319
rect 7406 10401 7434 10654
rect 7574 10626 7602 11550
rect 7630 10738 7658 10743
rect 7630 10691 7658 10710
rect 7574 10593 7602 10598
rect 7686 10514 7714 11943
rect 7854 11969 7882 12223
rect 7854 11943 7855 11969
rect 7881 11943 7882 11969
rect 7854 11937 7882 11943
rect 8246 11914 8274 12334
rect 8918 12362 8946 12367
rect 8918 12315 8946 12334
rect 9030 12361 9058 12367
rect 9030 12335 9031 12361
rect 9057 12335 9058 12361
rect 9030 11970 9058 12335
rect 8246 11689 8274 11886
rect 8246 11663 8247 11689
rect 8273 11663 8274 11689
rect 8246 11657 8274 11663
rect 8694 11942 9058 11970
rect 8694 11802 8722 11942
rect 9086 11914 9114 12558
rect 9422 12530 9450 12535
rect 9422 12473 9450 12502
rect 9422 12447 9423 12473
rect 9449 12447 9450 12473
rect 9422 12441 9450 12447
rect 9366 12418 9394 12423
rect 9366 12371 9394 12390
rect 9142 12362 9170 12367
rect 9142 12315 9170 12334
rect 9646 12361 9674 12367
rect 9646 12335 9647 12361
rect 9673 12335 9674 12361
rect 9086 11881 9114 11886
rect 8694 11689 8722 11774
rect 8694 11663 8695 11689
rect 8721 11663 8722 11689
rect 8358 11633 8386 11639
rect 8358 11607 8359 11633
rect 8385 11607 8386 11633
rect 7854 11578 7882 11583
rect 7854 11531 7882 11550
rect 7910 11130 7938 11135
rect 7910 11018 7938 11102
rect 7686 10481 7714 10486
rect 7742 10906 7770 10911
rect 7742 10514 7770 10878
rect 7742 10513 7882 10514
rect 7742 10487 7743 10513
rect 7769 10487 7882 10513
rect 7742 10486 7882 10487
rect 7742 10481 7770 10486
rect 7406 10375 7407 10401
rect 7433 10375 7434 10401
rect 7406 10346 7434 10375
rect 7406 10122 7434 10318
rect 7518 10402 7546 10407
rect 7462 10122 7490 10127
rect 7406 10121 7490 10122
rect 7406 10095 7463 10121
rect 7489 10095 7490 10121
rect 7406 10094 7490 10095
rect 7462 10089 7490 10094
rect 7518 10094 7546 10374
rect 7854 10122 7882 10486
rect 7518 10066 7826 10094
rect 6734 10065 6818 10066
rect 6734 10039 6735 10065
rect 6761 10039 6818 10065
rect 6734 10038 6818 10039
rect 6734 10033 6762 10038
rect 7742 10010 7770 10015
rect 7742 9963 7770 9982
rect 2238 9814 2370 9819
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2238 9781 2370 9786
rect 7798 9617 7826 10066
rect 7854 9842 7882 10094
rect 7910 10065 7938 10990
rect 8022 11074 8050 11079
rect 8022 10793 8050 11046
rect 8302 10906 8330 10911
rect 8358 10906 8386 11607
rect 8302 10905 8386 10906
rect 8302 10879 8303 10905
rect 8329 10879 8386 10905
rect 8302 10878 8386 10879
rect 8414 11578 8442 11583
rect 8022 10767 8023 10793
rect 8049 10767 8050 10793
rect 8022 10761 8050 10767
rect 8134 10793 8162 10799
rect 8134 10767 8135 10793
rect 8161 10767 8162 10793
rect 8134 10570 8162 10767
rect 8134 10537 8162 10542
rect 8302 10738 8330 10878
rect 8246 10514 8274 10519
rect 8246 10457 8274 10486
rect 8246 10431 8247 10457
rect 8273 10431 8274 10457
rect 8246 10425 8274 10431
rect 7966 10346 7994 10351
rect 7966 10299 7994 10318
rect 7910 10039 7911 10065
rect 7937 10039 7938 10065
rect 7910 10033 7938 10039
rect 8078 10010 8106 10015
rect 8078 9963 8106 9982
rect 7966 9954 7994 9959
rect 7854 9814 7938 9842
rect 7798 9591 7799 9617
rect 7825 9591 7826 9617
rect 7798 9585 7826 9591
rect 7742 9562 7770 9567
rect 7686 9534 7742 9562
rect 7630 9506 7658 9511
rect 5894 9226 5922 9231
rect 6230 9226 6258 9231
rect 5894 9225 6090 9226
rect 5894 9199 5895 9225
rect 5921 9199 6090 9225
rect 5894 9198 6090 9199
rect 5894 9193 5922 9198
rect 6062 9170 6090 9198
rect 6230 9179 6258 9198
rect 2238 9030 2370 9035
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2238 8997 2370 9002
rect 6062 8441 6090 9142
rect 7014 9170 7042 9175
rect 6454 8778 6482 8783
rect 6454 8497 6482 8750
rect 6454 8471 6455 8497
rect 6481 8471 6482 8497
rect 6454 8465 6482 8471
rect 6062 8415 6063 8441
rect 6089 8415 6090 8441
rect 6062 8409 6090 8415
rect 2238 8246 2370 8251
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2238 8213 2370 8218
rect 7014 7658 7042 9142
rect 7294 9169 7322 9175
rect 7294 9143 7295 9169
rect 7321 9143 7322 9169
rect 7294 8834 7322 9143
rect 7574 9170 7602 9175
rect 7518 8834 7546 8839
rect 7294 8833 7546 8834
rect 7294 8807 7519 8833
rect 7545 8807 7546 8833
rect 7294 8806 7546 8807
rect 7518 8666 7546 8806
rect 7518 8633 7546 8638
rect 7518 8498 7546 8503
rect 7518 8385 7546 8470
rect 7574 8442 7602 9142
rect 7630 8777 7658 9478
rect 7686 9281 7714 9534
rect 7742 9529 7770 9534
rect 7686 9255 7687 9281
rect 7713 9255 7714 9281
rect 7686 9249 7714 9255
rect 7854 9226 7882 9231
rect 7910 9226 7938 9814
rect 7966 9561 7994 9926
rect 7966 9535 7967 9561
rect 7993 9535 7994 9561
rect 7966 9529 7994 9535
rect 8134 9953 8162 9959
rect 8134 9927 8135 9953
rect 8161 9927 8162 9953
rect 8134 9729 8162 9927
rect 8134 9703 8135 9729
rect 8161 9703 8162 9729
rect 8134 9562 8162 9703
rect 8134 9529 8162 9534
rect 8190 9786 8218 9791
rect 7854 9225 7938 9226
rect 7854 9199 7855 9225
rect 7881 9199 7938 9225
rect 7854 9198 7938 9199
rect 7966 9225 7994 9231
rect 7966 9199 7967 9225
rect 7993 9199 7994 9225
rect 7854 9193 7882 9198
rect 7630 8751 7631 8777
rect 7657 8751 7658 8777
rect 7630 8745 7658 8751
rect 7742 9169 7770 9175
rect 7742 9143 7743 9169
rect 7769 9143 7770 9169
rect 7742 8778 7770 9143
rect 7966 9058 7994 9199
rect 7966 9025 7994 9030
rect 8134 9225 8162 9231
rect 8134 9199 8135 9225
rect 8161 9199 8162 9225
rect 8134 8834 8162 9199
rect 7742 8745 7770 8750
rect 7966 8806 8162 8834
rect 7966 8777 7994 8806
rect 7966 8751 7967 8777
rect 7993 8751 7994 8777
rect 7966 8498 7994 8751
rect 8022 8721 8050 8727
rect 8022 8695 8023 8721
rect 8049 8695 8050 8721
rect 8022 8554 8050 8695
rect 8078 8721 8106 8727
rect 8078 8695 8079 8721
rect 8105 8695 8106 8721
rect 8078 8666 8106 8695
rect 8078 8633 8106 8638
rect 8190 8554 8218 9758
rect 8302 9730 8330 10710
rect 8414 9786 8442 11550
rect 8526 11074 8554 11079
rect 8526 11027 8554 11046
rect 8694 10849 8722 11663
rect 8806 11858 8834 11863
rect 8806 11242 8834 11830
rect 9590 11690 9618 11695
rect 9198 11634 9226 11639
rect 9198 11633 9506 11634
rect 9198 11607 9199 11633
rect 9225 11607 9506 11633
rect 9198 11606 9506 11607
rect 9198 11601 9226 11606
rect 8862 11578 8890 11583
rect 8862 11531 8890 11550
rect 9030 11577 9058 11583
rect 9030 11551 9031 11577
rect 9057 11551 9058 11577
rect 8806 11241 8890 11242
rect 8806 11215 8807 11241
rect 8833 11215 8890 11241
rect 8806 11214 8890 11215
rect 8806 11209 8834 11214
rect 8694 10823 8695 10849
rect 8721 10823 8722 10849
rect 8694 10817 8722 10823
rect 8750 10850 8778 10855
rect 8750 10849 8834 10850
rect 8750 10823 8751 10849
rect 8777 10823 8834 10849
rect 8750 10822 8834 10823
rect 8750 10817 8778 10822
rect 8414 9753 8442 9758
rect 8470 10738 8498 10743
rect 8302 9697 8330 9702
rect 8302 9617 8330 9623
rect 8302 9591 8303 9617
rect 8329 9591 8330 9617
rect 8302 9562 8330 9591
rect 8302 9529 8330 9534
rect 8414 9562 8442 9567
rect 8470 9562 8498 10710
rect 8750 10681 8778 10687
rect 8750 10655 8751 10681
rect 8777 10655 8778 10681
rect 8582 10514 8610 10519
rect 8414 9561 8498 9562
rect 8414 9535 8415 9561
rect 8441 9535 8498 9561
rect 8414 9534 8498 9535
rect 8526 9618 8554 9623
rect 8414 9506 8442 9534
rect 8414 9473 8442 9478
rect 8414 9282 8442 9287
rect 8358 9254 8414 9282
rect 8358 9169 8386 9254
rect 8414 9249 8442 9254
rect 8358 9143 8359 9169
rect 8385 9143 8386 9169
rect 8358 9137 8386 9143
rect 8414 8833 8442 8839
rect 8414 8807 8415 8833
rect 8441 8807 8442 8833
rect 8414 8722 8442 8807
rect 8414 8689 8442 8694
rect 8526 8777 8554 9590
rect 8582 9114 8610 10486
rect 8750 10402 8778 10655
rect 8806 10682 8834 10822
rect 8806 10649 8834 10654
rect 8862 10458 8890 11214
rect 8918 11130 8946 11135
rect 8918 10905 8946 11102
rect 8918 10879 8919 10905
rect 8945 10879 8946 10905
rect 8918 10873 8946 10879
rect 8974 11130 9002 11135
rect 9030 11130 9058 11551
rect 8974 11129 9058 11130
rect 8974 11103 8975 11129
rect 9001 11103 9058 11129
rect 8974 11102 9058 11103
rect 9086 11185 9114 11191
rect 9086 11159 9087 11185
rect 9113 11159 9114 11185
rect 8974 10570 9002 11102
rect 9086 11074 9114 11159
rect 9478 11186 9506 11606
rect 9478 11153 9506 11158
rect 9534 11577 9562 11583
rect 9534 11551 9535 11577
rect 9561 11551 9562 11577
rect 9254 11074 9282 11079
rect 9114 11046 9226 11074
rect 9086 11041 9114 11046
rect 9198 10906 9226 11046
rect 9254 11027 9282 11046
rect 9478 11074 9506 11079
rect 9254 10906 9282 10911
rect 9198 10905 9282 10906
rect 9198 10879 9255 10905
rect 9281 10879 9282 10905
rect 9198 10878 9282 10879
rect 9254 10873 9282 10878
rect 9030 10849 9058 10855
rect 9030 10823 9031 10849
rect 9057 10823 9058 10849
rect 9030 10738 9058 10823
rect 9422 10849 9450 10855
rect 9422 10823 9423 10849
rect 9449 10823 9450 10849
rect 9086 10794 9114 10799
rect 9086 10793 9226 10794
rect 9086 10767 9087 10793
rect 9113 10767 9226 10793
rect 9086 10766 9226 10767
rect 9086 10761 9114 10766
rect 9030 10682 9058 10710
rect 9030 10654 9170 10682
rect 9030 10570 9058 10575
rect 8974 10542 9030 10570
rect 9058 10542 9114 10570
rect 9030 10537 9058 10542
rect 8750 10369 8778 10374
rect 8806 10430 9058 10458
rect 8806 10094 8834 10430
rect 9030 10401 9058 10430
rect 9030 10375 9031 10401
rect 9057 10375 9058 10401
rect 9030 10369 9058 10375
rect 9086 10345 9114 10542
rect 9142 10458 9170 10654
rect 9142 10425 9170 10430
rect 9086 10319 9087 10345
rect 9113 10319 9114 10345
rect 9086 10313 9114 10319
rect 9142 10346 9170 10351
rect 8862 10290 8890 10295
rect 8890 10262 8946 10290
rect 8862 10243 8890 10262
rect 8638 10066 8834 10094
rect 8638 9170 8666 10066
rect 8862 10065 8890 10071
rect 8862 10039 8863 10065
rect 8889 10039 8890 10065
rect 8694 10009 8722 10015
rect 8694 9983 8695 10009
rect 8721 9983 8722 10009
rect 8694 9282 8722 9983
rect 8806 10010 8834 10015
rect 8806 9506 8834 9982
rect 8862 9562 8890 10039
rect 8918 10010 8946 10262
rect 9030 10010 9058 10015
rect 8918 10009 9058 10010
rect 8918 9983 9031 10009
rect 9057 9983 9058 10009
rect 8918 9982 9058 9983
rect 9030 9977 9058 9982
rect 9142 9729 9170 10318
rect 9142 9703 9143 9729
rect 9169 9703 9170 9729
rect 9142 9697 9170 9703
rect 9198 9730 9226 10766
rect 9422 10682 9450 10823
rect 9422 10649 9450 10654
rect 9478 10289 9506 11046
rect 9478 10263 9479 10289
rect 9505 10263 9506 10289
rect 9478 10178 9506 10263
rect 9366 10150 9506 10178
rect 9198 9702 9282 9730
rect 8974 9618 9002 9623
rect 9198 9618 9226 9623
rect 9002 9617 9226 9618
rect 9002 9591 9199 9617
rect 9225 9591 9226 9617
rect 9002 9590 9226 9591
rect 8974 9571 9002 9590
rect 9198 9585 9226 9590
rect 8862 9515 8890 9534
rect 8806 9473 8834 9478
rect 9086 9506 9114 9511
rect 9254 9506 9282 9702
rect 9086 9459 9114 9478
rect 9142 9478 9282 9506
rect 9310 9618 9338 9623
rect 8694 9249 8722 9254
rect 8974 9226 9002 9231
rect 8638 9137 8666 9142
rect 8750 9225 9002 9226
rect 8750 9199 8975 9225
rect 9001 9199 9002 9225
rect 8750 9198 9002 9199
rect 8582 9081 8610 9086
rect 8526 8751 8527 8777
rect 8553 8751 8554 8777
rect 8022 8526 8218 8554
rect 8358 8554 8386 8559
rect 8358 8507 8386 8526
rect 7966 8465 7994 8470
rect 8302 8498 8330 8503
rect 8302 8451 8330 8470
rect 7742 8442 7770 8447
rect 7574 8414 7742 8442
rect 7742 8395 7770 8414
rect 7518 8359 7519 8385
rect 7545 8359 7546 8385
rect 7518 8353 7546 8359
rect 8526 8162 8554 8751
rect 8750 8833 8778 9198
rect 8974 9193 9002 9198
rect 8862 9114 8890 9119
rect 9142 9114 9170 9478
rect 9254 9282 9282 9287
rect 9254 9235 9282 9254
rect 8890 9086 9002 9114
rect 8862 9081 8890 9086
rect 8750 8807 8751 8833
rect 8777 8807 8778 8833
rect 8750 8722 8778 8807
rect 8862 8778 8890 8783
rect 8862 8731 8890 8750
rect 8582 8666 8610 8671
rect 8610 8638 8666 8666
rect 8582 8633 8610 8638
rect 8638 8498 8666 8638
rect 8750 8553 8778 8694
rect 8750 8527 8751 8553
rect 8777 8527 8778 8553
rect 8750 8521 8778 8527
rect 8694 8498 8722 8503
rect 8638 8497 8722 8498
rect 8638 8471 8695 8497
rect 8721 8471 8722 8497
rect 8638 8470 8722 8471
rect 8694 8465 8722 8470
rect 8918 8386 8946 8391
rect 8526 8129 8554 8134
rect 8862 8162 8890 8167
rect 8862 8115 8890 8134
rect 8750 8050 8778 8055
rect 8526 8049 8778 8050
rect 8526 8023 8751 8049
rect 8777 8023 8778 8049
rect 8526 8022 8778 8023
rect 7014 7657 7322 7658
rect 7014 7631 7015 7657
rect 7041 7631 7322 7657
rect 7014 7630 7322 7631
rect 7014 7625 7042 7630
rect 7294 7490 7322 7630
rect 7350 7602 7378 7607
rect 7350 7555 7378 7574
rect 8414 7602 8442 7607
rect 8414 7601 8498 7602
rect 8414 7575 8415 7601
rect 8441 7575 8498 7601
rect 8414 7574 8498 7575
rect 8526 7574 8554 8022
rect 8750 8017 8778 8022
rect 8750 7770 8778 7775
rect 8918 7770 8946 8358
rect 8974 8049 9002 9086
rect 9142 9002 9170 9086
rect 9086 8974 9170 9002
rect 9198 9170 9226 9175
rect 9030 8721 9058 8727
rect 9030 8695 9031 8721
rect 9057 8695 9058 8721
rect 9030 8554 9058 8695
rect 9086 8722 9114 8974
rect 9086 8689 9114 8694
rect 9142 8890 9170 8895
rect 9030 8521 9058 8526
rect 8974 8023 8975 8049
rect 9001 8023 9002 8049
rect 8974 8017 9002 8023
rect 9142 8049 9170 8862
rect 9198 8834 9226 9142
rect 9198 8806 9282 8834
rect 9198 8722 9226 8727
rect 9198 8675 9226 8694
rect 9254 8610 9282 8806
rect 9198 8582 9282 8610
rect 9198 8497 9226 8582
rect 9198 8471 9199 8497
rect 9225 8471 9226 8497
rect 9198 8465 9226 8471
rect 9254 8498 9282 8503
rect 9310 8498 9338 9590
rect 9366 9058 9394 10150
rect 9534 10066 9562 11551
rect 9590 10682 9618 11662
rect 9646 11018 9674 12335
rect 9702 11410 9730 13118
rect 9758 13145 9786 13426
rect 9918 13342 10050 13347
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 9918 13309 10050 13314
rect 10206 13258 10234 13263
rect 9758 13119 9759 13145
rect 9785 13119 9786 13145
rect 9758 12418 9786 13119
rect 10094 13257 10234 13258
rect 10094 13231 10207 13257
rect 10233 13231 10234 13257
rect 10094 13230 10234 13231
rect 9814 12642 9842 12647
rect 9814 12474 9842 12614
rect 9918 12558 10050 12563
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 9918 12525 10050 12530
rect 9814 12446 9898 12474
rect 9758 12385 9786 12390
rect 9814 12361 9842 12367
rect 9814 12335 9815 12361
rect 9841 12335 9842 12361
rect 9758 12306 9786 12311
rect 9814 12306 9842 12335
rect 9786 12278 9842 12306
rect 9758 12273 9786 12278
rect 9870 12250 9898 12446
rect 9814 12222 9898 12250
rect 10094 12417 10122 13230
rect 10206 13225 10234 13230
rect 10262 13257 10290 13454
rect 10262 13231 10263 13257
rect 10289 13231 10290 13257
rect 10262 13225 10290 13231
rect 10318 13202 10346 13207
rect 10094 12391 10095 12417
rect 10121 12391 10122 12417
rect 9814 11774 9842 12222
rect 10094 12194 10122 12391
rect 10094 12161 10122 12166
rect 10150 13146 10178 13151
rect 10150 12362 10178 13118
rect 10318 13145 10346 13174
rect 10318 13119 10319 13145
rect 10345 13119 10346 13145
rect 10318 12642 10346 13119
rect 10374 13145 10402 13454
rect 10598 13435 10626 13454
rect 10374 13119 10375 13145
rect 10401 13119 10402 13145
rect 10374 13113 10402 13119
rect 10654 13145 10682 13566
rect 10710 13481 10738 13566
rect 10710 13455 10711 13481
rect 10737 13455 10738 13481
rect 10710 13449 10738 13455
rect 10766 13481 10794 13487
rect 10766 13455 10767 13481
rect 10793 13455 10794 13481
rect 10766 13202 10794 13455
rect 10766 13169 10794 13174
rect 10654 13119 10655 13145
rect 10681 13119 10682 13145
rect 10654 13113 10682 13119
rect 11214 13146 11242 13151
rect 11046 13090 11074 13095
rect 10990 13089 11074 13090
rect 10990 13063 11047 13089
rect 11073 13063 11074 13089
rect 10990 13062 11074 13063
rect 10822 12754 10850 12759
rect 10318 12609 10346 12614
rect 10766 12753 10850 12754
rect 10766 12727 10823 12753
rect 10849 12727 10850 12753
rect 10766 12726 10850 12727
rect 10766 12642 10794 12726
rect 10822 12721 10850 12726
rect 10934 12753 10962 12759
rect 10934 12727 10935 12753
rect 10961 12727 10962 12753
rect 10094 12082 10122 12087
rect 9982 11913 10010 11919
rect 9982 11887 9983 11913
rect 10009 11887 10010 11913
rect 9982 11858 10010 11887
rect 9982 11825 10010 11830
rect 9758 11746 9842 11774
rect 9918 11774 10050 11779
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 9758 11522 9786 11746
rect 9918 11741 10050 11746
rect 9758 11489 9786 11494
rect 9702 11382 9786 11410
rect 9758 11241 9786 11382
rect 9758 11215 9759 11241
rect 9785 11215 9786 11241
rect 9758 11209 9786 11215
rect 10094 11241 10122 12054
rect 10150 12081 10178 12334
rect 10150 12055 10151 12081
rect 10177 12055 10178 12081
rect 10150 12049 10178 12055
rect 10598 12418 10626 12423
rect 10150 11970 10178 11975
rect 10150 11969 10234 11970
rect 10150 11943 10151 11969
rect 10177 11943 10234 11969
rect 10150 11942 10234 11943
rect 10150 11937 10178 11942
rect 10094 11215 10095 11241
rect 10121 11215 10122 11241
rect 10094 11209 10122 11215
rect 9702 11129 9730 11135
rect 9702 11103 9703 11129
rect 9729 11103 9730 11129
rect 9702 11018 9730 11103
rect 9814 11073 9842 11079
rect 9814 11047 9815 11073
rect 9841 11047 9842 11073
rect 9674 10990 9730 11018
rect 9758 11018 9786 11023
rect 9646 10985 9674 10990
rect 9702 10906 9730 10911
rect 9646 10794 9674 10799
rect 9646 10747 9674 10766
rect 9702 10793 9730 10878
rect 9702 10767 9703 10793
rect 9729 10767 9730 10793
rect 9702 10761 9730 10767
rect 9590 10654 9730 10682
rect 9478 10038 9534 10066
rect 9366 9025 9394 9030
rect 9422 9506 9450 9511
rect 9366 8721 9394 8727
rect 9366 8695 9367 8721
rect 9393 8695 9394 8721
rect 9366 8554 9394 8695
rect 9366 8521 9394 8526
rect 9254 8497 9338 8498
rect 9254 8471 9255 8497
rect 9281 8471 9338 8497
rect 9254 8470 9338 8471
rect 9142 8023 9143 8049
rect 9169 8023 9170 8049
rect 9142 8017 9170 8023
rect 9086 7937 9114 7943
rect 9086 7911 9087 7937
rect 9113 7911 9114 7937
rect 8750 7769 9058 7770
rect 8750 7743 8751 7769
rect 8777 7743 9058 7769
rect 8750 7742 9058 7743
rect 8750 7574 8778 7742
rect 8974 7658 9002 7663
rect 8414 7569 8442 7574
rect 8470 7546 8554 7574
rect 2238 7462 2370 7467
rect 7294 7462 7434 7490
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2238 7429 2370 7434
rect 7406 7265 7434 7462
rect 7406 7239 7407 7265
rect 7433 7239 7434 7265
rect 7406 7233 7434 7239
rect 7798 7210 7826 7215
rect 7798 7209 8274 7210
rect 7798 7183 7799 7209
rect 7825 7183 8274 7209
rect 7798 7182 8274 7183
rect 7798 7177 7826 7182
rect 8246 6817 8274 7182
rect 8302 6930 8330 6935
rect 8302 6883 8330 6902
rect 8414 6874 8442 6879
rect 8414 6827 8442 6846
rect 8246 6791 8247 6817
rect 8273 6791 8274 6817
rect 8246 6785 8274 6791
rect 2238 6678 2370 6683
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2238 6645 2370 6650
rect 2238 5894 2370 5899
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2238 5861 2370 5866
rect 2238 5110 2370 5115
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2238 5077 2370 5082
rect 2238 4326 2370 4331
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2238 4293 2370 4298
rect 2238 3542 2370 3547
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2238 3509 2370 3514
rect 2238 2758 2370 2763
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2238 2725 2370 2730
rect 8526 2170 8554 7546
rect 8694 7546 8778 7574
rect 8918 7602 8946 7621
rect 8918 7569 8946 7574
rect 8694 6762 8722 7546
rect 8694 6481 8722 6734
rect 8694 6455 8695 6481
rect 8721 6455 8722 6481
rect 8694 6449 8722 6455
rect 8862 7321 8890 7327
rect 8862 7295 8863 7321
rect 8889 7295 8890 7321
rect 8862 6426 8890 7295
rect 8974 6929 9002 7630
rect 9030 7574 9058 7742
rect 9086 7657 9114 7911
rect 9086 7631 9087 7657
rect 9113 7631 9114 7657
rect 9086 7625 9114 7631
rect 9254 7658 9282 8470
rect 9366 8442 9394 8447
rect 9422 8442 9450 9478
rect 9366 8441 9450 8442
rect 9366 8415 9367 8441
rect 9393 8415 9450 8441
rect 9366 8414 9450 8415
rect 9478 8441 9506 10038
rect 9534 10033 9562 10038
rect 9590 10401 9618 10407
rect 9590 10375 9591 10401
rect 9617 10375 9618 10401
rect 9590 9786 9618 10375
rect 9534 9758 9618 9786
rect 9646 10290 9674 10295
rect 9534 9282 9562 9758
rect 9646 9673 9674 10262
rect 9646 9647 9647 9673
rect 9673 9647 9674 9673
rect 9590 9617 9618 9623
rect 9590 9591 9591 9617
rect 9617 9591 9618 9617
rect 9590 9450 9618 9591
rect 9590 9417 9618 9422
rect 9534 9249 9562 9254
rect 9478 8415 9479 8441
rect 9505 8415 9506 8441
rect 9366 8409 9394 8414
rect 9478 8409 9506 8415
rect 9534 9058 9562 9063
rect 9310 8162 9338 8167
rect 9310 8049 9338 8134
rect 9478 8162 9506 8167
rect 9534 8162 9562 9030
rect 9646 8890 9674 9647
rect 9646 8843 9674 8862
rect 9702 9337 9730 10654
rect 9758 9729 9786 10990
rect 9814 10850 9842 11047
rect 10038 11074 10066 11093
rect 10038 11041 10066 11046
rect 10150 11074 10178 11079
rect 9918 10990 10050 10995
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 9918 10957 10050 10962
rect 10150 10906 10178 11046
rect 10150 10873 10178 10878
rect 9870 10850 9898 10855
rect 9814 10849 9898 10850
rect 9814 10823 9871 10849
rect 9897 10823 9898 10849
rect 9814 10822 9898 10823
rect 9870 10817 9898 10822
rect 9814 10682 9842 10687
rect 9814 10635 9842 10654
rect 10038 10458 10066 10463
rect 9758 9703 9759 9729
rect 9785 9703 9786 9729
rect 9758 9697 9786 9703
rect 9814 10457 10066 10458
rect 9814 10431 10039 10457
rect 10065 10431 10066 10457
rect 9814 10430 10066 10431
rect 9702 9311 9703 9337
rect 9729 9311 9730 9337
rect 9478 8161 9562 8162
rect 9478 8135 9479 8161
rect 9505 8135 9562 8161
rect 9478 8134 9562 8135
rect 9478 8129 9506 8134
rect 9310 8023 9311 8049
rect 9337 8023 9338 8049
rect 9310 8017 9338 8023
rect 9422 8050 9450 8055
rect 9254 7625 9282 7630
rect 9142 7602 9170 7621
rect 9422 7574 9450 8022
rect 9702 7714 9730 9311
rect 9702 7657 9730 7686
rect 9702 7631 9703 7657
rect 9729 7631 9730 7657
rect 9702 7625 9730 7631
rect 9758 7938 9786 7943
rect 9030 7546 9114 7574
rect 9142 7569 9170 7574
rect 9086 7321 9114 7546
rect 9086 7295 9087 7321
rect 9113 7295 9114 7321
rect 9086 7289 9114 7295
rect 9310 7546 9450 7574
rect 9758 7574 9786 7910
rect 9814 7770 9842 10430
rect 10038 10425 10066 10430
rect 10094 10402 10122 10407
rect 9982 10346 10010 10351
rect 9982 10299 10010 10318
rect 9918 10206 10050 10211
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 9918 10173 10050 10178
rect 10094 10010 10122 10374
rect 10206 10402 10234 11942
rect 10430 11914 10458 11919
rect 10430 11634 10458 11886
rect 10430 11587 10458 11606
rect 10262 11130 10290 11135
rect 10262 11083 10290 11102
rect 10598 11018 10626 12390
rect 10654 12417 10682 12423
rect 10654 12391 10655 12417
rect 10681 12391 10682 12417
rect 10654 12306 10682 12391
rect 10654 12273 10682 12278
rect 10710 12082 10738 12087
rect 10766 12082 10794 12614
rect 10878 12698 10906 12703
rect 10710 12081 10794 12082
rect 10710 12055 10711 12081
rect 10737 12055 10794 12081
rect 10710 12054 10794 12055
rect 10822 12362 10850 12367
rect 10878 12362 10906 12670
rect 10822 12361 10906 12362
rect 10822 12335 10823 12361
rect 10849 12335 10906 12361
rect 10822 12334 10906 12335
rect 10710 12049 10738 12054
rect 10654 11913 10682 11919
rect 10654 11887 10655 11913
rect 10681 11887 10682 11913
rect 10654 11186 10682 11887
rect 10654 11153 10682 11158
rect 10710 11857 10738 11863
rect 10710 11831 10711 11857
rect 10737 11831 10738 11857
rect 10710 11074 10738 11831
rect 10710 11041 10738 11046
rect 10598 10985 10626 10990
rect 10710 10906 10738 10911
rect 10710 10877 10738 10878
rect 10374 10849 10402 10855
rect 10374 10823 10375 10849
rect 10401 10823 10402 10849
rect 10710 10851 10711 10877
rect 10737 10851 10738 10877
rect 10710 10845 10738 10851
rect 10262 10793 10290 10799
rect 10262 10767 10263 10793
rect 10289 10767 10290 10793
rect 10262 10458 10290 10767
rect 10374 10738 10402 10823
rect 10654 10793 10682 10799
rect 10654 10767 10655 10793
rect 10681 10767 10682 10793
rect 10654 10738 10682 10767
rect 10374 10705 10402 10710
rect 10430 10710 10682 10738
rect 10262 10430 10346 10458
rect 10150 10066 10178 10071
rect 10150 10019 10178 10038
rect 10094 9977 10122 9982
rect 10206 9954 10234 10374
rect 10318 10290 10346 10430
rect 10374 10290 10402 10295
rect 10318 10262 10374 10290
rect 10374 10257 10402 10262
rect 10206 9921 10234 9926
rect 10206 9842 10234 9847
rect 10094 9786 10122 9791
rect 10094 9617 10122 9758
rect 10094 9591 10095 9617
rect 10121 9591 10122 9617
rect 10094 9585 10122 9591
rect 10206 9674 10234 9814
rect 10206 9617 10234 9646
rect 10206 9591 10207 9617
rect 10233 9591 10234 9617
rect 10206 9585 10234 9591
rect 10262 9673 10290 9679
rect 10262 9647 10263 9673
rect 10289 9647 10290 9673
rect 9918 9422 10050 9427
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 9918 9389 10050 9394
rect 9870 9338 9898 9343
rect 9870 9225 9898 9310
rect 9870 9199 9871 9225
rect 9897 9199 9898 9225
rect 9870 9193 9898 9199
rect 10094 9170 10122 9175
rect 9870 8778 9898 8783
rect 9870 8731 9898 8750
rect 10094 8777 10122 9142
rect 10094 8751 10095 8777
rect 10121 8751 10122 8777
rect 10094 8745 10122 8751
rect 9918 8638 10050 8643
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 9918 8605 10050 8610
rect 10038 8554 10066 8559
rect 10038 8049 10066 8526
rect 10262 8106 10290 9647
rect 10374 9674 10402 9679
rect 10374 9562 10402 9646
rect 10318 9506 10346 9511
rect 10318 9459 10346 9478
rect 10374 8833 10402 9534
rect 10374 8807 10375 8833
rect 10401 8807 10402 8833
rect 10374 8801 10402 8807
rect 10430 8889 10458 10710
rect 10710 10681 10738 10687
rect 10710 10655 10711 10681
rect 10737 10655 10738 10681
rect 10710 10570 10738 10655
rect 10710 10537 10738 10542
rect 10822 10513 10850 12334
rect 10878 11858 10906 11863
rect 10878 11130 10906 11830
rect 10934 11746 10962 12727
rect 10990 12641 11018 13062
rect 11046 13057 11074 13062
rect 11046 12754 11074 12759
rect 11046 12753 11186 12754
rect 11046 12727 11047 12753
rect 11073 12727 11186 12753
rect 11046 12726 11186 12727
rect 11046 12721 11074 12726
rect 10990 12615 10991 12641
rect 11017 12615 11018 12641
rect 10990 12609 11018 12615
rect 11158 12586 11186 12726
rect 11214 12697 11242 13118
rect 11942 13090 11970 13846
rect 12054 13454 12082 15946
rect 17598 15302 17730 15307
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17598 15269 17730 15274
rect 17598 14518 17730 14523
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17598 14485 17730 14490
rect 17598 13734 17730 13739
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17598 13701 17730 13706
rect 20006 13593 20034 13599
rect 20006 13567 20007 13593
rect 20033 13567 20034 13593
rect 13454 13538 13482 13543
rect 13454 13491 13482 13510
rect 14238 13538 14266 13543
rect 12222 13482 12250 13487
rect 12054 13426 12138 13454
rect 11214 12671 11215 12697
rect 11241 12671 11242 12697
rect 11214 12665 11242 12671
rect 11326 12753 11354 12759
rect 11326 12727 11327 12753
rect 11353 12727 11354 12753
rect 11326 12698 11354 12727
rect 11494 12754 11522 12759
rect 11494 12707 11522 12726
rect 11326 12665 11354 12670
rect 11270 12641 11298 12647
rect 11270 12615 11271 12641
rect 11297 12615 11298 12641
rect 11270 12586 11298 12615
rect 11158 12558 11298 12586
rect 11942 12641 11970 13062
rect 12110 13089 12138 13426
rect 12110 13063 12111 13089
rect 12137 13063 12138 13089
rect 12110 12754 12138 13063
rect 12110 12721 12138 12726
rect 12222 12697 12250 13454
rect 13398 13482 13426 13487
rect 13398 13435 13426 13454
rect 12446 13425 12474 13431
rect 12446 13399 12447 13425
rect 12473 13399 12474 13425
rect 12222 12671 12223 12697
rect 12249 12671 12250 12697
rect 12222 12665 12250 12671
rect 12278 13202 12306 13207
rect 12278 12697 12306 13174
rect 12446 13146 12474 13399
rect 14238 13258 14266 13510
rect 18830 13538 18858 13543
rect 18830 13491 18858 13510
rect 14070 13257 14266 13258
rect 14070 13231 14239 13257
rect 14265 13231 14266 13257
rect 14070 13230 14266 13231
rect 12614 13146 12642 13151
rect 12446 13145 12642 13146
rect 12446 13119 12615 13145
rect 12641 13119 12642 13145
rect 12446 13118 12642 13119
rect 12334 13090 12362 13095
rect 12446 13090 12474 13118
rect 12362 13062 12474 13090
rect 12334 13043 12362 13062
rect 12502 12810 12530 12815
rect 12502 12763 12530 12782
rect 12278 12671 12279 12697
rect 12305 12671 12306 12697
rect 12278 12665 12306 12671
rect 12446 12753 12474 12759
rect 12446 12727 12447 12753
rect 12473 12727 12474 12753
rect 11942 12615 11943 12641
rect 11969 12615 11970 12641
rect 11718 12194 11746 12199
rect 11662 11970 11690 11975
rect 11438 11913 11466 11919
rect 11438 11887 11439 11913
rect 11465 11887 11466 11913
rect 11270 11858 11298 11863
rect 11270 11811 11298 11830
rect 11326 11857 11354 11863
rect 11326 11831 11327 11857
rect 11353 11831 11354 11857
rect 10934 11713 10962 11718
rect 10934 11634 10962 11639
rect 10934 11185 10962 11606
rect 11270 11242 11298 11247
rect 11326 11242 11354 11831
rect 11270 11241 11354 11242
rect 11270 11215 11271 11241
rect 11297 11215 11354 11241
rect 11270 11214 11354 11215
rect 11382 11857 11410 11863
rect 11382 11831 11383 11857
rect 11409 11831 11410 11857
rect 11270 11209 11298 11214
rect 10934 11159 10935 11185
rect 10961 11159 10962 11185
rect 10934 11153 10962 11159
rect 10878 10850 10906 11102
rect 11382 10850 11410 11831
rect 11438 11354 11466 11887
rect 11494 11354 11522 11359
rect 11438 11326 11494 11354
rect 11494 11321 11522 11326
rect 10878 10817 10906 10822
rect 11214 10822 11410 10850
rect 11606 11074 11634 11079
rect 11606 10850 11634 11046
rect 10934 10794 10962 10799
rect 10934 10747 10962 10766
rect 11214 10793 11242 10822
rect 11214 10767 11215 10793
rect 11241 10767 11242 10793
rect 11214 10761 11242 10767
rect 10822 10487 10823 10513
rect 10849 10487 10850 10513
rect 10822 10481 10850 10487
rect 11214 10626 11242 10631
rect 11158 10458 11186 10463
rect 11046 10402 11074 10407
rect 11046 10355 11074 10374
rect 10654 10345 10682 10351
rect 10654 10319 10655 10345
rect 10681 10319 10682 10345
rect 10654 9674 10682 10319
rect 10766 10290 10794 10295
rect 10654 9641 10682 9646
rect 10710 9730 10738 9735
rect 10598 9618 10626 9623
rect 10542 9394 10570 9399
rect 10542 9337 10570 9366
rect 10542 9311 10543 9337
rect 10569 9311 10570 9337
rect 10542 9305 10570 9311
rect 10598 9338 10626 9590
rect 10710 9617 10738 9702
rect 10710 9591 10711 9617
rect 10737 9591 10738 9617
rect 10710 9585 10738 9591
rect 10654 9562 10682 9567
rect 10654 9506 10682 9534
rect 10710 9506 10738 9511
rect 10654 9505 10738 9506
rect 10654 9479 10711 9505
rect 10737 9479 10738 9505
rect 10654 9478 10738 9479
rect 10710 9473 10738 9478
rect 10654 9338 10682 9343
rect 10598 9337 10682 9338
rect 10598 9311 10655 9337
rect 10681 9311 10682 9337
rect 10598 9310 10682 9311
rect 10654 9305 10682 9310
rect 10430 8863 10431 8889
rect 10457 8863 10458 8889
rect 10430 8554 10458 8863
rect 10038 8023 10039 8049
rect 10065 8023 10066 8049
rect 10038 8017 10066 8023
rect 10094 8078 10262 8106
rect 9982 7938 10010 7957
rect 9982 7905 10010 7910
rect 9918 7854 10050 7859
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 9918 7821 10050 7826
rect 9814 7742 10066 7770
rect 9814 7658 9842 7677
rect 9814 7625 9842 7630
rect 8974 6903 8975 6929
rect 9001 6903 9002 6929
rect 8974 6897 9002 6903
rect 9142 6985 9170 6991
rect 9142 6959 9143 6985
rect 9169 6959 9170 6985
rect 9142 6930 9170 6959
rect 9142 6897 9170 6902
rect 9310 6930 9338 7546
rect 9086 6873 9114 6879
rect 9086 6847 9087 6873
rect 9113 6847 9114 6873
rect 9030 6818 9058 6823
rect 9030 6537 9058 6790
rect 9030 6511 9031 6537
rect 9057 6511 9058 6537
rect 9030 6505 9058 6511
rect 9086 6426 9114 6847
rect 9310 6873 9338 6902
rect 9310 6847 9311 6873
rect 9337 6847 9338 6873
rect 9310 6841 9338 6847
rect 9534 7545 9562 7551
rect 9758 7546 9842 7574
rect 9534 7519 9535 7545
rect 9561 7519 9562 7545
rect 9534 7266 9562 7519
rect 9534 6874 9562 7238
rect 9814 6930 9842 7546
rect 10038 7377 10066 7742
rect 10094 7713 10122 8078
rect 10262 8049 10290 8078
rect 10262 8023 10263 8049
rect 10289 8023 10290 8049
rect 10262 8017 10290 8023
rect 10318 8526 10430 8554
rect 10150 7994 10178 7999
rect 10178 7966 10234 7994
rect 10150 7947 10178 7966
rect 10206 7769 10234 7966
rect 10206 7743 10207 7769
rect 10233 7743 10234 7769
rect 10206 7737 10234 7743
rect 10318 7769 10346 8526
rect 10430 8521 10458 8526
rect 10598 9169 10626 9175
rect 10598 9143 10599 9169
rect 10625 9143 10626 9169
rect 10374 8050 10402 8055
rect 10598 8050 10626 9143
rect 10710 8778 10738 8783
rect 10766 8778 10794 10262
rect 11158 9730 11186 10430
rect 11214 10346 11242 10598
rect 11270 10514 11298 10822
rect 11550 10793 11578 10799
rect 11550 10767 11551 10793
rect 11577 10767 11578 10793
rect 11494 10738 11522 10743
rect 11270 10481 11298 10486
rect 11438 10710 11494 10738
rect 11382 10458 11410 10463
rect 11382 10401 11410 10430
rect 11382 10375 11383 10401
rect 11409 10375 11410 10401
rect 11382 10369 11410 10375
rect 11214 10299 11242 10318
rect 11382 10122 11410 10127
rect 11326 10066 11354 10071
rect 11158 9702 11242 9730
rect 10934 9562 10962 9567
rect 10962 9534 11018 9562
rect 10934 9515 10962 9534
rect 10990 9338 11018 9534
rect 11102 9561 11130 9567
rect 11102 9535 11103 9561
rect 11129 9535 11130 9561
rect 11046 9338 11074 9343
rect 10878 9337 11074 9338
rect 10878 9311 11047 9337
rect 11073 9311 11074 9337
rect 10878 9310 11074 9311
rect 10878 9225 10906 9310
rect 11046 9305 11074 9310
rect 10878 9199 10879 9225
rect 10905 9199 10906 9225
rect 10878 9193 10906 9199
rect 11046 9114 11074 9119
rect 11102 9114 11130 9535
rect 11074 9086 11130 9114
rect 11158 9338 11186 9343
rect 11046 9081 11074 9086
rect 10822 9058 10850 9063
rect 10822 8945 10850 9030
rect 10822 8919 10823 8945
rect 10849 8919 10850 8945
rect 10822 8913 10850 8919
rect 11158 8833 11186 9310
rect 11214 9225 11242 9702
rect 11214 9199 11215 9225
rect 11241 9199 11242 9225
rect 11214 9193 11242 9199
rect 11326 9394 11354 10038
rect 11158 8807 11159 8833
rect 11185 8807 11186 8833
rect 11158 8801 11186 8807
rect 10738 8750 10794 8778
rect 11326 8777 11354 9366
rect 11382 9506 11410 10094
rect 11382 9337 11410 9478
rect 11382 9311 11383 9337
rect 11409 9311 11410 9337
rect 11382 9305 11410 9311
rect 11438 9338 11466 10710
rect 11494 10705 11522 10710
rect 11550 10570 11578 10767
rect 11494 10542 11578 10570
rect 11494 10402 11522 10542
rect 11494 10369 11522 10374
rect 11550 10346 11578 10351
rect 11606 10346 11634 10822
rect 11662 10737 11690 11942
rect 11718 11018 11746 12166
rect 11942 11634 11970 12615
rect 12110 12642 12138 12647
rect 12110 12595 12138 12614
rect 12446 12474 12474 12727
rect 12614 12754 12642 13118
rect 13006 13089 13034 13095
rect 13006 13063 13007 13089
rect 13033 13063 13034 13089
rect 13006 12810 13034 13063
rect 14070 13089 14098 13230
rect 14238 13225 14266 13230
rect 19950 13426 19978 13431
rect 14406 13202 14434 13207
rect 14406 13155 14434 13174
rect 18830 13146 18858 13151
rect 18830 13099 18858 13118
rect 14070 13063 14071 13089
rect 14097 13063 14098 13089
rect 14070 13057 14098 13063
rect 19950 13089 19978 13398
rect 20006 13146 20034 13567
rect 20006 13113 20034 13118
rect 19950 13063 19951 13089
rect 19977 13063 19978 13089
rect 19950 13057 19978 13063
rect 17598 12950 17730 12955
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17598 12917 17730 12922
rect 13006 12777 13034 12782
rect 14126 12809 14154 12815
rect 14126 12783 14127 12809
rect 14153 12783 14154 12809
rect 12670 12754 12698 12759
rect 12614 12753 12698 12754
rect 12614 12727 12671 12753
rect 12697 12727 12698 12753
rect 12614 12726 12698 12727
rect 12670 12721 12698 12726
rect 13678 12754 13706 12759
rect 13062 12698 13090 12703
rect 13062 12697 13146 12698
rect 13062 12671 13063 12697
rect 13089 12671 13146 12697
rect 13062 12670 13146 12671
rect 13062 12665 13090 12670
rect 12446 12441 12474 12446
rect 12726 12642 12754 12647
rect 12726 12473 12754 12614
rect 12726 12447 12727 12473
rect 12753 12447 12754 12473
rect 12726 12441 12754 12447
rect 12950 12474 12978 12479
rect 12838 12418 12866 12423
rect 12838 12371 12866 12390
rect 12894 12417 12922 12423
rect 12894 12391 12895 12417
rect 12921 12391 12922 12417
rect 12838 12306 12866 12311
rect 12838 11858 12866 12278
rect 12894 11970 12922 12391
rect 12950 12417 12978 12446
rect 12950 12391 12951 12417
rect 12977 12391 12978 12417
rect 12950 12081 12978 12391
rect 13118 12305 13146 12670
rect 13622 12418 13650 12423
rect 13622 12371 13650 12390
rect 13678 12417 13706 12726
rect 14126 12754 14154 12783
rect 20006 12809 20034 12815
rect 20006 12783 20007 12809
rect 20033 12783 20034 12809
rect 14126 12721 14154 12726
rect 18830 12754 18858 12759
rect 18830 12707 18858 12726
rect 20006 12474 20034 12783
rect 20006 12441 20034 12446
rect 13678 12391 13679 12417
rect 13705 12391 13706 12417
rect 13678 12385 13706 12391
rect 13118 12279 13119 12305
rect 13145 12279 13146 12305
rect 13118 12273 13146 12279
rect 17598 12166 17730 12171
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17598 12133 17730 12138
rect 12950 12055 12951 12081
rect 12977 12055 12978 12081
rect 12950 12049 12978 12055
rect 12894 11937 12922 11942
rect 13006 11913 13034 11919
rect 13006 11887 13007 11913
rect 13033 11887 13034 11913
rect 12950 11858 12978 11863
rect 12838 11857 12978 11858
rect 12838 11831 12951 11857
rect 12977 11831 12978 11857
rect 12838 11830 12978 11831
rect 11942 11601 11970 11606
rect 12558 11634 12586 11639
rect 11998 11354 12026 11359
rect 11718 10990 11802 11018
rect 11662 10711 11663 10737
rect 11689 10711 11690 10737
rect 11662 10705 11690 10711
rect 11718 10906 11746 10911
rect 11718 10849 11746 10878
rect 11718 10823 11719 10849
rect 11745 10823 11746 10849
rect 11718 10738 11746 10823
rect 11718 10705 11746 10710
rect 11774 10402 11802 10990
rect 11998 10905 12026 11326
rect 11998 10879 11999 10905
rect 12025 10879 12026 10905
rect 11998 10873 12026 10879
rect 12334 11298 12362 11303
rect 12334 11241 12362 11270
rect 12334 11215 12335 11241
rect 12361 11215 12362 11241
rect 12054 10849 12082 10855
rect 12054 10823 12055 10849
rect 12081 10823 12082 10849
rect 11942 10794 11970 10799
rect 11830 10402 11858 10407
rect 11550 10345 11634 10346
rect 11550 10319 11551 10345
rect 11577 10319 11634 10345
rect 11550 10318 11634 10319
rect 11718 10401 11858 10402
rect 11718 10375 11831 10401
rect 11857 10375 11858 10401
rect 11718 10374 11858 10375
rect 11550 10313 11578 10318
rect 11718 9730 11746 10374
rect 11830 10369 11858 10374
rect 11886 10346 11914 10351
rect 11886 9954 11914 10318
rect 11942 10066 11970 10766
rect 12054 10682 12082 10823
rect 12110 10850 12138 10855
rect 12110 10803 12138 10822
rect 12334 10793 12362 11215
rect 12558 11241 12586 11606
rect 12558 11215 12559 11241
rect 12585 11215 12586 11241
rect 12558 11186 12586 11215
rect 12894 11186 12922 11191
rect 12586 11158 12698 11186
rect 12558 11153 12586 11158
rect 12334 10767 12335 10793
rect 12361 10767 12362 10793
rect 12334 10761 12362 10767
rect 12670 10905 12698 11158
rect 12894 11139 12922 11158
rect 12950 11018 12978 11830
rect 13006 11074 13034 11887
rect 13734 11634 13762 11639
rect 13678 11633 13762 11634
rect 13678 11607 13735 11633
rect 13761 11607 13762 11633
rect 13678 11606 13762 11607
rect 13510 11577 13538 11583
rect 13510 11551 13511 11577
rect 13537 11551 13538 11577
rect 13230 11186 13258 11191
rect 13230 11185 13370 11186
rect 13230 11159 13231 11185
rect 13257 11159 13370 11185
rect 13230 11158 13370 11159
rect 13230 11153 13258 11158
rect 13006 11046 13314 11074
rect 12950 10990 13258 11018
rect 12670 10879 12671 10905
rect 12697 10879 12698 10905
rect 11998 10402 12026 10407
rect 12054 10402 12082 10654
rect 12670 10458 12698 10879
rect 13230 10458 13258 10990
rect 13286 10794 13314 11046
rect 13342 10905 13370 11158
rect 13342 10879 13343 10905
rect 13369 10879 13370 10905
rect 13342 10873 13370 10879
rect 13510 10906 13538 11551
rect 13622 11577 13650 11583
rect 13622 11551 13623 11577
rect 13649 11551 13650 11577
rect 13454 10850 13482 10855
rect 13510 10850 13538 10878
rect 13454 10849 13538 10850
rect 13454 10823 13455 10849
rect 13481 10823 13538 10849
rect 13454 10822 13538 10823
rect 13566 11521 13594 11527
rect 13566 11495 13567 11521
rect 13593 11495 13594 11521
rect 13566 10849 13594 11495
rect 13622 11186 13650 11551
rect 13622 11153 13650 11158
rect 13566 10823 13567 10849
rect 13593 10823 13594 10849
rect 13454 10817 13482 10822
rect 13566 10817 13594 10823
rect 13678 10794 13706 11606
rect 13734 11601 13762 11606
rect 18830 11577 18858 11583
rect 18830 11551 18831 11577
rect 18857 11551 18858 11577
rect 17598 11382 17730 11387
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17598 11349 17730 11354
rect 18830 11298 18858 11551
rect 20006 11466 20034 11471
rect 20006 11419 20034 11438
rect 18830 11265 18858 11270
rect 14294 11241 14322 11247
rect 14294 11215 14295 11241
rect 14321 11215 14322 11241
rect 14294 11186 14322 11215
rect 20006 11241 20034 11247
rect 20006 11215 20007 11241
rect 20033 11215 20034 11241
rect 14294 11153 14322 11158
rect 18830 11186 18858 11191
rect 18830 11139 18858 11158
rect 20006 11130 20034 11215
rect 20006 11097 20034 11102
rect 18830 10794 18858 10799
rect 13286 10793 13370 10794
rect 13286 10767 13287 10793
rect 13313 10767 13370 10793
rect 13286 10766 13370 10767
rect 13286 10761 13314 10766
rect 12670 10457 12866 10458
rect 12670 10431 12671 10457
rect 12697 10431 12866 10457
rect 12670 10430 12866 10431
rect 13230 10430 13314 10458
rect 12670 10425 12698 10430
rect 11998 10401 12082 10402
rect 11998 10375 11999 10401
rect 12025 10375 12082 10401
rect 11998 10374 12082 10375
rect 12838 10401 12866 10430
rect 12838 10375 12839 10401
rect 12865 10375 12866 10401
rect 11998 10369 12026 10374
rect 12838 10369 12866 10375
rect 12110 10346 12138 10351
rect 13230 10346 13258 10351
rect 12110 10299 12138 10318
rect 12950 10345 13258 10346
rect 12950 10319 13231 10345
rect 13257 10319 13258 10345
rect 12950 10318 13258 10319
rect 11942 10033 11970 10038
rect 12166 10289 12194 10295
rect 12166 10263 12167 10289
rect 12193 10263 12194 10289
rect 11942 9954 11970 9959
rect 11886 9926 11942 9954
rect 11942 9907 11970 9926
rect 11718 9702 11970 9730
rect 11550 9673 11578 9679
rect 11550 9647 11551 9673
rect 11577 9647 11578 9673
rect 11494 9338 11522 9343
rect 11438 9337 11522 9338
rect 11438 9311 11495 9337
rect 11521 9311 11522 9337
rect 11438 9310 11522 9311
rect 11494 9305 11522 9310
rect 11438 9226 11466 9231
rect 11438 9179 11466 9198
rect 11550 9114 11578 9647
rect 11662 9617 11690 9623
rect 11662 9591 11663 9617
rect 11689 9591 11690 9617
rect 11662 9562 11690 9591
rect 11662 9529 11690 9534
rect 11718 9505 11746 9702
rect 11718 9479 11719 9505
rect 11745 9479 11746 9505
rect 11718 9473 11746 9479
rect 11774 9618 11802 9623
rect 11774 9282 11802 9590
rect 11942 9617 11970 9702
rect 11942 9591 11943 9617
rect 11969 9591 11970 9617
rect 11942 9585 11970 9591
rect 12110 9618 12138 9623
rect 12110 9571 12138 9590
rect 11998 9506 12026 9511
rect 11998 9459 12026 9478
rect 11718 9254 11802 9282
rect 11718 9225 11746 9254
rect 11718 9199 11719 9225
rect 11745 9199 11746 9225
rect 11718 9193 11746 9199
rect 11578 9086 11690 9114
rect 11550 9081 11578 9086
rect 11662 8833 11690 9086
rect 11662 8807 11663 8833
rect 11689 8807 11690 8833
rect 11662 8801 11690 8807
rect 11326 8751 11327 8777
rect 11353 8751 11354 8777
rect 10710 8731 10738 8750
rect 11326 8745 11354 8751
rect 10990 8722 11018 8727
rect 10990 8721 11130 8722
rect 10990 8695 10991 8721
rect 11017 8695 11130 8721
rect 10990 8694 11130 8695
rect 10990 8689 11018 8694
rect 10934 8497 10962 8503
rect 10934 8471 10935 8497
rect 10961 8471 10962 8497
rect 10934 8442 10962 8471
rect 10766 8106 10794 8111
rect 10654 8050 10682 8055
rect 10374 8049 10682 8050
rect 10374 8023 10375 8049
rect 10401 8023 10655 8049
rect 10681 8023 10682 8049
rect 10374 8022 10682 8023
rect 10374 8017 10402 8022
rect 10654 8017 10682 8022
rect 10766 8049 10794 8078
rect 10766 8023 10767 8049
rect 10793 8023 10794 8049
rect 10766 8017 10794 8023
rect 10822 7937 10850 7943
rect 10822 7911 10823 7937
rect 10849 7911 10850 7937
rect 10822 7770 10850 7911
rect 10878 7938 10906 7943
rect 10878 7891 10906 7910
rect 10318 7743 10319 7769
rect 10345 7743 10346 7769
rect 10318 7737 10346 7743
rect 10766 7742 10850 7770
rect 10094 7687 10095 7713
rect 10121 7687 10122 7713
rect 10094 7681 10122 7687
rect 10038 7351 10039 7377
rect 10065 7351 10066 7377
rect 10038 7345 10066 7351
rect 10150 7602 10178 7607
rect 10150 7545 10178 7574
rect 10150 7519 10151 7545
rect 10177 7519 10178 7545
rect 10150 7377 10178 7519
rect 10150 7351 10151 7377
rect 10177 7351 10178 7377
rect 10150 7345 10178 7351
rect 10766 7322 10794 7742
rect 10934 7574 10962 8414
rect 10990 8050 11018 8055
rect 10990 8003 11018 8022
rect 10766 7289 10794 7294
rect 10822 7546 10962 7574
rect 11102 7574 11130 8694
rect 11830 8721 11858 8727
rect 11830 8695 11831 8721
rect 11857 8695 11858 8721
rect 11830 7994 11858 8695
rect 12166 8050 12194 10263
rect 12950 10121 12978 10318
rect 13230 10313 13258 10318
rect 12950 10095 12951 10121
rect 12977 10095 12978 10121
rect 12950 10089 12978 10095
rect 12894 10010 12922 10015
rect 12894 9963 12922 9982
rect 13006 10009 13034 10015
rect 13006 9983 13007 10009
rect 13033 9983 13034 10009
rect 12782 9954 12810 9959
rect 12782 9907 12810 9926
rect 13006 9954 13034 9983
rect 13230 10010 13258 10015
rect 13230 9963 13258 9982
rect 13006 9921 13034 9926
rect 13062 9898 13090 9903
rect 13062 9842 13090 9870
rect 13006 9814 13090 9842
rect 12894 9618 12922 9623
rect 12894 9571 12922 9590
rect 12390 9562 12418 9567
rect 12390 9515 12418 9534
rect 12558 9506 12586 9511
rect 12558 9459 12586 9478
rect 12838 9225 12866 9231
rect 12838 9199 12839 9225
rect 12865 9199 12866 9225
rect 12726 9170 12754 9175
rect 12838 9170 12866 9199
rect 12726 9169 12866 9170
rect 12726 9143 12727 9169
rect 12753 9143 12866 9169
rect 12726 9142 12866 9143
rect 12166 8017 12194 8022
rect 12670 8386 12698 8391
rect 12726 8386 12754 9142
rect 13006 8833 13034 9814
rect 13230 9618 13258 9623
rect 13286 9618 13314 10430
rect 13342 9898 13370 10766
rect 13678 10094 13706 10766
rect 18718 10793 18858 10794
rect 18718 10767 18831 10793
rect 18857 10767 18858 10793
rect 18718 10766 18858 10767
rect 17598 10598 17730 10603
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17598 10565 17730 10570
rect 14294 10457 14322 10463
rect 14294 10431 14295 10457
rect 14321 10431 14322 10457
rect 13566 10066 13706 10094
rect 13790 10346 13818 10351
rect 13566 10065 13594 10066
rect 13566 10039 13567 10065
rect 13593 10039 13594 10065
rect 13566 10033 13594 10039
rect 13790 10065 13818 10318
rect 14294 10346 14322 10431
rect 14294 10313 14322 10318
rect 14630 10401 14658 10407
rect 14630 10375 14631 10401
rect 14657 10375 14658 10401
rect 14630 10346 14658 10375
rect 14630 10313 14658 10318
rect 18718 10346 18746 10766
rect 18830 10761 18858 10766
rect 19950 10737 19978 10743
rect 19950 10711 19951 10737
rect 19977 10711 19978 10737
rect 19950 10458 19978 10711
rect 19950 10425 19978 10430
rect 20006 10457 20034 10463
rect 20006 10431 20007 10457
rect 20033 10431 20034 10457
rect 18830 10402 18858 10407
rect 18830 10355 18858 10374
rect 18718 10313 18746 10318
rect 14742 10290 14770 10295
rect 14742 10243 14770 10262
rect 20006 10122 20034 10431
rect 20006 10089 20034 10094
rect 13790 10039 13791 10065
rect 13817 10039 13818 10065
rect 13790 10033 13818 10039
rect 13678 10010 13706 10015
rect 13678 10009 13762 10010
rect 13678 9983 13679 10009
rect 13705 9983 13762 10009
rect 13678 9982 13762 9983
rect 13678 9977 13706 9982
rect 13622 9954 13650 9959
rect 13622 9907 13650 9926
rect 13342 9865 13370 9870
rect 13230 9617 13314 9618
rect 13230 9591 13231 9617
rect 13257 9591 13314 9617
rect 13230 9590 13314 9591
rect 13230 9585 13258 9590
rect 13118 9562 13146 9567
rect 13118 9515 13146 9534
rect 13062 9505 13090 9511
rect 13062 9479 13063 9505
rect 13089 9479 13090 9505
rect 13062 9338 13090 9479
rect 13062 9310 13258 9338
rect 13230 9281 13258 9310
rect 13230 9255 13231 9281
rect 13257 9255 13258 9281
rect 13230 9249 13258 9255
rect 13006 8807 13007 8833
rect 13033 8807 13034 8833
rect 13006 8801 13034 8807
rect 13230 8834 13258 8839
rect 13286 8834 13314 9590
rect 13678 9618 13706 9623
rect 13566 9562 13594 9567
rect 13566 9515 13594 9534
rect 13678 9561 13706 9590
rect 13678 9535 13679 9561
rect 13705 9535 13706 9561
rect 13678 9529 13706 9535
rect 13734 9561 13762 9982
rect 17598 9814 17730 9819
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17598 9781 17730 9786
rect 20006 9673 20034 9679
rect 20006 9647 20007 9673
rect 20033 9647 20034 9673
rect 13734 9535 13735 9561
rect 13761 9535 13762 9561
rect 13734 9506 13762 9535
rect 13230 8833 13314 8834
rect 13230 8807 13231 8833
rect 13257 8807 13314 8833
rect 13230 8806 13314 8807
rect 13342 8834 13370 8839
rect 13566 8834 13594 8839
rect 13342 8833 13594 8834
rect 13342 8807 13343 8833
rect 13369 8807 13567 8833
rect 13593 8807 13594 8833
rect 13342 8806 13594 8807
rect 13230 8801 13258 8806
rect 13342 8801 13370 8806
rect 13566 8801 13594 8806
rect 13622 8834 13650 8839
rect 13622 8787 13650 8806
rect 13174 8721 13202 8727
rect 13174 8695 13175 8721
rect 13201 8695 13202 8721
rect 13174 8498 13202 8695
rect 13510 8721 13538 8727
rect 13510 8695 13511 8721
rect 13537 8695 13538 8721
rect 13230 8498 13258 8503
rect 13174 8497 13258 8498
rect 13174 8471 13231 8497
rect 13257 8471 13258 8497
rect 13174 8470 13258 8471
rect 13230 8465 13258 8470
rect 12838 8441 12866 8447
rect 12838 8415 12839 8441
rect 12865 8415 12866 8441
rect 12838 8386 12866 8415
rect 13510 8442 13538 8695
rect 13510 8409 13538 8414
rect 13734 8721 13762 9478
rect 14294 9618 14322 9623
rect 14294 9169 14322 9590
rect 18830 9618 18858 9623
rect 18830 9571 18858 9590
rect 20006 9450 20034 9647
rect 20006 9417 20034 9422
rect 14294 9143 14295 9169
rect 14321 9143 14322 9169
rect 14294 9137 14322 9143
rect 17598 9030 17730 9035
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17598 8997 17730 9002
rect 20006 8889 20034 8895
rect 20006 8863 20007 8889
rect 20033 8863 20034 8889
rect 13734 8695 13735 8721
rect 13761 8695 13762 8721
rect 12670 8385 12866 8386
rect 12670 8359 12671 8385
rect 12697 8359 12866 8385
rect 12670 8358 12866 8359
rect 11830 7713 11858 7966
rect 11886 7938 11914 7943
rect 11886 7769 11914 7910
rect 11886 7743 11887 7769
rect 11913 7743 11914 7769
rect 11886 7737 11914 7743
rect 11830 7687 11831 7713
rect 11857 7687 11858 7713
rect 11830 7681 11858 7687
rect 11942 7713 11970 7719
rect 11942 7687 11943 7713
rect 11969 7687 11970 7713
rect 11942 7574 11970 7687
rect 12334 7657 12362 7663
rect 12334 7631 12335 7657
rect 12361 7631 12362 7657
rect 11102 7546 11242 7574
rect 10262 7266 10290 7271
rect 10262 7219 10290 7238
rect 10374 7266 10402 7271
rect 10374 7219 10402 7238
rect 10822 7265 10850 7546
rect 10934 7513 10962 7518
rect 11158 7322 11186 7327
rect 11158 7275 11186 7294
rect 10822 7239 10823 7265
rect 10849 7239 10850 7265
rect 10822 7233 10850 7239
rect 10318 7154 10346 7159
rect 10318 7153 10794 7154
rect 10318 7127 10319 7153
rect 10345 7127 10794 7153
rect 10318 7126 10794 7127
rect 10318 7121 10346 7126
rect 9918 7070 10050 7075
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 9918 7037 10050 7042
rect 9926 6930 9954 6935
rect 9814 6929 9954 6930
rect 9814 6903 9927 6929
rect 9953 6903 9954 6929
rect 9814 6902 9954 6903
rect 9926 6897 9954 6902
rect 10150 6929 10178 6935
rect 10150 6903 10151 6929
rect 10177 6903 10178 6929
rect 9646 6874 9674 6879
rect 9534 6846 9646 6874
rect 9646 6827 9674 6846
rect 9758 6874 9786 6879
rect 9758 6827 9786 6846
rect 10038 6874 10066 6879
rect 10038 6827 10066 6846
rect 9870 6818 9898 6823
rect 9870 6771 9898 6790
rect 10094 6538 10122 6543
rect 10150 6538 10178 6903
rect 10206 6930 10234 6935
rect 10206 6883 10234 6902
rect 10318 6762 10346 6767
rect 10318 6538 10346 6734
rect 10094 6537 10178 6538
rect 10094 6511 10095 6537
rect 10121 6511 10178 6537
rect 10094 6510 10178 6511
rect 10094 6505 10122 6510
rect 8862 6398 9114 6426
rect 8862 2170 8890 2175
rect 8526 2169 8890 2170
rect 8526 2143 8863 2169
rect 8889 2143 8890 2169
rect 8526 2142 8890 2143
rect 8862 2137 8890 2142
rect 8750 2058 8778 2063
rect 2238 1974 2370 1979
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2238 1941 2370 1946
rect 3486 1666 3514 1671
rect 3374 1665 3514 1666
rect 3374 1639 3487 1665
rect 3513 1639 3514 1665
rect 3374 1638 3514 1639
rect 3374 400 3402 1638
rect 3486 1633 3514 1638
rect 8750 400 8778 2030
rect 9030 1778 9058 1783
rect 9086 1778 9114 6398
rect 9918 6286 10050 6291
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 9918 6253 10050 6258
rect 9918 5502 10050 5507
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 9918 5469 10050 5474
rect 9918 4718 10050 4723
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 9918 4685 10050 4690
rect 9918 3934 10050 3939
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 9918 3901 10050 3906
rect 9918 3150 10050 3155
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 9918 3117 10050 3122
rect 9918 2366 10050 2371
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 9918 2333 10050 2338
rect 9366 2058 9394 2063
rect 9366 2011 9394 2030
rect 9030 1777 9114 1778
rect 9030 1751 9031 1777
rect 9057 1751 9114 1777
rect 9030 1750 9114 1751
rect 9310 1833 9338 1839
rect 9310 1807 9311 1833
rect 9337 1807 9338 1833
rect 9030 1745 9058 1750
rect 9310 1694 9338 1807
rect 10150 1778 10178 6510
rect 10262 6537 10346 6538
rect 10262 6511 10319 6537
rect 10345 6511 10346 6537
rect 10262 6510 10346 6511
rect 10262 6089 10290 6510
rect 10318 6505 10346 6510
rect 10766 6481 10794 7126
rect 11214 6874 11242 7546
rect 11830 7546 11858 7551
rect 11942 7546 12250 7574
rect 11270 7266 11298 7271
rect 11270 6985 11298 7238
rect 11270 6959 11271 6985
rect 11297 6959 11298 6985
rect 11270 6953 11298 6959
rect 11214 6827 11242 6846
rect 11382 6873 11410 6879
rect 11382 6847 11383 6873
rect 11409 6847 11410 6873
rect 10766 6455 10767 6481
rect 10793 6455 10794 6481
rect 10766 6449 10794 6455
rect 10654 6370 10682 6375
rect 10598 6369 10682 6370
rect 10598 6343 10655 6369
rect 10681 6343 10682 6369
rect 10598 6342 10682 6343
rect 10598 6145 10626 6342
rect 10654 6337 10682 6342
rect 10598 6119 10599 6145
rect 10625 6119 10626 6145
rect 10598 6113 10626 6119
rect 10262 6063 10263 6089
rect 10289 6063 10290 6089
rect 10262 6057 10290 6063
rect 11382 5922 11410 6847
rect 11830 6538 11858 7518
rect 12222 7321 12250 7546
rect 12334 7546 12362 7631
rect 12670 7574 12698 8358
rect 12950 8330 12978 8335
rect 12950 7994 12978 8302
rect 13062 8050 13090 8055
rect 13062 8003 13090 8022
rect 13286 8050 13314 8055
rect 13454 8050 13482 8055
rect 13286 8049 13482 8050
rect 13286 8023 13287 8049
rect 13313 8023 13455 8049
rect 13481 8023 13482 8049
rect 13286 8022 13482 8023
rect 13286 8017 13314 8022
rect 13454 8017 13482 8022
rect 13622 8050 13650 8055
rect 13734 8050 13762 8695
rect 14294 8834 14322 8839
rect 14294 8385 14322 8806
rect 18830 8834 18858 8839
rect 18830 8787 18858 8806
rect 20006 8778 20034 8863
rect 20006 8745 20034 8750
rect 14294 8359 14295 8385
rect 14321 8359 14322 8385
rect 14294 8353 14322 8359
rect 17598 8246 17730 8251
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17598 8213 17730 8218
rect 20006 8105 20034 8111
rect 20006 8079 20007 8105
rect 20033 8079 20034 8105
rect 13622 8049 13762 8050
rect 13622 8023 13623 8049
rect 13649 8023 13762 8049
rect 13622 8022 13762 8023
rect 18830 8049 18858 8055
rect 18830 8023 18831 8049
rect 18857 8023 18858 8049
rect 13622 8017 13650 8022
rect 12838 7966 12950 7994
rect 12782 7657 12810 7663
rect 12782 7631 12783 7657
rect 12809 7631 12810 7657
rect 12782 7574 12810 7631
rect 12446 7546 12810 7574
rect 12362 7518 12474 7546
rect 12334 7513 12362 7518
rect 12222 7295 12223 7321
rect 12249 7295 12250 7321
rect 12222 6762 12250 7295
rect 12446 7321 12474 7518
rect 12782 7378 12810 7383
rect 12838 7378 12866 7966
rect 12950 7947 12978 7966
rect 13174 7937 13202 7943
rect 13174 7911 13175 7937
rect 13201 7911 13202 7937
rect 13174 7713 13202 7911
rect 13174 7687 13175 7713
rect 13201 7687 13202 7713
rect 13174 7681 13202 7687
rect 13566 7937 13594 7943
rect 13566 7911 13567 7937
rect 13593 7911 13594 7937
rect 13566 7602 13594 7911
rect 13566 7569 13594 7574
rect 14238 7602 14266 7607
rect 14238 7555 14266 7574
rect 18830 7602 18858 8023
rect 20006 7770 20034 8079
rect 20006 7737 20034 7742
rect 18830 7569 18858 7574
rect 17598 7462 17730 7467
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17598 7429 17730 7434
rect 12782 7377 12866 7378
rect 12782 7351 12783 7377
rect 12809 7351 12866 7377
rect 12782 7350 12866 7351
rect 12782 7345 12810 7350
rect 12446 7295 12447 7321
rect 12473 7295 12474 7321
rect 12446 7289 12474 7295
rect 12838 7153 12866 7159
rect 12838 7127 12839 7153
rect 12865 7127 12866 7153
rect 12782 6930 12810 6935
rect 12838 6930 12866 7127
rect 12894 7154 12922 7159
rect 12894 7107 12922 7126
rect 13454 7154 13482 7159
rect 12782 6929 12866 6930
rect 12782 6903 12783 6929
rect 12809 6903 12866 6929
rect 12782 6902 12866 6903
rect 12782 6897 12810 6902
rect 12614 6874 12642 6893
rect 12614 6841 12642 6846
rect 12614 6762 12642 6767
rect 12222 6729 12250 6734
rect 12390 6761 12642 6762
rect 12390 6735 12615 6761
rect 12641 6735 12642 6761
rect 12390 6734 12642 6735
rect 11830 6537 12026 6538
rect 11830 6511 11831 6537
rect 11857 6511 12026 6537
rect 11830 6510 12026 6511
rect 11830 6505 11858 6510
rect 11886 6201 11914 6510
rect 11998 6481 12026 6510
rect 12390 6537 12418 6734
rect 12614 6729 12642 6734
rect 12670 6762 12698 6767
rect 12390 6511 12391 6537
rect 12417 6511 12418 6537
rect 12390 6505 12418 6511
rect 11998 6455 11999 6481
rect 12025 6455 12026 6481
rect 11998 6449 12026 6455
rect 11886 6175 11887 6201
rect 11913 6175 11914 6201
rect 11886 6169 11914 6175
rect 11382 5889 11410 5894
rect 11662 6033 11690 6039
rect 11662 6007 11663 6033
rect 11689 6007 11690 6033
rect 11662 5922 11690 6007
rect 11662 5889 11690 5894
rect 12278 5922 12306 5927
rect 12110 2058 12138 2063
rect 11438 1834 11466 1839
rect 10374 1778 10402 1783
rect 10150 1777 10402 1778
rect 10150 1751 10375 1777
rect 10401 1751 10402 1777
rect 10150 1750 10402 1751
rect 10374 1745 10402 1750
rect 9086 1666 9338 1694
rect 10094 1722 10122 1727
rect 9086 400 9114 1666
rect 9918 1582 10050 1587
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 9918 1549 10050 1554
rect 10094 400 10122 1694
rect 10878 1722 10906 1727
rect 10878 1665 10906 1694
rect 10878 1639 10879 1665
rect 10905 1639 10906 1665
rect 10878 1633 10906 1639
rect 11438 400 11466 1806
rect 12110 400 12138 2030
rect 12278 1777 12306 5894
rect 12670 2169 12698 6734
rect 13454 6538 13482 7126
rect 17598 6678 17730 6683
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17598 6645 17730 6650
rect 13454 6491 13482 6510
rect 14294 6538 14322 6543
rect 12670 2143 12671 2169
rect 12697 2143 12698 2169
rect 12670 2137 12698 2143
rect 13118 2058 13146 2063
rect 13118 2011 13146 2030
rect 12782 1834 12810 1839
rect 12782 1787 12810 1806
rect 13174 1834 13202 1839
rect 12278 1751 12279 1777
rect 12305 1751 12306 1777
rect 12278 1745 12306 1751
rect 13174 1694 13202 1806
rect 14294 1777 14322 6510
rect 17598 5894 17730 5899
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17598 5861 17730 5866
rect 17598 5110 17730 5115
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17598 5077 17730 5082
rect 17598 4326 17730 4331
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17598 4293 17730 4298
rect 17598 3542 17730 3547
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17598 3509 17730 3514
rect 17598 2758 17730 2763
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17598 2725 17730 2730
rect 17598 1974 17730 1979
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17598 1941 17730 1946
rect 14686 1834 14714 1839
rect 14686 1787 14714 1806
rect 14294 1751 14295 1777
rect 14321 1751 14322 1777
rect 14294 1745 14322 1751
rect 13118 1666 13202 1694
rect 13118 400 13146 1666
rect 3360 0 3416 400
rect 8736 0 8792 400
rect 9072 0 9128 400
rect 10080 0 10136 400
rect 11424 0 11480 400
rect 12096 0 12152 400
rect 13104 0 13160 400
<< via2 >>
rect 2238 19221 2266 19222
rect 2238 19195 2239 19221
rect 2239 19195 2265 19221
rect 2265 19195 2266 19221
rect 2238 19194 2266 19195
rect 2290 19221 2318 19222
rect 2290 19195 2291 19221
rect 2291 19195 2317 19221
rect 2317 19195 2318 19221
rect 2290 19194 2318 19195
rect 2342 19221 2370 19222
rect 2342 19195 2343 19221
rect 2343 19195 2369 19221
rect 2369 19195 2370 19221
rect 2342 19194 2370 19195
rect 8750 18718 8778 18746
rect 9366 18745 9394 18746
rect 9366 18719 9367 18745
rect 9367 18719 9393 18745
rect 9393 18719 9394 18745
rect 9366 18718 9394 18719
rect 2238 18437 2266 18438
rect 2238 18411 2239 18437
rect 2239 18411 2265 18437
rect 2265 18411 2266 18437
rect 2238 18410 2266 18411
rect 2290 18437 2318 18438
rect 2290 18411 2291 18437
rect 2291 18411 2317 18437
rect 2317 18411 2318 18437
rect 2290 18410 2318 18411
rect 2342 18437 2370 18438
rect 2342 18411 2343 18437
rect 2343 18411 2369 18437
rect 2369 18411 2370 18437
rect 2342 18410 2370 18411
rect 2238 17653 2266 17654
rect 2238 17627 2239 17653
rect 2239 17627 2265 17653
rect 2265 17627 2266 17653
rect 2238 17626 2266 17627
rect 2290 17653 2318 17654
rect 2290 17627 2291 17653
rect 2291 17627 2317 17653
rect 2317 17627 2318 17653
rect 2290 17626 2318 17627
rect 2342 17653 2370 17654
rect 2342 17627 2343 17653
rect 2343 17627 2369 17653
rect 2369 17627 2370 17653
rect 2342 17626 2370 17627
rect 2238 16869 2266 16870
rect 2238 16843 2239 16869
rect 2239 16843 2265 16869
rect 2265 16843 2266 16869
rect 2238 16842 2266 16843
rect 2290 16869 2318 16870
rect 2290 16843 2291 16869
rect 2291 16843 2317 16869
rect 2317 16843 2318 16869
rect 2290 16842 2318 16843
rect 2342 16869 2370 16870
rect 2342 16843 2343 16869
rect 2343 16843 2369 16869
rect 2369 16843 2370 16869
rect 2342 16842 2370 16843
rect 2238 16085 2266 16086
rect 2238 16059 2239 16085
rect 2239 16059 2265 16085
rect 2265 16059 2266 16085
rect 2238 16058 2266 16059
rect 2290 16085 2318 16086
rect 2290 16059 2291 16085
rect 2291 16059 2317 16085
rect 2317 16059 2318 16085
rect 2290 16058 2318 16059
rect 2342 16085 2370 16086
rect 2342 16059 2343 16085
rect 2343 16059 2369 16085
rect 2369 16059 2370 16085
rect 2342 16058 2370 16059
rect 2238 15301 2266 15302
rect 2238 15275 2239 15301
rect 2239 15275 2265 15301
rect 2265 15275 2266 15301
rect 2238 15274 2266 15275
rect 2290 15301 2318 15302
rect 2290 15275 2291 15301
rect 2291 15275 2317 15301
rect 2317 15275 2318 15301
rect 2290 15274 2318 15275
rect 2342 15301 2370 15302
rect 2342 15275 2343 15301
rect 2343 15275 2369 15301
rect 2369 15275 2370 15301
rect 2342 15274 2370 15275
rect 2238 14517 2266 14518
rect 2238 14491 2239 14517
rect 2239 14491 2265 14517
rect 2265 14491 2266 14517
rect 2238 14490 2266 14491
rect 2290 14517 2318 14518
rect 2290 14491 2291 14517
rect 2291 14491 2317 14517
rect 2317 14491 2318 14517
rect 2290 14490 2318 14491
rect 2342 14517 2370 14518
rect 2342 14491 2343 14517
rect 2343 14491 2369 14517
rect 2369 14491 2370 14517
rect 2342 14490 2370 14491
rect 2086 13790 2114 13818
rect 966 12782 994 12810
rect 1022 12446 1050 12474
rect 2238 13733 2266 13734
rect 2238 13707 2239 13733
rect 2239 13707 2265 13733
rect 2265 13707 2266 13733
rect 2238 13706 2266 13707
rect 2290 13733 2318 13734
rect 2290 13707 2291 13733
rect 2291 13707 2317 13733
rect 2317 13707 2318 13733
rect 2290 13706 2318 13707
rect 2342 13733 2370 13734
rect 2342 13707 2343 13733
rect 2343 13707 2369 13733
rect 2369 13707 2370 13733
rect 2342 13706 2370 13707
rect 9422 13929 9450 13930
rect 9422 13903 9423 13929
rect 9423 13903 9449 13929
rect 9449 13903 9450 13929
rect 9422 13902 9450 13903
rect 9918 18829 9946 18830
rect 9918 18803 9919 18829
rect 9919 18803 9945 18829
rect 9945 18803 9946 18829
rect 9918 18802 9946 18803
rect 9970 18829 9998 18830
rect 9970 18803 9971 18829
rect 9971 18803 9997 18829
rect 9997 18803 9998 18829
rect 9970 18802 9998 18803
rect 10022 18829 10050 18830
rect 10022 18803 10023 18829
rect 10023 18803 10049 18829
rect 10049 18803 10050 18829
rect 10022 18802 10050 18803
rect 10766 19110 10794 19138
rect 10542 18969 10570 18970
rect 10542 18943 10543 18969
rect 10543 18943 10569 18969
rect 10569 18943 10570 18969
rect 10542 18942 10570 18943
rect 10430 18718 10458 18746
rect 9918 18045 9946 18046
rect 9918 18019 9919 18045
rect 9919 18019 9945 18045
rect 9945 18019 9946 18045
rect 9918 18018 9946 18019
rect 9970 18045 9998 18046
rect 9970 18019 9971 18045
rect 9971 18019 9997 18045
rect 9997 18019 9998 18045
rect 9970 18018 9998 18019
rect 10022 18045 10050 18046
rect 10022 18019 10023 18045
rect 10023 18019 10049 18045
rect 10049 18019 10050 18045
rect 10022 18018 10050 18019
rect 9918 17261 9946 17262
rect 9918 17235 9919 17261
rect 9919 17235 9945 17261
rect 9945 17235 9946 17261
rect 9918 17234 9946 17235
rect 9970 17261 9998 17262
rect 9970 17235 9971 17261
rect 9971 17235 9997 17261
rect 9997 17235 9998 17261
rect 9970 17234 9998 17235
rect 10022 17261 10050 17262
rect 10022 17235 10023 17261
rect 10023 17235 10049 17261
rect 10049 17235 10050 17261
rect 10022 17234 10050 17235
rect 9918 16477 9946 16478
rect 9918 16451 9919 16477
rect 9919 16451 9945 16477
rect 9945 16451 9946 16477
rect 9918 16450 9946 16451
rect 9970 16477 9998 16478
rect 9970 16451 9971 16477
rect 9971 16451 9997 16477
rect 9997 16451 9998 16477
rect 9970 16450 9998 16451
rect 10022 16477 10050 16478
rect 10022 16451 10023 16477
rect 10023 16451 10049 16477
rect 10049 16451 10050 16477
rect 10022 16450 10050 16451
rect 9918 15693 9946 15694
rect 9918 15667 9919 15693
rect 9919 15667 9945 15693
rect 9945 15667 9946 15693
rect 9918 15666 9946 15667
rect 9970 15693 9998 15694
rect 9970 15667 9971 15693
rect 9971 15667 9997 15693
rect 9997 15667 9998 15693
rect 9970 15666 9998 15667
rect 10022 15693 10050 15694
rect 10022 15667 10023 15693
rect 10023 15667 10049 15693
rect 10049 15667 10050 15693
rect 10022 15666 10050 15667
rect 9918 14909 9946 14910
rect 9918 14883 9919 14909
rect 9919 14883 9945 14909
rect 9945 14883 9946 14909
rect 9918 14882 9946 14883
rect 9970 14909 9998 14910
rect 9970 14883 9971 14909
rect 9971 14883 9997 14909
rect 9997 14883 9998 14909
rect 9970 14882 9998 14883
rect 10022 14909 10050 14910
rect 10022 14883 10023 14909
rect 10023 14883 10049 14909
rect 10049 14883 10050 14909
rect 10022 14882 10050 14883
rect 9918 14125 9946 14126
rect 9918 14099 9919 14125
rect 9919 14099 9945 14125
rect 9945 14099 9946 14125
rect 9918 14098 9946 14099
rect 9970 14125 9998 14126
rect 9970 14099 9971 14125
rect 9971 14099 9997 14125
rect 9997 14099 9998 14125
rect 9970 14098 9998 14099
rect 10022 14125 10050 14126
rect 10022 14099 10023 14125
rect 10023 14099 10049 14125
rect 10049 14099 10050 14125
rect 10022 14098 10050 14099
rect 10318 14014 10346 14042
rect 9814 13593 9842 13594
rect 9814 13567 9815 13593
rect 9815 13567 9841 13593
rect 9841 13567 9842 13593
rect 9814 13566 9842 13567
rect 2142 13145 2170 13146
rect 2142 13119 2143 13145
rect 2143 13119 2169 13145
rect 2169 13119 2170 13145
rect 2142 13118 2170 13119
rect 5950 13118 5978 13146
rect 2238 12949 2266 12950
rect 2238 12923 2239 12949
rect 2239 12923 2265 12949
rect 2265 12923 2266 12949
rect 2238 12922 2266 12923
rect 2290 12949 2318 12950
rect 2290 12923 2291 12949
rect 2291 12923 2317 12949
rect 2317 12923 2318 12949
rect 2290 12922 2318 12923
rect 2342 12949 2370 12950
rect 2342 12923 2343 12949
rect 2343 12923 2369 12949
rect 2369 12923 2370 12949
rect 2342 12922 2370 12923
rect 2142 12753 2170 12754
rect 2142 12727 2143 12753
rect 2143 12727 2169 12753
rect 2169 12727 2170 12753
rect 2142 12726 2170 12727
rect 5446 12726 5474 12754
rect 2238 12165 2266 12166
rect 2238 12139 2239 12165
rect 2239 12139 2265 12165
rect 2265 12139 2266 12165
rect 2238 12138 2266 12139
rect 2290 12165 2318 12166
rect 2290 12139 2291 12165
rect 2291 12139 2317 12165
rect 2317 12139 2318 12165
rect 2290 12138 2318 12139
rect 2342 12165 2370 12166
rect 2342 12139 2343 12165
rect 2343 12139 2369 12165
rect 2369 12139 2370 12165
rect 2342 12138 2370 12139
rect 5950 12390 5978 12418
rect 7350 13089 7378 13090
rect 7350 13063 7351 13089
rect 7351 13063 7377 13089
rect 7377 13063 7378 13089
rect 7350 13062 7378 13063
rect 8134 13062 8162 13090
rect 6902 12278 6930 12306
rect 6958 12054 6986 12082
rect 7126 12278 7154 12306
rect 5446 11998 5474 12026
rect 6734 12025 6762 12026
rect 6734 11999 6735 12025
rect 6735 11999 6761 12025
rect 6761 11999 6762 12025
rect 6734 11998 6762 11999
rect 7070 11913 7098 11914
rect 7070 11887 7071 11913
rect 7071 11887 7097 11913
rect 7097 11887 7098 11913
rect 7070 11886 7098 11887
rect 6510 11830 6538 11858
rect 7182 12081 7210 12082
rect 7182 12055 7183 12081
rect 7183 12055 7209 12081
rect 7209 12055 7210 12081
rect 7182 12054 7210 12055
rect 7182 11857 7210 11858
rect 7182 11831 7183 11857
rect 7183 11831 7209 11857
rect 7209 11831 7210 11857
rect 7182 11830 7210 11831
rect 7294 11774 7322 11802
rect 7630 12558 7658 12586
rect 8302 12502 8330 12530
rect 7406 12278 7434 12306
rect 7798 12417 7826 12418
rect 7798 12391 7799 12417
rect 7799 12391 7825 12417
rect 7825 12391 7826 12417
rect 7798 12390 7826 12391
rect 8750 13342 8778 13370
rect 9478 13454 9506 13482
rect 11214 19137 11242 19138
rect 11214 19111 11215 19137
rect 11215 19111 11241 19137
rect 11241 19111 11242 19137
rect 11214 19110 11242 19111
rect 17598 19221 17626 19222
rect 17598 19195 17599 19221
rect 17599 19195 17625 19221
rect 17625 19195 17626 19221
rect 17598 19194 17626 19195
rect 17650 19221 17678 19222
rect 17650 19195 17651 19221
rect 17651 19195 17677 19221
rect 17677 19195 17678 19221
rect 17650 19194 17678 19195
rect 17702 19221 17730 19222
rect 17702 19195 17703 19221
rect 17703 19195 17729 19221
rect 17729 19195 17730 19221
rect 17702 19194 17730 19195
rect 12110 19110 12138 19138
rect 12782 19137 12810 19138
rect 12782 19111 12783 19137
rect 12783 19111 12809 19137
rect 12809 19111 12810 19137
rect 12782 19110 12810 19111
rect 11102 18942 11130 18970
rect 11046 18745 11074 18746
rect 11046 18719 11047 18745
rect 11047 18719 11073 18745
rect 11073 18719 11074 18745
rect 11046 18718 11074 18719
rect 10710 13958 10738 13986
rect 17598 18437 17626 18438
rect 17598 18411 17599 18437
rect 17599 18411 17625 18437
rect 17625 18411 17626 18437
rect 17598 18410 17626 18411
rect 17650 18437 17678 18438
rect 17650 18411 17651 18437
rect 17651 18411 17677 18437
rect 17677 18411 17678 18437
rect 17650 18410 17678 18411
rect 17702 18437 17730 18438
rect 17702 18411 17703 18437
rect 17703 18411 17729 18437
rect 17729 18411 17730 18437
rect 17702 18410 17730 18411
rect 17598 17653 17626 17654
rect 17598 17627 17599 17653
rect 17599 17627 17625 17653
rect 17625 17627 17626 17653
rect 17598 17626 17626 17627
rect 17650 17653 17678 17654
rect 17650 17627 17651 17653
rect 17651 17627 17677 17653
rect 17677 17627 17678 17653
rect 17650 17626 17678 17627
rect 17702 17653 17730 17654
rect 17702 17627 17703 17653
rect 17703 17627 17729 17653
rect 17729 17627 17730 17653
rect 17702 17626 17730 17627
rect 20118 17150 20146 17178
rect 17598 16869 17626 16870
rect 17598 16843 17599 16869
rect 17599 16843 17625 16869
rect 17625 16843 17626 16869
rect 17598 16842 17626 16843
rect 17650 16869 17678 16870
rect 17650 16843 17651 16869
rect 17651 16843 17677 16869
rect 17677 16843 17678 16869
rect 17650 16842 17678 16843
rect 17702 16869 17730 16870
rect 17702 16843 17703 16869
rect 17703 16843 17729 16869
rect 17729 16843 17730 16869
rect 17702 16842 17730 16843
rect 17598 16085 17626 16086
rect 17598 16059 17599 16085
rect 17599 16059 17625 16085
rect 17625 16059 17626 16085
rect 17598 16058 17626 16059
rect 17650 16085 17678 16086
rect 17650 16059 17651 16085
rect 17651 16059 17677 16085
rect 17677 16059 17678 16085
rect 17650 16058 17678 16059
rect 17702 16085 17730 16086
rect 17702 16059 17703 16085
rect 17703 16059 17729 16085
rect 17729 16059 17730 16085
rect 17702 16058 17730 16059
rect 10822 14014 10850 14042
rect 10374 13846 10402 13874
rect 11158 14041 11186 14042
rect 11158 14015 11159 14041
rect 11159 14015 11185 14041
rect 11185 14015 11186 14041
rect 11158 14014 11186 14015
rect 10990 13985 11018 13986
rect 10990 13959 10991 13985
rect 10991 13959 11017 13985
rect 11017 13959 11018 13985
rect 10990 13958 11018 13959
rect 11438 13873 11466 13874
rect 11438 13847 11439 13873
rect 11439 13847 11465 13873
rect 11465 13847 11466 13873
rect 11438 13846 11466 13847
rect 11942 13846 11970 13874
rect 9534 13342 9562 13370
rect 8470 12558 8498 12586
rect 9086 12558 9114 12586
rect 8974 12417 9002 12418
rect 8974 12391 8975 12417
rect 8975 12391 9001 12417
rect 9001 12391 9002 12417
rect 8974 12390 9002 12391
rect 7630 12278 7658 12306
rect 8246 12334 8274 12362
rect 2238 11381 2266 11382
rect 2238 11355 2239 11381
rect 2239 11355 2265 11381
rect 2265 11355 2266 11381
rect 2238 11354 2266 11355
rect 2290 11381 2318 11382
rect 2290 11355 2291 11381
rect 2291 11355 2317 11381
rect 2317 11355 2318 11381
rect 2290 11354 2318 11355
rect 2342 11381 2370 11382
rect 2342 11355 2343 11381
rect 2343 11355 2369 11381
rect 2369 11355 2370 11381
rect 2342 11354 2370 11355
rect 5390 11326 5418 11354
rect 6454 11241 6482 11242
rect 6454 11215 6455 11241
rect 6455 11215 6481 11241
rect 6481 11215 6482 11241
rect 6454 11214 6482 11215
rect 5054 10934 5082 10962
rect 2238 10597 2266 10598
rect 2238 10571 2239 10597
rect 2239 10571 2265 10597
rect 2265 10571 2266 10597
rect 2238 10570 2266 10571
rect 2290 10597 2318 10598
rect 2290 10571 2291 10597
rect 2291 10571 2317 10597
rect 2317 10571 2318 10597
rect 2290 10570 2318 10571
rect 2342 10597 2370 10598
rect 2342 10571 2343 10597
rect 2343 10571 2369 10597
rect 2369 10571 2370 10597
rect 2342 10570 2370 10571
rect 6958 11326 6986 11354
rect 7070 11214 7098 11242
rect 6790 10934 6818 10962
rect 5390 10598 5418 10626
rect 6566 10598 6594 10626
rect 6454 10457 6482 10458
rect 6454 10431 6455 10457
rect 6455 10431 6481 10457
rect 6481 10431 6482 10457
rect 6454 10430 6482 10431
rect 2086 10262 2114 10290
rect 7294 11214 7322 11242
rect 7574 11774 7602 11802
rect 7518 11577 7546 11578
rect 7518 11551 7519 11577
rect 7519 11551 7545 11577
rect 7545 11551 7546 11577
rect 7518 11550 7546 11551
rect 7574 11550 7602 11578
rect 7462 11326 7490 11354
rect 7350 11102 7378 11130
rect 7462 11073 7490 11074
rect 7462 11047 7463 11073
rect 7463 11047 7489 11073
rect 7489 11047 7490 11073
rect 7462 11046 7490 11047
rect 7518 10905 7546 10906
rect 7518 10879 7519 10905
rect 7519 10879 7545 10905
rect 7545 10879 7546 10905
rect 7518 10878 7546 10879
rect 7238 10542 7266 10570
rect 6846 10457 6874 10458
rect 6846 10431 6847 10457
rect 6847 10431 6873 10457
rect 6873 10431 6874 10457
rect 6846 10430 6874 10431
rect 7126 10430 7154 10458
rect 6902 10401 6930 10402
rect 6902 10375 6903 10401
rect 6903 10375 6929 10401
rect 6929 10375 6930 10401
rect 6902 10374 6930 10375
rect 7630 10737 7658 10738
rect 7630 10711 7631 10737
rect 7631 10711 7657 10737
rect 7657 10711 7658 10737
rect 7630 10710 7658 10711
rect 7574 10598 7602 10626
rect 8918 12361 8946 12362
rect 8918 12335 8919 12361
rect 8919 12335 8945 12361
rect 8945 12335 8946 12361
rect 8918 12334 8946 12335
rect 8246 11886 8274 11914
rect 9422 12502 9450 12530
rect 9366 12417 9394 12418
rect 9366 12391 9367 12417
rect 9367 12391 9393 12417
rect 9393 12391 9394 12417
rect 9366 12390 9394 12391
rect 9142 12361 9170 12362
rect 9142 12335 9143 12361
rect 9143 12335 9169 12361
rect 9169 12335 9170 12361
rect 9142 12334 9170 12335
rect 9086 11886 9114 11914
rect 8694 11774 8722 11802
rect 7854 11577 7882 11578
rect 7854 11551 7855 11577
rect 7855 11551 7881 11577
rect 7881 11551 7882 11577
rect 7854 11550 7882 11551
rect 7910 11102 7938 11130
rect 7910 10990 7938 11018
rect 7686 10486 7714 10514
rect 7742 10878 7770 10906
rect 7406 10318 7434 10346
rect 7518 10401 7546 10402
rect 7518 10375 7519 10401
rect 7519 10375 7545 10401
rect 7545 10375 7546 10401
rect 7518 10374 7546 10375
rect 7854 10094 7882 10122
rect 7742 10009 7770 10010
rect 7742 9983 7743 10009
rect 7743 9983 7769 10009
rect 7769 9983 7770 10009
rect 7742 9982 7770 9983
rect 2238 9813 2266 9814
rect 2238 9787 2239 9813
rect 2239 9787 2265 9813
rect 2265 9787 2266 9813
rect 2238 9786 2266 9787
rect 2290 9813 2318 9814
rect 2290 9787 2291 9813
rect 2291 9787 2317 9813
rect 2317 9787 2318 9813
rect 2290 9786 2318 9787
rect 2342 9813 2370 9814
rect 2342 9787 2343 9813
rect 2343 9787 2369 9813
rect 2369 9787 2370 9813
rect 2342 9786 2370 9787
rect 8022 11046 8050 11074
rect 8414 11577 8442 11578
rect 8414 11551 8415 11577
rect 8415 11551 8441 11577
rect 8441 11551 8442 11577
rect 8414 11550 8442 11551
rect 8134 10542 8162 10570
rect 8302 10710 8330 10738
rect 8246 10486 8274 10514
rect 7966 10345 7994 10346
rect 7966 10319 7967 10345
rect 7967 10319 7993 10345
rect 7993 10319 7994 10345
rect 7966 10318 7994 10319
rect 8078 10009 8106 10010
rect 8078 9983 8079 10009
rect 8079 9983 8105 10009
rect 8105 9983 8106 10009
rect 8078 9982 8106 9983
rect 7966 9926 7994 9954
rect 7742 9534 7770 9562
rect 7630 9478 7658 9506
rect 6230 9225 6258 9226
rect 6230 9199 6231 9225
rect 6231 9199 6257 9225
rect 6257 9199 6258 9225
rect 6230 9198 6258 9199
rect 6062 9142 6090 9170
rect 2238 9029 2266 9030
rect 2238 9003 2239 9029
rect 2239 9003 2265 9029
rect 2265 9003 2266 9029
rect 2238 9002 2266 9003
rect 2290 9029 2318 9030
rect 2290 9003 2291 9029
rect 2291 9003 2317 9029
rect 2317 9003 2318 9029
rect 2290 9002 2318 9003
rect 2342 9029 2370 9030
rect 2342 9003 2343 9029
rect 2343 9003 2369 9029
rect 2369 9003 2370 9029
rect 2342 9002 2370 9003
rect 7014 9142 7042 9170
rect 6454 8750 6482 8778
rect 2238 8245 2266 8246
rect 2238 8219 2239 8245
rect 2239 8219 2265 8245
rect 2265 8219 2266 8245
rect 2238 8218 2266 8219
rect 2290 8245 2318 8246
rect 2290 8219 2291 8245
rect 2291 8219 2317 8245
rect 2317 8219 2318 8245
rect 2290 8218 2318 8219
rect 2342 8245 2370 8246
rect 2342 8219 2343 8245
rect 2343 8219 2369 8245
rect 2369 8219 2370 8245
rect 2342 8218 2370 8219
rect 7574 9169 7602 9170
rect 7574 9143 7575 9169
rect 7575 9143 7601 9169
rect 7601 9143 7602 9169
rect 7574 9142 7602 9143
rect 7518 8638 7546 8666
rect 7518 8470 7546 8498
rect 8134 9534 8162 9562
rect 8190 9758 8218 9786
rect 7966 9030 7994 9058
rect 7742 8750 7770 8778
rect 8078 8638 8106 8666
rect 8526 11073 8554 11074
rect 8526 11047 8527 11073
rect 8527 11047 8553 11073
rect 8553 11047 8554 11073
rect 8526 11046 8554 11047
rect 8806 11830 8834 11858
rect 9590 11662 9618 11690
rect 8862 11577 8890 11578
rect 8862 11551 8863 11577
rect 8863 11551 8889 11577
rect 8889 11551 8890 11577
rect 8862 11550 8890 11551
rect 8414 9758 8442 9786
rect 8470 10710 8498 10738
rect 8302 9702 8330 9730
rect 8302 9534 8330 9562
rect 8582 10486 8610 10514
rect 8526 9590 8554 9618
rect 8414 9478 8442 9506
rect 8414 9254 8442 9282
rect 8414 8694 8442 8722
rect 8806 10654 8834 10682
rect 8918 11102 8946 11130
rect 9478 11185 9506 11186
rect 9478 11159 9479 11185
rect 9479 11159 9505 11185
rect 9505 11159 9506 11185
rect 9478 11158 9506 11159
rect 9086 11046 9114 11074
rect 9254 11073 9282 11074
rect 9254 11047 9255 11073
rect 9255 11047 9281 11073
rect 9281 11047 9282 11073
rect 9254 11046 9282 11047
rect 9478 11046 9506 11074
rect 9030 10710 9058 10738
rect 9030 10542 9058 10570
rect 8750 10374 8778 10402
rect 9142 10430 9170 10458
rect 9142 10318 9170 10346
rect 8862 10289 8890 10290
rect 8862 10263 8863 10289
rect 8863 10263 8889 10289
rect 8889 10263 8890 10289
rect 8862 10262 8890 10263
rect 8806 9982 8834 10010
rect 9422 10654 9450 10682
rect 8974 9617 9002 9618
rect 8974 9591 8975 9617
rect 8975 9591 9001 9617
rect 9001 9591 9002 9617
rect 8974 9590 9002 9591
rect 8862 9561 8890 9562
rect 8862 9535 8863 9561
rect 8863 9535 8889 9561
rect 8889 9535 8890 9561
rect 8862 9534 8890 9535
rect 8806 9478 8834 9506
rect 9086 9505 9114 9506
rect 9086 9479 9087 9505
rect 9087 9479 9113 9505
rect 9113 9479 9114 9505
rect 9086 9478 9114 9479
rect 9310 9590 9338 9618
rect 8694 9254 8722 9282
rect 8638 9142 8666 9170
rect 8582 9086 8610 9114
rect 8358 8553 8386 8554
rect 8358 8527 8359 8553
rect 8359 8527 8385 8553
rect 8385 8527 8386 8553
rect 8358 8526 8386 8527
rect 7966 8470 7994 8498
rect 8302 8497 8330 8498
rect 8302 8471 8303 8497
rect 8303 8471 8329 8497
rect 8329 8471 8330 8497
rect 8302 8470 8330 8471
rect 7742 8441 7770 8442
rect 7742 8415 7743 8441
rect 7743 8415 7769 8441
rect 7769 8415 7770 8441
rect 7742 8414 7770 8415
rect 9254 9281 9282 9282
rect 9254 9255 9255 9281
rect 9255 9255 9281 9281
rect 9281 9255 9282 9281
rect 9254 9254 9282 9255
rect 8862 9086 8890 9114
rect 8862 8777 8890 8778
rect 8862 8751 8863 8777
rect 8863 8751 8889 8777
rect 8889 8751 8890 8777
rect 8862 8750 8890 8751
rect 8750 8694 8778 8722
rect 8582 8638 8610 8666
rect 8918 8358 8946 8386
rect 8526 8134 8554 8162
rect 8862 8161 8890 8162
rect 8862 8135 8863 8161
rect 8863 8135 8889 8161
rect 8889 8135 8890 8161
rect 8862 8134 8890 8135
rect 7350 7601 7378 7602
rect 7350 7575 7351 7601
rect 7351 7575 7377 7601
rect 7377 7575 7378 7601
rect 7350 7574 7378 7575
rect 9142 9086 9170 9114
rect 9198 9142 9226 9170
rect 9086 8694 9114 8722
rect 9142 8862 9170 8890
rect 9030 8526 9058 8554
rect 9198 8721 9226 8722
rect 9198 8695 9199 8721
rect 9199 8695 9225 8721
rect 9225 8695 9226 8721
rect 9198 8694 9226 8695
rect 9918 13341 9946 13342
rect 9918 13315 9919 13341
rect 9919 13315 9945 13341
rect 9945 13315 9946 13341
rect 9918 13314 9946 13315
rect 9970 13341 9998 13342
rect 9970 13315 9971 13341
rect 9971 13315 9997 13341
rect 9997 13315 9998 13341
rect 9970 13314 9998 13315
rect 10022 13341 10050 13342
rect 10022 13315 10023 13341
rect 10023 13315 10049 13341
rect 10049 13315 10050 13341
rect 10022 13314 10050 13315
rect 9814 12614 9842 12642
rect 9918 12557 9946 12558
rect 9918 12531 9919 12557
rect 9919 12531 9945 12557
rect 9945 12531 9946 12557
rect 9918 12530 9946 12531
rect 9970 12557 9998 12558
rect 9970 12531 9971 12557
rect 9971 12531 9997 12557
rect 9997 12531 9998 12557
rect 9970 12530 9998 12531
rect 10022 12557 10050 12558
rect 10022 12531 10023 12557
rect 10023 12531 10049 12557
rect 10049 12531 10050 12557
rect 10022 12530 10050 12531
rect 9758 12390 9786 12418
rect 9758 12278 9786 12306
rect 10318 13174 10346 13202
rect 10094 12166 10122 12194
rect 10150 13145 10178 13146
rect 10150 13119 10151 13145
rect 10151 13119 10177 13145
rect 10177 13119 10178 13145
rect 10150 13118 10178 13119
rect 10598 13481 10626 13482
rect 10598 13455 10599 13481
rect 10599 13455 10625 13481
rect 10625 13455 10626 13481
rect 10598 13454 10626 13455
rect 10710 13566 10738 13594
rect 10766 13174 10794 13202
rect 11214 13118 11242 13146
rect 10318 12614 10346 12642
rect 10766 12614 10794 12642
rect 10150 12334 10178 12362
rect 10094 12054 10122 12082
rect 9982 11830 10010 11858
rect 9918 11773 9946 11774
rect 9918 11747 9919 11773
rect 9919 11747 9945 11773
rect 9945 11747 9946 11773
rect 9918 11746 9946 11747
rect 9970 11773 9998 11774
rect 9970 11747 9971 11773
rect 9971 11747 9997 11773
rect 9997 11747 9998 11773
rect 9970 11746 9998 11747
rect 10022 11773 10050 11774
rect 10022 11747 10023 11773
rect 10023 11747 10049 11773
rect 10049 11747 10050 11773
rect 10022 11746 10050 11747
rect 9758 11494 9786 11522
rect 10598 12390 10626 12418
rect 9646 10990 9674 11018
rect 9758 10990 9786 11018
rect 9702 10878 9730 10906
rect 9646 10793 9674 10794
rect 9646 10767 9647 10793
rect 9647 10767 9673 10793
rect 9673 10767 9674 10793
rect 9646 10766 9674 10767
rect 9534 10038 9562 10066
rect 9366 9030 9394 9058
rect 9422 9478 9450 9506
rect 9366 8526 9394 8554
rect 8974 7657 9002 7658
rect 8974 7631 8975 7657
rect 8975 7631 9001 7657
rect 9001 7631 9002 7657
rect 8974 7630 9002 7631
rect 2238 7461 2266 7462
rect 2238 7435 2239 7461
rect 2239 7435 2265 7461
rect 2265 7435 2266 7461
rect 2238 7434 2266 7435
rect 2290 7461 2318 7462
rect 2290 7435 2291 7461
rect 2291 7435 2317 7461
rect 2317 7435 2318 7461
rect 2290 7434 2318 7435
rect 2342 7461 2370 7462
rect 2342 7435 2343 7461
rect 2343 7435 2369 7461
rect 2369 7435 2370 7461
rect 2342 7434 2370 7435
rect 8302 6929 8330 6930
rect 8302 6903 8303 6929
rect 8303 6903 8329 6929
rect 8329 6903 8330 6929
rect 8302 6902 8330 6903
rect 8414 6873 8442 6874
rect 8414 6847 8415 6873
rect 8415 6847 8441 6873
rect 8441 6847 8442 6873
rect 8414 6846 8442 6847
rect 2238 6677 2266 6678
rect 2238 6651 2239 6677
rect 2239 6651 2265 6677
rect 2265 6651 2266 6677
rect 2238 6650 2266 6651
rect 2290 6677 2318 6678
rect 2290 6651 2291 6677
rect 2291 6651 2317 6677
rect 2317 6651 2318 6677
rect 2290 6650 2318 6651
rect 2342 6677 2370 6678
rect 2342 6651 2343 6677
rect 2343 6651 2369 6677
rect 2369 6651 2370 6677
rect 2342 6650 2370 6651
rect 2238 5893 2266 5894
rect 2238 5867 2239 5893
rect 2239 5867 2265 5893
rect 2265 5867 2266 5893
rect 2238 5866 2266 5867
rect 2290 5893 2318 5894
rect 2290 5867 2291 5893
rect 2291 5867 2317 5893
rect 2317 5867 2318 5893
rect 2290 5866 2318 5867
rect 2342 5893 2370 5894
rect 2342 5867 2343 5893
rect 2343 5867 2369 5893
rect 2369 5867 2370 5893
rect 2342 5866 2370 5867
rect 2238 5109 2266 5110
rect 2238 5083 2239 5109
rect 2239 5083 2265 5109
rect 2265 5083 2266 5109
rect 2238 5082 2266 5083
rect 2290 5109 2318 5110
rect 2290 5083 2291 5109
rect 2291 5083 2317 5109
rect 2317 5083 2318 5109
rect 2290 5082 2318 5083
rect 2342 5109 2370 5110
rect 2342 5083 2343 5109
rect 2343 5083 2369 5109
rect 2369 5083 2370 5109
rect 2342 5082 2370 5083
rect 2238 4325 2266 4326
rect 2238 4299 2239 4325
rect 2239 4299 2265 4325
rect 2265 4299 2266 4325
rect 2238 4298 2266 4299
rect 2290 4325 2318 4326
rect 2290 4299 2291 4325
rect 2291 4299 2317 4325
rect 2317 4299 2318 4325
rect 2290 4298 2318 4299
rect 2342 4325 2370 4326
rect 2342 4299 2343 4325
rect 2343 4299 2369 4325
rect 2369 4299 2370 4325
rect 2342 4298 2370 4299
rect 2238 3541 2266 3542
rect 2238 3515 2239 3541
rect 2239 3515 2265 3541
rect 2265 3515 2266 3541
rect 2238 3514 2266 3515
rect 2290 3541 2318 3542
rect 2290 3515 2291 3541
rect 2291 3515 2317 3541
rect 2317 3515 2318 3541
rect 2290 3514 2318 3515
rect 2342 3541 2370 3542
rect 2342 3515 2343 3541
rect 2343 3515 2369 3541
rect 2369 3515 2370 3541
rect 2342 3514 2370 3515
rect 2238 2757 2266 2758
rect 2238 2731 2239 2757
rect 2239 2731 2265 2757
rect 2265 2731 2266 2757
rect 2238 2730 2266 2731
rect 2290 2757 2318 2758
rect 2290 2731 2291 2757
rect 2291 2731 2317 2757
rect 2317 2731 2318 2757
rect 2290 2730 2318 2731
rect 2342 2757 2370 2758
rect 2342 2731 2343 2757
rect 2343 2731 2369 2757
rect 2369 2731 2370 2757
rect 2342 2730 2370 2731
rect 8918 7601 8946 7602
rect 8918 7575 8919 7601
rect 8919 7575 8945 7601
rect 8945 7575 8946 7601
rect 8918 7574 8946 7575
rect 8694 6734 8722 6762
rect 9646 10262 9674 10290
rect 9590 9422 9618 9450
rect 9534 9254 9562 9282
rect 9534 9030 9562 9058
rect 9310 8134 9338 8162
rect 9646 8889 9674 8890
rect 9646 8863 9647 8889
rect 9647 8863 9673 8889
rect 9673 8863 9674 8889
rect 9646 8862 9674 8863
rect 10038 11073 10066 11074
rect 10038 11047 10039 11073
rect 10039 11047 10065 11073
rect 10065 11047 10066 11073
rect 10038 11046 10066 11047
rect 10150 11073 10178 11074
rect 10150 11047 10151 11073
rect 10151 11047 10177 11073
rect 10177 11047 10178 11073
rect 10150 11046 10178 11047
rect 9918 10989 9946 10990
rect 9918 10963 9919 10989
rect 9919 10963 9945 10989
rect 9945 10963 9946 10989
rect 9918 10962 9946 10963
rect 9970 10989 9998 10990
rect 9970 10963 9971 10989
rect 9971 10963 9997 10989
rect 9997 10963 9998 10989
rect 9970 10962 9998 10963
rect 10022 10989 10050 10990
rect 10022 10963 10023 10989
rect 10023 10963 10049 10989
rect 10049 10963 10050 10989
rect 10022 10962 10050 10963
rect 10150 10878 10178 10906
rect 9814 10681 9842 10682
rect 9814 10655 9815 10681
rect 9815 10655 9841 10681
rect 9841 10655 9842 10681
rect 9814 10654 9842 10655
rect 9422 8049 9450 8050
rect 9422 8023 9423 8049
rect 9423 8023 9449 8049
rect 9449 8023 9450 8049
rect 9422 8022 9450 8023
rect 9254 7630 9282 7658
rect 9142 7601 9170 7602
rect 9142 7575 9143 7601
rect 9143 7575 9169 7601
rect 9169 7575 9170 7601
rect 9142 7574 9170 7575
rect 9702 7686 9730 7714
rect 9758 7910 9786 7938
rect 10094 10401 10122 10402
rect 10094 10375 10095 10401
rect 10095 10375 10121 10401
rect 10121 10375 10122 10401
rect 10094 10374 10122 10375
rect 9982 10345 10010 10346
rect 9982 10319 9983 10345
rect 9983 10319 10009 10345
rect 10009 10319 10010 10345
rect 9982 10318 10010 10319
rect 9918 10205 9946 10206
rect 9918 10179 9919 10205
rect 9919 10179 9945 10205
rect 9945 10179 9946 10205
rect 9918 10178 9946 10179
rect 9970 10205 9998 10206
rect 9970 10179 9971 10205
rect 9971 10179 9997 10205
rect 9997 10179 9998 10205
rect 9970 10178 9998 10179
rect 10022 10205 10050 10206
rect 10022 10179 10023 10205
rect 10023 10179 10049 10205
rect 10049 10179 10050 10205
rect 10022 10178 10050 10179
rect 10430 11886 10458 11914
rect 10430 11633 10458 11634
rect 10430 11607 10431 11633
rect 10431 11607 10457 11633
rect 10457 11607 10458 11633
rect 10430 11606 10458 11607
rect 10262 11129 10290 11130
rect 10262 11103 10263 11129
rect 10263 11103 10289 11129
rect 10289 11103 10290 11129
rect 10262 11102 10290 11103
rect 10654 12278 10682 12306
rect 10878 12670 10906 12698
rect 10654 11158 10682 11186
rect 10710 11046 10738 11074
rect 10598 10990 10626 11018
rect 10710 10878 10738 10906
rect 10374 10710 10402 10738
rect 10206 10401 10234 10402
rect 10206 10375 10207 10401
rect 10207 10375 10233 10401
rect 10233 10375 10234 10401
rect 10206 10374 10234 10375
rect 10150 10065 10178 10066
rect 10150 10039 10151 10065
rect 10151 10039 10177 10065
rect 10177 10039 10178 10065
rect 10150 10038 10178 10039
rect 10094 9982 10122 10010
rect 10374 10262 10402 10290
rect 10206 9926 10234 9954
rect 10206 9814 10234 9842
rect 10094 9758 10122 9786
rect 10206 9646 10234 9674
rect 9918 9421 9946 9422
rect 9918 9395 9919 9421
rect 9919 9395 9945 9421
rect 9945 9395 9946 9421
rect 9918 9394 9946 9395
rect 9970 9421 9998 9422
rect 9970 9395 9971 9421
rect 9971 9395 9997 9421
rect 9997 9395 9998 9421
rect 9970 9394 9998 9395
rect 10022 9421 10050 9422
rect 10022 9395 10023 9421
rect 10023 9395 10049 9421
rect 10049 9395 10050 9421
rect 10022 9394 10050 9395
rect 9870 9310 9898 9338
rect 10094 9142 10122 9170
rect 9870 8777 9898 8778
rect 9870 8751 9871 8777
rect 9871 8751 9897 8777
rect 9897 8751 9898 8777
rect 9870 8750 9898 8751
rect 9918 8637 9946 8638
rect 9918 8611 9919 8637
rect 9919 8611 9945 8637
rect 9945 8611 9946 8637
rect 9918 8610 9946 8611
rect 9970 8637 9998 8638
rect 9970 8611 9971 8637
rect 9971 8611 9997 8637
rect 9997 8611 9998 8637
rect 9970 8610 9998 8611
rect 10022 8637 10050 8638
rect 10022 8611 10023 8637
rect 10023 8611 10049 8637
rect 10049 8611 10050 8637
rect 10022 8610 10050 8611
rect 10038 8526 10066 8554
rect 10374 9646 10402 9674
rect 10374 9534 10402 9562
rect 10318 9505 10346 9506
rect 10318 9479 10319 9505
rect 10319 9479 10345 9505
rect 10345 9479 10346 9505
rect 10318 9478 10346 9479
rect 10710 10542 10738 10570
rect 10878 11830 10906 11858
rect 17598 15301 17626 15302
rect 17598 15275 17599 15301
rect 17599 15275 17625 15301
rect 17625 15275 17626 15301
rect 17598 15274 17626 15275
rect 17650 15301 17678 15302
rect 17650 15275 17651 15301
rect 17651 15275 17677 15301
rect 17677 15275 17678 15301
rect 17650 15274 17678 15275
rect 17702 15301 17730 15302
rect 17702 15275 17703 15301
rect 17703 15275 17729 15301
rect 17729 15275 17730 15301
rect 17702 15274 17730 15275
rect 17598 14517 17626 14518
rect 17598 14491 17599 14517
rect 17599 14491 17625 14517
rect 17625 14491 17626 14517
rect 17598 14490 17626 14491
rect 17650 14517 17678 14518
rect 17650 14491 17651 14517
rect 17651 14491 17677 14517
rect 17677 14491 17678 14517
rect 17650 14490 17678 14491
rect 17702 14517 17730 14518
rect 17702 14491 17703 14517
rect 17703 14491 17729 14517
rect 17729 14491 17730 14517
rect 17702 14490 17730 14491
rect 17598 13733 17626 13734
rect 17598 13707 17599 13733
rect 17599 13707 17625 13733
rect 17625 13707 17626 13733
rect 17598 13706 17626 13707
rect 17650 13733 17678 13734
rect 17650 13707 17651 13733
rect 17651 13707 17677 13733
rect 17677 13707 17678 13733
rect 17650 13706 17678 13707
rect 17702 13733 17730 13734
rect 17702 13707 17703 13733
rect 17703 13707 17729 13733
rect 17729 13707 17730 13733
rect 17702 13706 17730 13707
rect 13454 13537 13482 13538
rect 13454 13511 13455 13537
rect 13455 13511 13481 13537
rect 13481 13511 13482 13537
rect 13454 13510 13482 13511
rect 14238 13510 14266 13538
rect 12222 13454 12250 13482
rect 11942 13062 11970 13090
rect 11494 12753 11522 12754
rect 11494 12727 11495 12753
rect 11495 12727 11521 12753
rect 11521 12727 11522 12753
rect 11494 12726 11522 12727
rect 11326 12670 11354 12698
rect 12110 12726 12138 12754
rect 13398 13481 13426 13482
rect 13398 13455 13399 13481
rect 13399 13455 13425 13481
rect 13425 13455 13426 13481
rect 13398 13454 13426 13455
rect 12278 13174 12306 13202
rect 18830 13537 18858 13538
rect 18830 13511 18831 13537
rect 18831 13511 18857 13537
rect 18857 13511 18858 13537
rect 18830 13510 18858 13511
rect 12334 13089 12362 13090
rect 12334 13063 12335 13089
rect 12335 13063 12361 13089
rect 12361 13063 12362 13089
rect 12334 13062 12362 13063
rect 12502 12809 12530 12810
rect 12502 12783 12503 12809
rect 12503 12783 12529 12809
rect 12529 12783 12530 12809
rect 12502 12782 12530 12783
rect 11718 12166 11746 12194
rect 11662 11969 11690 11970
rect 11662 11943 11663 11969
rect 11663 11943 11689 11969
rect 11689 11943 11690 11969
rect 11662 11942 11690 11943
rect 11270 11857 11298 11858
rect 11270 11831 11271 11857
rect 11271 11831 11297 11857
rect 11297 11831 11298 11857
rect 11270 11830 11298 11831
rect 10934 11718 10962 11746
rect 10934 11606 10962 11634
rect 10878 11102 10906 11130
rect 11494 11326 11522 11354
rect 10878 10822 10906 10850
rect 11606 11046 11634 11074
rect 11606 10822 11634 10850
rect 10934 10793 10962 10794
rect 10934 10767 10935 10793
rect 10935 10767 10961 10793
rect 10961 10767 10962 10793
rect 10934 10766 10962 10767
rect 11214 10598 11242 10626
rect 11158 10430 11186 10458
rect 11046 10401 11074 10402
rect 11046 10375 11047 10401
rect 11047 10375 11073 10401
rect 11073 10375 11074 10401
rect 11046 10374 11074 10375
rect 10766 10289 10794 10290
rect 10766 10263 10767 10289
rect 10767 10263 10793 10289
rect 10793 10263 10794 10289
rect 10766 10262 10794 10263
rect 10654 9646 10682 9674
rect 10710 9702 10738 9730
rect 10598 9590 10626 9618
rect 10542 9366 10570 9394
rect 10654 9534 10682 9562
rect 10262 8078 10290 8106
rect 9982 7937 10010 7938
rect 9982 7911 9983 7937
rect 9983 7911 10009 7937
rect 10009 7911 10010 7937
rect 9982 7910 10010 7911
rect 9918 7853 9946 7854
rect 9918 7827 9919 7853
rect 9919 7827 9945 7853
rect 9945 7827 9946 7853
rect 9918 7826 9946 7827
rect 9970 7853 9998 7854
rect 9970 7827 9971 7853
rect 9971 7827 9997 7853
rect 9997 7827 9998 7853
rect 9970 7826 9998 7827
rect 10022 7853 10050 7854
rect 10022 7827 10023 7853
rect 10023 7827 10049 7853
rect 10049 7827 10050 7853
rect 10022 7826 10050 7827
rect 9814 7657 9842 7658
rect 9814 7631 9815 7657
rect 9815 7631 9841 7657
rect 9841 7631 9842 7657
rect 9814 7630 9842 7631
rect 9142 6902 9170 6930
rect 9310 6902 9338 6930
rect 9030 6790 9058 6818
rect 9534 7238 9562 7266
rect 10430 8526 10458 8554
rect 10150 7993 10178 7994
rect 10150 7967 10151 7993
rect 10151 7967 10177 7993
rect 10177 7967 10178 7993
rect 10150 7966 10178 7967
rect 11270 10486 11298 10514
rect 11494 10710 11522 10738
rect 11382 10430 11410 10458
rect 11214 10345 11242 10346
rect 11214 10319 11215 10345
rect 11215 10319 11241 10345
rect 11241 10319 11242 10345
rect 11214 10318 11242 10319
rect 11382 10094 11410 10122
rect 11326 10038 11354 10066
rect 10934 9561 10962 9562
rect 10934 9535 10935 9561
rect 10935 9535 10961 9561
rect 10961 9535 10962 9561
rect 10934 9534 10962 9535
rect 11046 9086 11074 9114
rect 11158 9310 11186 9338
rect 10822 9030 10850 9058
rect 11326 9366 11354 9394
rect 10710 8777 10738 8778
rect 10710 8751 10711 8777
rect 10711 8751 10737 8777
rect 10737 8751 10738 8777
rect 10710 8750 10738 8751
rect 11382 9478 11410 9506
rect 11494 10374 11522 10402
rect 12110 12641 12138 12642
rect 12110 12615 12111 12641
rect 12111 12615 12137 12641
rect 12137 12615 12138 12641
rect 12110 12614 12138 12615
rect 19950 13398 19978 13426
rect 14406 13201 14434 13202
rect 14406 13175 14407 13201
rect 14407 13175 14433 13201
rect 14433 13175 14434 13201
rect 14406 13174 14434 13175
rect 18830 13145 18858 13146
rect 18830 13119 18831 13145
rect 18831 13119 18857 13145
rect 18857 13119 18858 13145
rect 18830 13118 18858 13119
rect 20006 13118 20034 13146
rect 17598 12949 17626 12950
rect 17598 12923 17599 12949
rect 17599 12923 17625 12949
rect 17625 12923 17626 12949
rect 17598 12922 17626 12923
rect 17650 12949 17678 12950
rect 17650 12923 17651 12949
rect 17651 12923 17677 12949
rect 17677 12923 17678 12949
rect 17650 12922 17678 12923
rect 17702 12949 17730 12950
rect 17702 12923 17703 12949
rect 17703 12923 17729 12949
rect 17729 12923 17730 12949
rect 17702 12922 17730 12923
rect 13006 12782 13034 12810
rect 13678 12726 13706 12754
rect 12446 12446 12474 12474
rect 12726 12614 12754 12642
rect 12950 12446 12978 12474
rect 12838 12417 12866 12418
rect 12838 12391 12839 12417
rect 12839 12391 12865 12417
rect 12865 12391 12866 12417
rect 12838 12390 12866 12391
rect 12838 12278 12866 12306
rect 13622 12417 13650 12418
rect 13622 12391 13623 12417
rect 13623 12391 13649 12417
rect 13649 12391 13650 12417
rect 13622 12390 13650 12391
rect 14126 12726 14154 12754
rect 18830 12753 18858 12754
rect 18830 12727 18831 12753
rect 18831 12727 18857 12753
rect 18857 12727 18858 12753
rect 18830 12726 18858 12727
rect 20006 12446 20034 12474
rect 17598 12165 17626 12166
rect 17598 12139 17599 12165
rect 17599 12139 17625 12165
rect 17625 12139 17626 12165
rect 17598 12138 17626 12139
rect 17650 12165 17678 12166
rect 17650 12139 17651 12165
rect 17651 12139 17677 12165
rect 17677 12139 17678 12165
rect 17650 12138 17678 12139
rect 17702 12165 17730 12166
rect 17702 12139 17703 12165
rect 17703 12139 17729 12165
rect 17729 12139 17730 12165
rect 17702 12138 17730 12139
rect 12894 11942 12922 11970
rect 11942 11606 11970 11634
rect 12558 11606 12586 11634
rect 11998 11326 12026 11354
rect 11718 10878 11746 10906
rect 11718 10710 11746 10738
rect 12334 11270 12362 11298
rect 11942 10793 11970 10794
rect 11942 10767 11943 10793
rect 11943 10767 11969 10793
rect 11969 10767 11970 10793
rect 11942 10766 11970 10767
rect 11886 10318 11914 10346
rect 12110 10849 12138 10850
rect 12110 10823 12111 10849
rect 12111 10823 12137 10849
rect 12137 10823 12138 10849
rect 12110 10822 12138 10823
rect 12558 11158 12586 11186
rect 12894 11185 12922 11186
rect 12894 11159 12895 11185
rect 12895 11159 12921 11185
rect 12921 11159 12922 11185
rect 12894 11158 12922 11159
rect 12054 10654 12082 10682
rect 13510 10878 13538 10906
rect 13622 11158 13650 11186
rect 17598 11381 17626 11382
rect 17598 11355 17599 11381
rect 17599 11355 17625 11381
rect 17625 11355 17626 11381
rect 17598 11354 17626 11355
rect 17650 11381 17678 11382
rect 17650 11355 17651 11381
rect 17651 11355 17677 11381
rect 17677 11355 17678 11381
rect 17650 11354 17678 11355
rect 17702 11381 17730 11382
rect 17702 11355 17703 11381
rect 17703 11355 17729 11381
rect 17729 11355 17730 11381
rect 17702 11354 17730 11355
rect 20006 11465 20034 11466
rect 20006 11439 20007 11465
rect 20007 11439 20033 11465
rect 20033 11439 20034 11465
rect 20006 11438 20034 11439
rect 18830 11270 18858 11298
rect 14294 11158 14322 11186
rect 18830 11185 18858 11186
rect 18830 11159 18831 11185
rect 18831 11159 18857 11185
rect 18857 11159 18858 11185
rect 18830 11158 18858 11159
rect 20006 11102 20034 11130
rect 12110 10345 12138 10346
rect 12110 10319 12111 10345
rect 12111 10319 12137 10345
rect 12137 10319 12138 10345
rect 12110 10318 12138 10319
rect 11942 10038 11970 10066
rect 11942 9953 11970 9954
rect 11942 9927 11943 9953
rect 11943 9927 11969 9953
rect 11969 9927 11970 9953
rect 11942 9926 11970 9927
rect 11438 9225 11466 9226
rect 11438 9199 11439 9225
rect 11439 9199 11465 9225
rect 11465 9199 11466 9225
rect 11438 9198 11466 9199
rect 11662 9534 11690 9562
rect 11774 9590 11802 9618
rect 12110 9617 12138 9618
rect 12110 9591 12111 9617
rect 12111 9591 12137 9617
rect 12137 9591 12138 9617
rect 12110 9590 12138 9591
rect 11998 9505 12026 9506
rect 11998 9479 11999 9505
rect 11999 9479 12025 9505
rect 12025 9479 12026 9505
rect 11998 9478 12026 9479
rect 11550 9086 11578 9114
rect 10934 8414 10962 8442
rect 10766 8078 10794 8106
rect 10878 7937 10906 7938
rect 10878 7911 10879 7937
rect 10879 7911 10905 7937
rect 10905 7911 10906 7937
rect 10878 7910 10906 7911
rect 10150 7574 10178 7602
rect 10990 8049 11018 8050
rect 10990 8023 10991 8049
rect 10991 8023 11017 8049
rect 11017 8023 11018 8049
rect 10990 8022 11018 8023
rect 10766 7294 10794 7322
rect 12894 10009 12922 10010
rect 12894 9983 12895 10009
rect 12895 9983 12921 10009
rect 12921 9983 12922 10009
rect 12894 9982 12922 9983
rect 12782 9953 12810 9954
rect 12782 9927 12783 9953
rect 12783 9927 12809 9953
rect 12809 9927 12810 9953
rect 12782 9926 12810 9927
rect 13230 10009 13258 10010
rect 13230 9983 13231 10009
rect 13231 9983 13257 10009
rect 13257 9983 13258 10009
rect 13230 9982 13258 9983
rect 13006 9926 13034 9954
rect 13062 9870 13090 9898
rect 12894 9617 12922 9618
rect 12894 9591 12895 9617
rect 12895 9591 12921 9617
rect 12921 9591 12922 9617
rect 12894 9590 12922 9591
rect 12390 9561 12418 9562
rect 12390 9535 12391 9561
rect 12391 9535 12417 9561
rect 12417 9535 12418 9561
rect 12390 9534 12418 9535
rect 12558 9505 12586 9506
rect 12558 9479 12559 9505
rect 12559 9479 12585 9505
rect 12585 9479 12586 9505
rect 12558 9478 12586 9479
rect 12166 8022 12194 8050
rect 13678 10766 13706 10794
rect 17598 10597 17626 10598
rect 17598 10571 17599 10597
rect 17599 10571 17625 10597
rect 17625 10571 17626 10597
rect 17598 10570 17626 10571
rect 17650 10597 17678 10598
rect 17650 10571 17651 10597
rect 17651 10571 17677 10597
rect 17677 10571 17678 10597
rect 17650 10570 17678 10571
rect 17702 10597 17730 10598
rect 17702 10571 17703 10597
rect 17703 10571 17729 10597
rect 17729 10571 17730 10597
rect 17702 10570 17730 10571
rect 13790 10318 13818 10346
rect 14294 10318 14322 10346
rect 14630 10318 14658 10346
rect 19950 10430 19978 10458
rect 18830 10401 18858 10402
rect 18830 10375 18831 10401
rect 18831 10375 18857 10401
rect 18857 10375 18858 10401
rect 18830 10374 18858 10375
rect 18718 10318 18746 10346
rect 14742 10289 14770 10290
rect 14742 10263 14743 10289
rect 14743 10263 14769 10289
rect 14769 10263 14770 10289
rect 14742 10262 14770 10263
rect 20006 10094 20034 10122
rect 13622 9953 13650 9954
rect 13622 9927 13623 9953
rect 13623 9927 13649 9953
rect 13649 9927 13650 9953
rect 13622 9926 13650 9927
rect 13342 9870 13370 9898
rect 13118 9561 13146 9562
rect 13118 9535 13119 9561
rect 13119 9535 13145 9561
rect 13145 9535 13146 9561
rect 13118 9534 13146 9535
rect 13678 9590 13706 9618
rect 13566 9561 13594 9562
rect 13566 9535 13567 9561
rect 13567 9535 13593 9561
rect 13593 9535 13594 9561
rect 13566 9534 13594 9535
rect 17598 9813 17626 9814
rect 17598 9787 17599 9813
rect 17599 9787 17625 9813
rect 17625 9787 17626 9813
rect 17598 9786 17626 9787
rect 17650 9813 17678 9814
rect 17650 9787 17651 9813
rect 17651 9787 17677 9813
rect 17677 9787 17678 9813
rect 17650 9786 17678 9787
rect 17702 9813 17730 9814
rect 17702 9787 17703 9813
rect 17703 9787 17729 9813
rect 17729 9787 17730 9813
rect 17702 9786 17730 9787
rect 13734 9478 13762 9506
rect 13622 8833 13650 8834
rect 13622 8807 13623 8833
rect 13623 8807 13649 8833
rect 13649 8807 13650 8833
rect 13622 8806 13650 8807
rect 13510 8414 13538 8442
rect 14294 9590 14322 9618
rect 18830 9617 18858 9618
rect 18830 9591 18831 9617
rect 18831 9591 18857 9617
rect 18857 9591 18858 9617
rect 18830 9590 18858 9591
rect 20006 9422 20034 9450
rect 17598 9029 17626 9030
rect 17598 9003 17599 9029
rect 17599 9003 17625 9029
rect 17625 9003 17626 9029
rect 17598 9002 17626 9003
rect 17650 9029 17678 9030
rect 17650 9003 17651 9029
rect 17651 9003 17677 9029
rect 17677 9003 17678 9029
rect 17650 9002 17678 9003
rect 17702 9029 17730 9030
rect 17702 9003 17703 9029
rect 17703 9003 17729 9029
rect 17729 9003 17730 9029
rect 17702 9002 17730 9003
rect 11830 7966 11858 7994
rect 11886 7910 11914 7938
rect 10262 7265 10290 7266
rect 10262 7239 10263 7265
rect 10263 7239 10289 7265
rect 10289 7239 10290 7265
rect 10262 7238 10290 7239
rect 10374 7265 10402 7266
rect 10374 7239 10375 7265
rect 10375 7239 10401 7265
rect 10401 7239 10402 7265
rect 10374 7238 10402 7239
rect 10934 7518 10962 7546
rect 11158 7321 11186 7322
rect 11158 7295 11159 7321
rect 11159 7295 11185 7321
rect 11185 7295 11186 7321
rect 11158 7294 11186 7295
rect 9918 7069 9946 7070
rect 9918 7043 9919 7069
rect 9919 7043 9945 7069
rect 9945 7043 9946 7069
rect 9918 7042 9946 7043
rect 9970 7069 9998 7070
rect 9970 7043 9971 7069
rect 9971 7043 9997 7069
rect 9997 7043 9998 7069
rect 9970 7042 9998 7043
rect 10022 7069 10050 7070
rect 10022 7043 10023 7069
rect 10023 7043 10049 7069
rect 10049 7043 10050 7069
rect 10022 7042 10050 7043
rect 9646 6873 9674 6874
rect 9646 6847 9647 6873
rect 9647 6847 9673 6873
rect 9673 6847 9674 6873
rect 9646 6846 9674 6847
rect 9758 6873 9786 6874
rect 9758 6847 9759 6873
rect 9759 6847 9785 6873
rect 9785 6847 9786 6873
rect 9758 6846 9786 6847
rect 10038 6873 10066 6874
rect 10038 6847 10039 6873
rect 10039 6847 10065 6873
rect 10065 6847 10066 6873
rect 10038 6846 10066 6847
rect 9870 6817 9898 6818
rect 9870 6791 9871 6817
rect 9871 6791 9897 6817
rect 9897 6791 9898 6817
rect 9870 6790 9898 6791
rect 10206 6929 10234 6930
rect 10206 6903 10207 6929
rect 10207 6903 10233 6929
rect 10233 6903 10234 6929
rect 10206 6902 10234 6903
rect 10318 6734 10346 6762
rect 8750 2030 8778 2058
rect 2238 1973 2266 1974
rect 2238 1947 2239 1973
rect 2239 1947 2265 1973
rect 2265 1947 2266 1973
rect 2238 1946 2266 1947
rect 2290 1973 2318 1974
rect 2290 1947 2291 1973
rect 2291 1947 2317 1973
rect 2317 1947 2318 1973
rect 2290 1946 2318 1947
rect 2342 1973 2370 1974
rect 2342 1947 2343 1973
rect 2343 1947 2369 1973
rect 2369 1947 2370 1973
rect 2342 1946 2370 1947
rect 9918 6285 9946 6286
rect 9918 6259 9919 6285
rect 9919 6259 9945 6285
rect 9945 6259 9946 6285
rect 9918 6258 9946 6259
rect 9970 6285 9998 6286
rect 9970 6259 9971 6285
rect 9971 6259 9997 6285
rect 9997 6259 9998 6285
rect 9970 6258 9998 6259
rect 10022 6285 10050 6286
rect 10022 6259 10023 6285
rect 10023 6259 10049 6285
rect 10049 6259 10050 6285
rect 10022 6258 10050 6259
rect 9918 5501 9946 5502
rect 9918 5475 9919 5501
rect 9919 5475 9945 5501
rect 9945 5475 9946 5501
rect 9918 5474 9946 5475
rect 9970 5501 9998 5502
rect 9970 5475 9971 5501
rect 9971 5475 9997 5501
rect 9997 5475 9998 5501
rect 9970 5474 9998 5475
rect 10022 5501 10050 5502
rect 10022 5475 10023 5501
rect 10023 5475 10049 5501
rect 10049 5475 10050 5501
rect 10022 5474 10050 5475
rect 9918 4717 9946 4718
rect 9918 4691 9919 4717
rect 9919 4691 9945 4717
rect 9945 4691 9946 4717
rect 9918 4690 9946 4691
rect 9970 4717 9998 4718
rect 9970 4691 9971 4717
rect 9971 4691 9997 4717
rect 9997 4691 9998 4717
rect 9970 4690 9998 4691
rect 10022 4717 10050 4718
rect 10022 4691 10023 4717
rect 10023 4691 10049 4717
rect 10049 4691 10050 4717
rect 10022 4690 10050 4691
rect 9918 3933 9946 3934
rect 9918 3907 9919 3933
rect 9919 3907 9945 3933
rect 9945 3907 9946 3933
rect 9918 3906 9946 3907
rect 9970 3933 9998 3934
rect 9970 3907 9971 3933
rect 9971 3907 9997 3933
rect 9997 3907 9998 3933
rect 9970 3906 9998 3907
rect 10022 3933 10050 3934
rect 10022 3907 10023 3933
rect 10023 3907 10049 3933
rect 10049 3907 10050 3933
rect 10022 3906 10050 3907
rect 9918 3149 9946 3150
rect 9918 3123 9919 3149
rect 9919 3123 9945 3149
rect 9945 3123 9946 3149
rect 9918 3122 9946 3123
rect 9970 3149 9998 3150
rect 9970 3123 9971 3149
rect 9971 3123 9997 3149
rect 9997 3123 9998 3149
rect 9970 3122 9998 3123
rect 10022 3149 10050 3150
rect 10022 3123 10023 3149
rect 10023 3123 10049 3149
rect 10049 3123 10050 3149
rect 10022 3122 10050 3123
rect 9918 2365 9946 2366
rect 9918 2339 9919 2365
rect 9919 2339 9945 2365
rect 9945 2339 9946 2365
rect 9918 2338 9946 2339
rect 9970 2365 9998 2366
rect 9970 2339 9971 2365
rect 9971 2339 9997 2365
rect 9997 2339 9998 2365
rect 9970 2338 9998 2339
rect 10022 2365 10050 2366
rect 10022 2339 10023 2365
rect 10023 2339 10049 2365
rect 10049 2339 10050 2365
rect 10022 2338 10050 2339
rect 9366 2057 9394 2058
rect 9366 2031 9367 2057
rect 9367 2031 9393 2057
rect 9393 2031 9394 2057
rect 9366 2030 9394 2031
rect 11830 7518 11858 7546
rect 11270 7238 11298 7266
rect 11214 6873 11242 6874
rect 11214 6847 11215 6873
rect 11215 6847 11241 6873
rect 11241 6847 11242 6873
rect 11214 6846 11242 6847
rect 12950 8302 12978 8330
rect 13062 8049 13090 8050
rect 13062 8023 13063 8049
rect 13063 8023 13089 8049
rect 13089 8023 13090 8049
rect 13062 8022 13090 8023
rect 14294 8806 14322 8834
rect 18830 8833 18858 8834
rect 18830 8807 18831 8833
rect 18831 8807 18857 8833
rect 18857 8807 18858 8833
rect 18830 8806 18858 8807
rect 20006 8750 20034 8778
rect 17598 8245 17626 8246
rect 17598 8219 17599 8245
rect 17599 8219 17625 8245
rect 17625 8219 17626 8245
rect 17598 8218 17626 8219
rect 17650 8245 17678 8246
rect 17650 8219 17651 8245
rect 17651 8219 17677 8245
rect 17677 8219 17678 8245
rect 17650 8218 17678 8219
rect 17702 8245 17730 8246
rect 17702 8219 17703 8245
rect 17703 8219 17729 8245
rect 17729 8219 17730 8245
rect 17702 8218 17730 8219
rect 12950 7993 12978 7994
rect 12950 7967 12951 7993
rect 12951 7967 12977 7993
rect 12977 7967 12978 7993
rect 12950 7966 12978 7967
rect 12334 7518 12362 7546
rect 13566 7574 13594 7602
rect 14238 7601 14266 7602
rect 14238 7575 14239 7601
rect 14239 7575 14265 7601
rect 14265 7575 14266 7601
rect 14238 7574 14266 7575
rect 20006 7742 20034 7770
rect 18830 7574 18858 7602
rect 17598 7461 17626 7462
rect 17598 7435 17599 7461
rect 17599 7435 17625 7461
rect 17625 7435 17626 7461
rect 17598 7434 17626 7435
rect 17650 7461 17678 7462
rect 17650 7435 17651 7461
rect 17651 7435 17677 7461
rect 17677 7435 17678 7461
rect 17650 7434 17678 7435
rect 17702 7461 17730 7462
rect 17702 7435 17703 7461
rect 17703 7435 17729 7461
rect 17729 7435 17730 7461
rect 17702 7434 17730 7435
rect 12894 7153 12922 7154
rect 12894 7127 12895 7153
rect 12895 7127 12921 7153
rect 12921 7127 12922 7153
rect 12894 7126 12922 7127
rect 13454 7126 13482 7154
rect 12614 6873 12642 6874
rect 12614 6847 12615 6873
rect 12615 6847 12641 6873
rect 12641 6847 12642 6873
rect 12614 6846 12642 6847
rect 12222 6734 12250 6762
rect 12670 6734 12698 6762
rect 11382 5894 11410 5922
rect 11662 5894 11690 5922
rect 12278 5894 12306 5922
rect 12110 2030 12138 2058
rect 11438 1806 11466 1834
rect 10094 1694 10122 1722
rect 9918 1581 9946 1582
rect 9918 1555 9919 1581
rect 9919 1555 9945 1581
rect 9945 1555 9946 1581
rect 9918 1554 9946 1555
rect 9970 1581 9998 1582
rect 9970 1555 9971 1581
rect 9971 1555 9997 1581
rect 9997 1555 9998 1581
rect 9970 1554 9998 1555
rect 10022 1581 10050 1582
rect 10022 1555 10023 1581
rect 10023 1555 10049 1581
rect 10049 1555 10050 1581
rect 10022 1554 10050 1555
rect 10878 1694 10906 1722
rect 17598 6677 17626 6678
rect 17598 6651 17599 6677
rect 17599 6651 17625 6677
rect 17625 6651 17626 6677
rect 17598 6650 17626 6651
rect 17650 6677 17678 6678
rect 17650 6651 17651 6677
rect 17651 6651 17677 6677
rect 17677 6651 17678 6677
rect 17650 6650 17678 6651
rect 17702 6677 17730 6678
rect 17702 6651 17703 6677
rect 17703 6651 17729 6677
rect 17729 6651 17730 6677
rect 17702 6650 17730 6651
rect 13454 6537 13482 6538
rect 13454 6511 13455 6537
rect 13455 6511 13481 6537
rect 13481 6511 13482 6537
rect 13454 6510 13482 6511
rect 14294 6510 14322 6538
rect 13118 2057 13146 2058
rect 13118 2031 13119 2057
rect 13119 2031 13145 2057
rect 13145 2031 13146 2057
rect 13118 2030 13146 2031
rect 12782 1833 12810 1834
rect 12782 1807 12783 1833
rect 12783 1807 12809 1833
rect 12809 1807 12810 1833
rect 12782 1806 12810 1807
rect 13174 1806 13202 1834
rect 17598 5893 17626 5894
rect 17598 5867 17599 5893
rect 17599 5867 17625 5893
rect 17625 5867 17626 5893
rect 17598 5866 17626 5867
rect 17650 5893 17678 5894
rect 17650 5867 17651 5893
rect 17651 5867 17677 5893
rect 17677 5867 17678 5893
rect 17650 5866 17678 5867
rect 17702 5893 17730 5894
rect 17702 5867 17703 5893
rect 17703 5867 17729 5893
rect 17729 5867 17730 5893
rect 17702 5866 17730 5867
rect 17598 5109 17626 5110
rect 17598 5083 17599 5109
rect 17599 5083 17625 5109
rect 17625 5083 17626 5109
rect 17598 5082 17626 5083
rect 17650 5109 17678 5110
rect 17650 5083 17651 5109
rect 17651 5083 17677 5109
rect 17677 5083 17678 5109
rect 17650 5082 17678 5083
rect 17702 5109 17730 5110
rect 17702 5083 17703 5109
rect 17703 5083 17729 5109
rect 17729 5083 17730 5109
rect 17702 5082 17730 5083
rect 17598 4325 17626 4326
rect 17598 4299 17599 4325
rect 17599 4299 17625 4325
rect 17625 4299 17626 4325
rect 17598 4298 17626 4299
rect 17650 4325 17678 4326
rect 17650 4299 17651 4325
rect 17651 4299 17677 4325
rect 17677 4299 17678 4325
rect 17650 4298 17678 4299
rect 17702 4325 17730 4326
rect 17702 4299 17703 4325
rect 17703 4299 17729 4325
rect 17729 4299 17730 4325
rect 17702 4298 17730 4299
rect 17598 3541 17626 3542
rect 17598 3515 17599 3541
rect 17599 3515 17625 3541
rect 17625 3515 17626 3541
rect 17598 3514 17626 3515
rect 17650 3541 17678 3542
rect 17650 3515 17651 3541
rect 17651 3515 17677 3541
rect 17677 3515 17678 3541
rect 17650 3514 17678 3515
rect 17702 3541 17730 3542
rect 17702 3515 17703 3541
rect 17703 3515 17729 3541
rect 17729 3515 17730 3541
rect 17702 3514 17730 3515
rect 17598 2757 17626 2758
rect 17598 2731 17599 2757
rect 17599 2731 17625 2757
rect 17625 2731 17626 2757
rect 17598 2730 17626 2731
rect 17650 2757 17678 2758
rect 17650 2731 17651 2757
rect 17651 2731 17677 2757
rect 17677 2731 17678 2757
rect 17650 2730 17678 2731
rect 17702 2757 17730 2758
rect 17702 2731 17703 2757
rect 17703 2731 17729 2757
rect 17729 2731 17730 2757
rect 17702 2730 17730 2731
rect 17598 1973 17626 1974
rect 17598 1947 17599 1973
rect 17599 1947 17625 1973
rect 17625 1947 17626 1973
rect 17598 1946 17626 1947
rect 17650 1973 17678 1974
rect 17650 1947 17651 1973
rect 17651 1947 17677 1973
rect 17677 1947 17678 1973
rect 17650 1946 17678 1947
rect 17702 1973 17730 1974
rect 17702 1947 17703 1973
rect 17703 1947 17729 1973
rect 17729 1947 17730 1973
rect 17702 1946 17730 1947
rect 14686 1833 14714 1834
rect 14686 1807 14687 1833
rect 14687 1807 14713 1833
rect 14713 1807 14714 1833
rect 14686 1806 14714 1807
<< metal3 >>
rect 2233 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2375 19222
rect 17593 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17735 19222
rect 10761 19110 10766 19138
rect 10794 19110 11214 19138
rect 11242 19110 11247 19138
rect 12105 19110 12110 19138
rect 12138 19110 12782 19138
rect 12810 19110 12815 19138
rect 10537 18942 10542 18970
rect 10570 18942 11102 18970
rect 11130 18942 11135 18970
rect 9913 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10055 18830
rect 8745 18718 8750 18746
rect 8778 18718 9366 18746
rect 9394 18718 9399 18746
rect 10425 18718 10430 18746
rect 10458 18718 11046 18746
rect 11074 18718 11079 18746
rect 2233 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2375 18438
rect 17593 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17735 18438
rect 9913 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10055 18046
rect 2233 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2375 17654
rect 17593 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17735 17654
rect 9913 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10055 17262
rect 20600 17178 21000 17192
rect 20113 17150 20118 17178
rect 20146 17150 21000 17178
rect 20600 17136 21000 17150
rect 2233 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2375 16870
rect 17593 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17735 16870
rect 9913 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10055 16478
rect 2233 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2375 16086
rect 17593 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17735 16086
rect 9913 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10055 15694
rect 2233 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2375 15302
rect 17593 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17735 15302
rect 9913 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10055 14910
rect 2233 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2375 14518
rect 17593 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17735 14518
rect 9913 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10055 14126
rect 10313 14014 10318 14042
rect 10346 14014 10822 14042
rect 10850 14014 11158 14042
rect 11186 14014 11191 14042
rect 10705 13958 10710 13986
rect 10738 13958 10990 13986
rect 11018 13958 11023 13986
rect 9417 13902 9422 13930
rect 9450 13902 10094 13930
rect 10066 13874 10094 13902
rect 10066 13846 10374 13874
rect 10402 13846 11438 13874
rect 11466 13846 11942 13874
rect 11970 13846 11975 13874
rect 0 13818 400 13832
rect 0 13790 2086 13818
rect 2114 13790 2119 13818
rect 0 13776 400 13790
rect 2233 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2375 13734
rect 17593 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17735 13734
rect 9809 13566 9814 13594
rect 9842 13566 10710 13594
rect 10738 13566 10743 13594
rect 13449 13510 13454 13538
rect 13482 13510 14238 13538
rect 14266 13510 18830 13538
rect 18858 13510 18863 13538
rect 20600 13482 21000 13496
rect 9473 13454 9478 13482
rect 9506 13454 10598 13482
rect 10626 13454 10631 13482
rect 12217 13454 12222 13482
rect 12250 13454 13398 13482
rect 13426 13454 13431 13482
rect 19950 13454 21000 13482
rect 19950 13426 19978 13454
rect 20600 13440 21000 13454
rect 19945 13398 19950 13426
rect 19978 13398 19983 13426
rect 8745 13342 8750 13370
rect 8778 13342 9534 13370
rect 9562 13342 9567 13370
rect 9913 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10055 13342
rect 10313 13174 10318 13202
rect 10346 13174 10766 13202
rect 10794 13174 12278 13202
rect 12306 13174 12311 13202
rect 14401 13174 14406 13202
rect 14434 13174 15974 13202
rect 15946 13146 15974 13174
rect 20600 13146 21000 13160
rect 2137 13118 2142 13146
rect 2170 13118 5950 13146
rect 5978 13118 5983 13146
rect 10145 13118 10150 13146
rect 10178 13118 11214 13146
rect 11242 13118 11247 13146
rect 15946 13118 18830 13146
rect 18858 13118 18863 13146
rect 20001 13118 20006 13146
rect 20034 13118 21000 13146
rect 20600 13104 21000 13118
rect 7345 13062 7350 13090
rect 7378 13062 8134 13090
rect 8162 13062 8167 13090
rect 11937 13062 11942 13090
rect 11970 13062 12334 13090
rect 12362 13062 12367 13090
rect 2233 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2375 12950
rect 17593 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17735 12950
rect 0 12810 400 12824
rect 0 12782 966 12810
rect 994 12782 999 12810
rect 12497 12782 12502 12810
rect 12530 12782 13006 12810
rect 13034 12782 13039 12810
rect 0 12768 400 12782
rect 2137 12726 2142 12754
rect 2170 12726 5446 12754
rect 5474 12726 5479 12754
rect 11489 12726 11494 12754
rect 11522 12726 12110 12754
rect 12138 12726 12143 12754
rect 13673 12726 13678 12754
rect 13706 12726 14126 12754
rect 14154 12726 18830 12754
rect 18858 12726 18863 12754
rect 10873 12670 10878 12698
rect 10906 12670 11326 12698
rect 11354 12670 11359 12698
rect 9809 12614 9814 12642
rect 9842 12614 10318 12642
rect 10346 12614 10351 12642
rect 10761 12614 10766 12642
rect 10794 12614 12110 12642
rect 12138 12614 12726 12642
rect 12754 12614 12759 12642
rect 7625 12558 7630 12586
rect 7658 12558 8470 12586
rect 8498 12558 9086 12586
rect 9114 12558 9119 12586
rect 9913 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10055 12558
rect 8297 12502 8302 12530
rect 8330 12502 9422 12530
rect 9450 12502 9455 12530
rect 0 12474 400 12488
rect 20600 12474 21000 12488
rect 0 12446 1022 12474
rect 1050 12446 1055 12474
rect 12441 12446 12446 12474
rect 12474 12446 12950 12474
rect 12978 12446 12983 12474
rect 20001 12446 20006 12474
rect 20034 12446 21000 12474
rect 0 12432 400 12446
rect 20600 12432 21000 12446
rect 5945 12390 5950 12418
rect 5978 12390 7798 12418
rect 7826 12390 7831 12418
rect 8969 12390 8974 12418
rect 9002 12390 9366 12418
rect 9394 12390 9399 12418
rect 9753 12390 9758 12418
rect 9786 12390 10598 12418
rect 10626 12390 10631 12418
rect 12833 12390 12838 12418
rect 12866 12390 13622 12418
rect 13650 12390 13655 12418
rect 8241 12334 8246 12362
rect 8274 12334 8918 12362
rect 8946 12334 8951 12362
rect 9137 12334 9142 12362
rect 9170 12334 10150 12362
rect 10178 12334 10183 12362
rect 6897 12278 6902 12306
rect 6930 12278 7126 12306
rect 7154 12278 7406 12306
rect 7434 12278 7630 12306
rect 7658 12278 7663 12306
rect 9753 12278 9758 12306
rect 9786 12278 10654 12306
rect 10682 12278 12838 12306
rect 12866 12278 12871 12306
rect 10089 12166 10094 12194
rect 10122 12166 11718 12194
rect 11746 12166 11751 12194
rect 2233 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2375 12166
rect 17593 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17735 12166
rect 6953 12054 6958 12082
rect 6986 12054 7182 12082
rect 7210 12054 10094 12082
rect 10122 12054 10127 12082
rect 5441 11998 5446 12026
rect 5474 11998 6734 12026
rect 6762 11998 6767 12026
rect 11657 11942 11662 11970
rect 11690 11942 12894 11970
rect 12922 11942 12927 11970
rect 7065 11886 7070 11914
rect 7098 11886 8246 11914
rect 8274 11886 8279 11914
rect 9081 11886 9086 11914
rect 9114 11886 10430 11914
rect 10458 11886 10463 11914
rect 6505 11830 6510 11858
rect 6538 11830 7182 11858
rect 7210 11830 7215 11858
rect 8801 11830 8806 11858
rect 8834 11830 9982 11858
rect 10010 11830 10015 11858
rect 10873 11830 10878 11858
rect 10906 11830 11270 11858
rect 11298 11830 11303 11858
rect 7289 11774 7294 11802
rect 7322 11774 7574 11802
rect 7602 11774 8694 11802
rect 8722 11774 8727 11802
rect 9913 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10055 11774
rect 10094 11718 10934 11746
rect 10962 11718 10967 11746
rect 10094 11690 10122 11718
rect 9585 11662 9590 11690
rect 9618 11662 10122 11690
rect 10425 11606 10430 11634
rect 10458 11606 10934 11634
rect 10962 11606 11942 11634
rect 11970 11606 12558 11634
rect 12586 11606 12591 11634
rect 7513 11550 7518 11578
rect 7546 11550 7574 11578
rect 7602 11550 7854 11578
rect 7882 11550 7887 11578
rect 8409 11550 8414 11578
rect 8442 11550 8862 11578
rect 8890 11550 8895 11578
rect 9753 11494 9758 11522
rect 9786 11494 9805 11522
rect 20600 11466 21000 11480
rect 20001 11438 20006 11466
rect 20034 11438 21000 11466
rect 20600 11424 21000 11438
rect 2233 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2375 11382
rect 17593 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17735 11382
rect 5385 11326 5390 11354
rect 5418 11326 6958 11354
rect 6986 11326 7462 11354
rect 7490 11326 7495 11354
rect 11489 11326 11494 11354
rect 11522 11326 11998 11354
rect 12026 11326 12031 11354
rect 12329 11270 12334 11298
rect 12362 11270 18830 11298
rect 18858 11270 18863 11298
rect 6449 11214 6454 11242
rect 6482 11214 7070 11242
rect 7098 11214 7294 11242
rect 7322 11214 7327 11242
rect 9459 11158 9478 11186
rect 9506 11158 9511 11186
rect 10635 11158 10654 11186
rect 10682 11158 10687 11186
rect 12553 11158 12558 11186
rect 12586 11158 12894 11186
rect 12922 11158 12927 11186
rect 13617 11158 13622 11186
rect 13650 11158 14294 11186
rect 14322 11158 18830 11186
rect 18858 11158 18863 11186
rect 20600 11130 21000 11144
rect 7345 11102 7350 11130
rect 7378 11102 7910 11130
rect 7938 11102 7943 11130
rect 8913 11102 8918 11130
rect 8946 11102 10262 11130
rect 10290 11102 10878 11130
rect 10906 11102 10911 11130
rect 20001 11102 20006 11130
rect 20034 11102 21000 11130
rect 20600 11088 21000 11102
rect 7457 11046 7462 11074
rect 7490 11046 8022 11074
rect 8050 11046 8526 11074
rect 8554 11046 9086 11074
rect 9114 11046 9119 11074
rect 9235 11046 9254 11074
rect 9282 11046 9287 11074
rect 9473 11046 9478 11074
rect 9506 11046 10038 11074
rect 10066 11046 10071 11074
rect 10145 11046 10150 11074
rect 10178 11046 10710 11074
rect 10738 11046 11606 11074
rect 11634 11046 11639 11074
rect 7905 10990 7910 11018
rect 7938 10990 9646 11018
rect 9674 10990 9679 11018
rect 9739 10990 9758 11018
rect 9786 10990 9791 11018
rect 10579 10990 10598 11018
rect 10626 10990 10631 11018
rect 9913 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10055 10990
rect 5049 10934 5054 10962
rect 5082 10934 6790 10962
rect 6818 10934 6823 10962
rect 7513 10878 7518 10906
rect 7546 10878 7742 10906
rect 7770 10878 7775 10906
rect 9697 10878 9702 10906
rect 9730 10878 10150 10906
rect 10178 10878 10183 10906
rect 10705 10878 10710 10906
rect 10738 10878 10743 10906
rect 11713 10878 11718 10906
rect 11746 10878 13510 10906
rect 13538 10878 13543 10906
rect 10710 10850 10738 10878
rect 10710 10822 10878 10850
rect 10906 10822 10911 10850
rect 11601 10822 11606 10850
rect 11634 10822 12110 10850
rect 12138 10822 12143 10850
rect 9641 10766 9646 10794
rect 9674 10766 9758 10794
rect 9786 10766 10934 10794
rect 10962 10766 10967 10794
rect 11937 10766 11942 10794
rect 11970 10766 13678 10794
rect 13706 10766 13711 10794
rect 7625 10710 7630 10738
rect 7658 10710 8302 10738
rect 8330 10710 8335 10738
rect 8465 10710 8470 10738
rect 8498 10710 9030 10738
rect 9058 10710 9063 10738
rect 10369 10710 10374 10738
rect 10402 10710 11494 10738
rect 11522 10710 11718 10738
rect 11746 10710 11751 10738
rect 8801 10654 8806 10682
rect 8834 10654 9422 10682
rect 9450 10654 9814 10682
rect 9842 10654 12054 10682
rect 12082 10654 12087 10682
rect 5385 10598 5390 10626
rect 5418 10598 6566 10626
rect 6594 10598 7574 10626
rect 7602 10598 11214 10626
rect 11242 10598 11247 10626
rect 2233 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2375 10598
rect 17593 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17735 10598
rect 7233 10542 7238 10570
rect 7266 10542 8134 10570
rect 8162 10542 9030 10570
rect 9058 10542 9063 10570
rect 10593 10542 10598 10570
rect 10626 10542 10710 10570
rect 10738 10542 10743 10570
rect 7681 10486 7686 10514
rect 7714 10486 8246 10514
rect 8274 10486 8582 10514
rect 8610 10486 11270 10514
rect 11298 10486 11303 10514
rect 20600 10458 21000 10472
rect 6449 10430 6454 10458
rect 6482 10430 6846 10458
rect 6874 10430 7126 10458
rect 7154 10430 7159 10458
rect 9137 10430 9142 10458
rect 9170 10430 11158 10458
rect 11186 10430 11382 10458
rect 11410 10430 11415 10458
rect 19945 10430 19950 10458
rect 19978 10430 21000 10458
rect 20600 10416 21000 10430
rect 6897 10374 6902 10402
rect 6930 10374 7518 10402
rect 7546 10374 7551 10402
rect 8745 10374 8750 10402
rect 8778 10374 10094 10402
rect 10122 10374 10127 10402
rect 10201 10374 10206 10402
rect 10234 10374 11046 10402
rect 11074 10374 11494 10402
rect 11522 10374 11527 10402
rect 18825 10374 18830 10402
rect 18858 10374 18863 10402
rect 7401 10318 7406 10346
rect 7434 10318 7966 10346
rect 7994 10318 7999 10346
rect 9137 10318 9142 10346
rect 9170 10318 9982 10346
rect 10010 10318 10015 10346
rect 11209 10318 11214 10346
rect 11242 10318 11886 10346
rect 11914 10318 12110 10346
rect 12138 10318 12143 10346
rect 13785 10318 13790 10346
rect 13818 10318 14294 10346
rect 14322 10318 14630 10346
rect 14658 10318 18718 10346
rect 18746 10318 18751 10346
rect 18830 10290 18858 10374
rect 2081 10262 2086 10290
rect 2114 10262 8862 10290
rect 8890 10262 8895 10290
rect 9641 10262 9646 10290
rect 9674 10262 9758 10290
rect 9786 10262 9791 10290
rect 10369 10262 10374 10290
rect 10402 10262 10766 10290
rect 10794 10262 10799 10290
rect 14737 10262 14742 10290
rect 14770 10262 18858 10290
rect 9913 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10055 10206
rect 20600 10122 21000 10136
rect 7849 10094 7854 10122
rect 7882 10094 11382 10122
rect 11410 10094 11415 10122
rect 20001 10094 20006 10122
rect 20034 10094 21000 10122
rect 20600 10080 21000 10094
rect 9529 10038 9534 10066
rect 9562 10038 10150 10066
rect 10178 10038 10183 10066
rect 11321 10038 11326 10066
rect 11354 10038 11942 10066
rect 11970 10038 11975 10066
rect 7737 9982 7742 10010
rect 7770 9982 8078 10010
rect 8106 9982 8806 10010
rect 8834 9982 8839 10010
rect 10089 9982 10094 10010
rect 10122 9982 12894 10010
rect 12922 9982 12927 10010
rect 13225 9982 13230 10010
rect 13258 9982 13454 10010
rect 13426 9954 13454 9982
rect 7961 9926 7966 9954
rect 7994 9926 10206 9954
rect 10234 9926 10239 9954
rect 11937 9926 11942 9954
rect 11970 9926 12782 9954
rect 12810 9926 13006 9954
rect 13034 9926 13039 9954
rect 13426 9926 13622 9954
rect 13650 9926 13655 9954
rect 11746 9870 13062 9898
rect 13090 9870 13342 9898
rect 13370 9870 13375 9898
rect 11746 9842 11774 9870
rect 10201 9814 10206 9842
rect 10234 9814 11774 9842
rect 2233 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2375 9814
rect 17593 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17735 9814
rect 8185 9758 8190 9786
rect 8218 9758 8414 9786
rect 8442 9758 10094 9786
rect 10122 9758 10127 9786
rect 8297 9702 8302 9730
rect 8330 9702 10710 9730
rect 10738 9702 10743 9730
rect 9249 9646 9254 9674
rect 9282 9646 10206 9674
rect 10234 9646 10239 9674
rect 10369 9646 10374 9674
rect 10402 9646 10654 9674
rect 10682 9646 10687 9674
rect 8521 9590 8526 9618
rect 8554 9590 8974 9618
rect 9002 9590 9007 9618
rect 9305 9590 9310 9618
rect 9338 9590 9478 9618
rect 9506 9590 10598 9618
rect 10626 9590 10631 9618
rect 11769 9590 11774 9618
rect 11802 9590 12110 9618
rect 12138 9590 12894 9618
rect 12922 9590 12927 9618
rect 13673 9590 13678 9618
rect 13706 9590 14294 9618
rect 14322 9590 18830 9618
rect 18858 9590 18863 9618
rect 7737 9534 7742 9562
rect 7770 9534 8134 9562
rect 8162 9534 8167 9562
rect 8297 9534 8302 9562
rect 8330 9534 8862 9562
rect 8890 9534 10374 9562
rect 10402 9534 10407 9562
rect 10635 9534 10654 9562
rect 10682 9534 10687 9562
rect 10929 9534 10934 9562
rect 10962 9534 11662 9562
rect 11690 9534 12390 9562
rect 12418 9534 12423 9562
rect 13113 9534 13118 9562
rect 13146 9534 13566 9562
rect 13594 9534 13599 9562
rect 7625 9478 7630 9506
rect 7658 9478 8414 9506
rect 8442 9478 8447 9506
rect 8801 9478 8806 9506
rect 8834 9478 9086 9506
rect 9114 9478 9119 9506
rect 9417 9478 9422 9506
rect 9450 9478 10318 9506
rect 10346 9478 10351 9506
rect 11377 9478 11382 9506
rect 11410 9478 11998 9506
rect 12026 9478 12031 9506
rect 12553 9478 12558 9506
rect 12586 9478 13734 9506
rect 13762 9478 13767 9506
rect 9086 9450 9114 9478
rect 20600 9450 21000 9464
rect 9086 9422 9590 9450
rect 9618 9422 9623 9450
rect 20001 9422 20006 9450
rect 20034 9422 21000 9450
rect 9590 9338 9618 9422
rect 9913 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10055 9422
rect 20600 9408 21000 9422
rect 10537 9366 10542 9394
rect 10570 9366 11326 9394
rect 11354 9366 11359 9394
rect 9590 9310 9870 9338
rect 9898 9310 9903 9338
rect 9982 9310 11158 9338
rect 11186 9310 11191 9338
rect 9982 9282 10010 9310
rect 8409 9254 8414 9282
rect 8442 9254 8694 9282
rect 8722 9254 9254 9282
rect 9282 9254 9534 9282
rect 9562 9254 10010 9282
rect 6225 9198 6230 9226
rect 6258 9198 11438 9226
rect 11466 9198 11471 9226
rect 6057 9142 6062 9170
rect 6090 9142 7014 9170
rect 7042 9142 7574 9170
rect 7602 9142 7607 9170
rect 8633 9142 8638 9170
rect 8666 9142 9198 9170
rect 9226 9142 10094 9170
rect 10122 9142 10127 9170
rect 8577 9086 8582 9114
rect 8610 9086 8862 9114
rect 8890 9086 8895 9114
rect 9137 9086 9142 9114
rect 9170 9086 11046 9114
rect 11074 9086 11550 9114
rect 11578 9086 11583 9114
rect 7961 9030 7966 9058
rect 7994 9030 9366 9058
rect 9394 9030 9534 9058
rect 9562 9030 10822 9058
rect 10850 9030 10855 9058
rect 2233 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2375 9030
rect 17593 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17735 9030
rect 9137 8862 9142 8890
rect 9170 8862 9646 8890
rect 9674 8862 9679 8890
rect 13617 8806 13622 8834
rect 13650 8806 14294 8834
rect 14322 8806 18830 8834
rect 18858 8806 18863 8834
rect 20600 8778 21000 8792
rect 6449 8750 6454 8778
rect 6482 8750 7742 8778
rect 7770 8750 7775 8778
rect 8857 8750 8862 8778
rect 8890 8750 9870 8778
rect 9898 8750 10710 8778
rect 10738 8750 10743 8778
rect 20001 8750 20006 8778
rect 20034 8750 21000 8778
rect 20600 8736 21000 8750
rect 8409 8694 8414 8722
rect 8442 8694 8750 8722
rect 8778 8694 8783 8722
rect 9081 8694 9086 8722
rect 9114 8694 9198 8722
rect 9226 8694 9231 8722
rect 7513 8638 7518 8666
rect 7546 8638 8078 8666
rect 8106 8638 8582 8666
rect 8610 8638 8615 8666
rect 9913 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10055 8638
rect 8353 8526 8358 8554
rect 8386 8526 9030 8554
rect 9058 8526 9366 8554
rect 9394 8526 9399 8554
rect 10033 8526 10038 8554
rect 10066 8526 10430 8554
rect 10458 8526 10463 8554
rect 7513 8470 7518 8498
rect 7546 8470 7966 8498
rect 7994 8470 8302 8498
rect 8330 8470 8335 8498
rect 7737 8414 7742 8442
rect 7770 8414 10934 8442
rect 10962 8414 10967 8442
rect 13426 8414 13510 8442
rect 13538 8414 13543 8442
rect 8918 8386 8946 8414
rect 8913 8358 8918 8386
rect 8946 8358 8951 8386
rect 13426 8330 13454 8414
rect 12945 8302 12950 8330
rect 12978 8302 13454 8330
rect 2233 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2375 8246
rect 17593 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17735 8246
rect 8521 8134 8526 8162
rect 8554 8134 8862 8162
rect 8890 8134 9310 8162
rect 9338 8134 9343 8162
rect 10257 8078 10262 8106
rect 10290 8078 10766 8106
rect 10794 8078 10799 8106
rect 9417 8022 9422 8050
rect 9450 8022 10990 8050
rect 11018 8022 11023 8050
rect 12161 8022 12166 8050
rect 12194 8022 13062 8050
rect 13090 8022 13095 8050
rect 10145 7966 10150 7994
rect 10178 7966 10654 7994
rect 10682 7966 10687 7994
rect 11825 7966 11830 7994
rect 11858 7966 12950 7994
rect 12978 7966 12983 7994
rect 9753 7910 9758 7938
rect 9786 7910 9982 7938
rect 10010 7910 10015 7938
rect 10873 7910 10878 7938
rect 10906 7910 11886 7938
rect 11914 7910 11919 7938
rect 9913 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10055 7854
rect 20600 7770 21000 7784
rect 20001 7742 20006 7770
rect 20034 7742 21000 7770
rect 20600 7728 21000 7742
rect 8974 7686 9702 7714
rect 9730 7686 9735 7714
rect 8974 7658 9002 7686
rect 8969 7630 8974 7658
rect 9002 7630 9007 7658
rect 9249 7630 9254 7658
rect 9282 7630 9814 7658
rect 9842 7630 9847 7658
rect 7345 7574 7350 7602
rect 7378 7574 8918 7602
rect 8946 7574 8951 7602
rect 9137 7574 9142 7602
rect 9170 7574 10150 7602
rect 10178 7574 10183 7602
rect 13561 7574 13566 7602
rect 13594 7574 14238 7602
rect 14266 7574 18830 7602
rect 18858 7574 18863 7602
rect 10929 7518 10934 7546
rect 10962 7518 11830 7546
rect 11858 7518 12334 7546
rect 12362 7518 12367 7546
rect 2233 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2375 7462
rect 17593 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17735 7462
rect 10761 7294 10766 7322
rect 10794 7294 11158 7322
rect 11186 7294 11191 7322
rect 9529 7238 9534 7266
rect 9562 7238 10262 7266
rect 10290 7238 10295 7266
rect 10369 7238 10374 7266
rect 10402 7238 11270 7266
rect 11298 7238 11303 7266
rect 12889 7126 12894 7154
rect 12922 7126 13454 7154
rect 13482 7126 13487 7154
rect 9913 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10055 7070
rect 8297 6902 8302 6930
rect 8330 6902 9142 6930
rect 9170 6902 9175 6930
rect 9305 6902 9310 6930
rect 9338 6902 10206 6930
rect 10234 6902 10239 6930
rect 8409 6846 8414 6874
rect 8442 6846 9646 6874
rect 9674 6846 9679 6874
rect 9753 6846 9758 6874
rect 9786 6846 10038 6874
rect 10066 6846 10071 6874
rect 11209 6846 11214 6874
rect 11242 6846 12614 6874
rect 12642 6846 12647 6874
rect 9025 6790 9030 6818
rect 9058 6790 9870 6818
rect 9898 6790 9903 6818
rect 8689 6734 8694 6762
rect 8722 6734 10318 6762
rect 10346 6734 10351 6762
rect 12217 6734 12222 6762
rect 12250 6734 12670 6762
rect 12698 6734 12703 6762
rect 2233 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2375 6678
rect 17593 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17735 6678
rect 13449 6510 13454 6538
rect 13482 6510 14294 6538
rect 14322 6510 14327 6538
rect 9913 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10055 6286
rect 11377 5894 11382 5922
rect 11410 5894 11662 5922
rect 11690 5894 12278 5922
rect 12306 5894 12311 5922
rect 2233 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2375 5894
rect 17593 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17735 5894
rect 9913 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10055 5502
rect 2233 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2375 5110
rect 17593 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17735 5110
rect 9913 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10055 4718
rect 2233 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2375 4326
rect 17593 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17735 4326
rect 9913 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10055 3934
rect 2233 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2375 3542
rect 17593 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17735 3542
rect 9913 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10055 3150
rect 2233 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2375 2758
rect 17593 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17735 2758
rect 9913 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10055 2366
rect 8745 2030 8750 2058
rect 8778 2030 9366 2058
rect 9394 2030 9399 2058
rect 12105 2030 12110 2058
rect 12138 2030 13118 2058
rect 13146 2030 13151 2058
rect 2233 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2375 1974
rect 17593 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17735 1974
rect 11433 1806 11438 1834
rect 11466 1806 12782 1834
rect 12810 1806 12815 1834
rect 13169 1806 13174 1834
rect 13202 1806 14686 1834
rect 14714 1806 14719 1834
rect 10089 1694 10094 1722
rect 10122 1694 10878 1722
rect 10906 1694 10911 1722
rect 9913 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10055 1582
<< via3 >>
rect 2238 19194 2266 19222
rect 2290 19194 2318 19222
rect 2342 19194 2370 19222
rect 17598 19194 17626 19222
rect 17650 19194 17678 19222
rect 17702 19194 17730 19222
rect 9918 18802 9946 18830
rect 9970 18802 9998 18830
rect 10022 18802 10050 18830
rect 2238 18410 2266 18438
rect 2290 18410 2318 18438
rect 2342 18410 2370 18438
rect 17598 18410 17626 18438
rect 17650 18410 17678 18438
rect 17702 18410 17730 18438
rect 9918 18018 9946 18046
rect 9970 18018 9998 18046
rect 10022 18018 10050 18046
rect 2238 17626 2266 17654
rect 2290 17626 2318 17654
rect 2342 17626 2370 17654
rect 17598 17626 17626 17654
rect 17650 17626 17678 17654
rect 17702 17626 17730 17654
rect 9918 17234 9946 17262
rect 9970 17234 9998 17262
rect 10022 17234 10050 17262
rect 2238 16842 2266 16870
rect 2290 16842 2318 16870
rect 2342 16842 2370 16870
rect 17598 16842 17626 16870
rect 17650 16842 17678 16870
rect 17702 16842 17730 16870
rect 9918 16450 9946 16478
rect 9970 16450 9998 16478
rect 10022 16450 10050 16478
rect 2238 16058 2266 16086
rect 2290 16058 2318 16086
rect 2342 16058 2370 16086
rect 17598 16058 17626 16086
rect 17650 16058 17678 16086
rect 17702 16058 17730 16086
rect 9918 15666 9946 15694
rect 9970 15666 9998 15694
rect 10022 15666 10050 15694
rect 2238 15274 2266 15302
rect 2290 15274 2318 15302
rect 2342 15274 2370 15302
rect 17598 15274 17626 15302
rect 17650 15274 17678 15302
rect 17702 15274 17730 15302
rect 9918 14882 9946 14910
rect 9970 14882 9998 14910
rect 10022 14882 10050 14910
rect 2238 14490 2266 14518
rect 2290 14490 2318 14518
rect 2342 14490 2370 14518
rect 17598 14490 17626 14518
rect 17650 14490 17678 14518
rect 17702 14490 17730 14518
rect 9918 14098 9946 14126
rect 9970 14098 9998 14126
rect 10022 14098 10050 14126
rect 2238 13706 2266 13734
rect 2290 13706 2318 13734
rect 2342 13706 2370 13734
rect 17598 13706 17626 13734
rect 17650 13706 17678 13734
rect 17702 13706 17730 13734
rect 9918 13314 9946 13342
rect 9970 13314 9998 13342
rect 10022 13314 10050 13342
rect 2238 12922 2266 12950
rect 2290 12922 2318 12950
rect 2342 12922 2370 12950
rect 17598 12922 17626 12950
rect 17650 12922 17678 12950
rect 17702 12922 17730 12950
rect 9918 12530 9946 12558
rect 9970 12530 9998 12558
rect 10022 12530 10050 12558
rect 2238 12138 2266 12166
rect 2290 12138 2318 12166
rect 2342 12138 2370 12166
rect 17598 12138 17626 12166
rect 17650 12138 17678 12166
rect 17702 12138 17730 12166
rect 9918 11746 9946 11774
rect 9970 11746 9998 11774
rect 10022 11746 10050 11774
rect 9758 11494 9786 11522
rect 2238 11354 2266 11382
rect 2290 11354 2318 11382
rect 2342 11354 2370 11382
rect 17598 11354 17626 11382
rect 17650 11354 17678 11382
rect 17702 11354 17730 11382
rect 9478 11158 9506 11186
rect 10654 11158 10682 11186
rect 9254 11046 9282 11074
rect 9758 10990 9786 11018
rect 10598 10990 10626 11018
rect 9918 10962 9946 10990
rect 9970 10962 9998 10990
rect 10022 10962 10050 10990
rect 9758 10766 9786 10794
rect 2238 10570 2266 10598
rect 2290 10570 2318 10598
rect 2342 10570 2370 10598
rect 17598 10570 17626 10598
rect 17650 10570 17678 10598
rect 17702 10570 17730 10598
rect 10598 10542 10626 10570
rect 9758 10262 9786 10290
rect 9918 10178 9946 10206
rect 9970 10178 9998 10206
rect 10022 10178 10050 10206
rect 2238 9786 2266 9814
rect 2290 9786 2318 9814
rect 2342 9786 2370 9814
rect 17598 9786 17626 9814
rect 17650 9786 17678 9814
rect 17702 9786 17730 9814
rect 9254 9646 9282 9674
rect 9478 9590 9506 9618
rect 10654 9534 10682 9562
rect 9918 9394 9946 9422
rect 9970 9394 9998 9422
rect 10022 9394 10050 9422
rect 2238 9002 2266 9030
rect 2290 9002 2318 9030
rect 2342 9002 2370 9030
rect 17598 9002 17626 9030
rect 17650 9002 17678 9030
rect 17702 9002 17730 9030
rect 9918 8610 9946 8638
rect 9970 8610 9998 8638
rect 10022 8610 10050 8638
rect 2238 8218 2266 8246
rect 2290 8218 2318 8246
rect 2342 8218 2370 8246
rect 17598 8218 17626 8246
rect 17650 8218 17678 8246
rect 17702 8218 17730 8246
rect 10654 7966 10682 7994
rect 9918 7826 9946 7854
rect 9970 7826 9998 7854
rect 10022 7826 10050 7854
rect 2238 7434 2266 7462
rect 2290 7434 2318 7462
rect 2342 7434 2370 7462
rect 17598 7434 17626 7462
rect 17650 7434 17678 7462
rect 17702 7434 17730 7462
rect 9918 7042 9946 7070
rect 9970 7042 9998 7070
rect 10022 7042 10050 7070
rect 2238 6650 2266 6678
rect 2290 6650 2318 6678
rect 2342 6650 2370 6678
rect 17598 6650 17626 6678
rect 17650 6650 17678 6678
rect 17702 6650 17730 6678
rect 9918 6258 9946 6286
rect 9970 6258 9998 6286
rect 10022 6258 10050 6286
rect 2238 5866 2266 5894
rect 2290 5866 2318 5894
rect 2342 5866 2370 5894
rect 17598 5866 17626 5894
rect 17650 5866 17678 5894
rect 17702 5866 17730 5894
rect 9918 5474 9946 5502
rect 9970 5474 9998 5502
rect 10022 5474 10050 5502
rect 2238 5082 2266 5110
rect 2290 5082 2318 5110
rect 2342 5082 2370 5110
rect 17598 5082 17626 5110
rect 17650 5082 17678 5110
rect 17702 5082 17730 5110
rect 9918 4690 9946 4718
rect 9970 4690 9998 4718
rect 10022 4690 10050 4718
rect 2238 4298 2266 4326
rect 2290 4298 2318 4326
rect 2342 4298 2370 4326
rect 17598 4298 17626 4326
rect 17650 4298 17678 4326
rect 17702 4298 17730 4326
rect 9918 3906 9946 3934
rect 9970 3906 9998 3934
rect 10022 3906 10050 3934
rect 2238 3514 2266 3542
rect 2290 3514 2318 3542
rect 2342 3514 2370 3542
rect 17598 3514 17626 3542
rect 17650 3514 17678 3542
rect 17702 3514 17730 3542
rect 9918 3122 9946 3150
rect 9970 3122 9998 3150
rect 10022 3122 10050 3150
rect 2238 2730 2266 2758
rect 2290 2730 2318 2758
rect 2342 2730 2370 2758
rect 17598 2730 17626 2758
rect 17650 2730 17678 2758
rect 17702 2730 17730 2758
rect 9918 2338 9946 2366
rect 9970 2338 9998 2366
rect 10022 2338 10050 2366
rect 2238 1946 2266 1974
rect 2290 1946 2318 1974
rect 2342 1946 2370 1974
rect 17598 1946 17626 1974
rect 17650 1946 17678 1974
rect 17702 1946 17730 1974
rect 9918 1554 9946 1582
rect 9970 1554 9998 1582
rect 10022 1554 10050 1582
<< metal4 >>
rect 2224 19222 2384 19238
rect 2224 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2384 19222
rect 2224 18438 2384 19194
rect 2224 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2384 18438
rect 2224 17654 2384 18410
rect 2224 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2384 17654
rect 2224 16870 2384 17626
rect 2224 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2384 16870
rect 2224 16086 2384 16842
rect 2224 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2384 16086
rect 2224 15302 2384 16058
rect 2224 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2384 15302
rect 2224 14518 2384 15274
rect 2224 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2384 14518
rect 2224 13734 2384 14490
rect 2224 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2384 13734
rect 2224 12950 2384 13706
rect 2224 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2384 12950
rect 2224 12166 2384 12922
rect 2224 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2384 12166
rect 2224 11382 2384 12138
rect 9904 18830 10064 19238
rect 9904 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10064 18830
rect 9904 18046 10064 18802
rect 9904 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10064 18046
rect 9904 17262 10064 18018
rect 9904 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10064 17262
rect 9904 16478 10064 17234
rect 9904 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10064 16478
rect 9904 15694 10064 16450
rect 9904 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10064 15694
rect 9904 14910 10064 15666
rect 9904 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10064 14910
rect 9904 14126 10064 14882
rect 9904 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10064 14126
rect 9904 13342 10064 14098
rect 9904 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10064 13342
rect 9904 12558 10064 13314
rect 9904 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10064 12558
rect 9904 11774 10064 12530
rect 9904 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10064 11774
rect 2224 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2384 11382
rect 2224 10598 2384 11354
rect 9758 11522 9786 11527
rect 9478 11186 9506 11191
rect 2224 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2384 10598
rect 2224 9814 2384 10570
rect 2224 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2384 9814
rect 2224 9030 2384 9786
rect 9254 11074 9282 11079
rect 9254 9674 9282 11046
rect 9254 9641 9282 9646
rect 9478 9618 9506 11158
rect 9758 11018 9786 11494
rect 9758 10985 9786 10990
rect 9904 10990 10064 11746
rect 17584 19222 17744 19238
rect 17584 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17744 19222
rect 17584 18438 17744 19194
rect 17584 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17744 18438
rect 17584 17654 17744 18410
rect 17584 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17744 17654
rect 17584 16870 17744 17626
rect 17584 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17744 16870
rect 17584 16086 17744 16842
rect 17584 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17744 16086
rect 17584 15302 17744 16058
rect 17584 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17744 15302
rect 17584 14518 17744 15274
rect 17584 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17744 14518
rect 17584 13734 17744 14490
rect 17584 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17744 13734
rect 17584 12950 17744 13706
rect 17584 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17744 12950
rect 17584 12166 17744 12922
rect 17584 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17744 12166
rect 17584 11382 17744 12138
rect 17584 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17744 11382
rect 10654 11186 10682 11191
rect 9904 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10064 10990
rect 9758 10794 9786 10799
rect 9758 10290 9786 10766
rect 9758 10257 9786 10262
rect 9478 9585 9506 9590
rect 9904 10206 10064 10962
rect 10598 11018 10626 11023
rect 10598 10570 10626 10990
rect 10598 10537 10626 10542
rect 9904 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10064 10206
rect 2224 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2384 9030
rect 2224 8246 2384 9002
rect 2224 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2384 8246
rect 2224 7462 2384 8218
rect 2224 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2384 7462
rect 2224 6678 2384 7434
rect 2224 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2384 6678
rect 2224 5894 2384 6650
rect 2224 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2384 5894
rect 2224 5110 2384 5866
rect 2224 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2384 5110
rect 2224 4326 2384 5082
rect 2224 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2384 4326
rect 2224 3542 2384 4298
rect 2224 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2384 3542
rect 2224 2758 2384 3514
rect 2224 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2384 2758
rect 2224 1974 2384 2730
rect 2224 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2384 1974
rect 2224 1538 2384 1946
rect 9904 9422 10064 10178
rect 9904 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10064 9422
rect 9904 8638 10064 9394
rect 9904 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10064 8638
rect 9904 7854 10064 8610
rect 10654 9562 10682 11158
rect 10654 7994 10682 9534
rect 10654 7961 10682 7966
rect 17584 10598 17744 11354
rect 17584 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17744 10598
rect 17584 9814 17744 10570
rect 17584 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17744 9814
rect 17584 9030 17744 9786
rect 17584 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17744 9030
rect 17584 8246 17744 9002
rect 17584 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17744 8246
rect 9904 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10064 7854
rect 9904 7070 10064 7826
rect 9904 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10064 7070
rect 9904 6286 10064 7042
rect 9904 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10064 6286
rect 9904 5502 10064 6258
rect 9904 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10064 5502
rect 9904 4718 10064 5474
rect 9904 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10064 4718
rect 9904 3934 10064 4690
rect 9904 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10064 3934
rect 9904 3150 10064 3906
rect 9904 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10064 3150
rect 9904 2366 10064 3122
rect 9904 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10064 2366
rect 9904 1582 10064 2338
rect 9904 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10064 1582
rect 9904 1538 10064 1554
rect 17584 7462 17744 8218
rect 17584 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17744 7462
rect 17584 6678 17744 7434
rect 17584 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17744 6678
rect 17584 5894 17744 6650
rect 17584 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17744 5894
rect 17584 5110 17744 5866
rect 17584 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17744 5110
rect 17584 4326 17744 5082
rect 17584 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17744 4326
rect 17584 3542 17744 4298
rect 17584 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17744 3542
rect 17584 2758 17744 3514
rect 17584 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17744 2758
rect 17584 1974 17744 2730
rect 17584 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17744 1974
rect 17584 1538 17744 1946
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _112_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7392 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _113_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11312 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _114_
timestamp 1698175906
transform 1 0 12320 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _115_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 13832 0 1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _116_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 6776 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _117_
timestamp 1698175906
transform 1 0 7000 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _118_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7336 0 1 10192
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _119_
timestamp 1698175906
transform 1 0 8232 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _120_
timestamp 1698175906
transform 1 0 8960 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _121_
timestamp 1698175906
transform -1 0 11872 0 1 9408
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _122_
timestamp 1698175906
transform 1 0 11872 0 1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _123_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _124_
timestamp 1698175906
transform 1 0 8624 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _125_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8064 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _126_
timestamp 1698175906
transform 1 0 8624 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _127_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10584 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _128_
timestamp 1698175906
transform -1 0 10920 0 -1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _129_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12880 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _130_
timestamp 1698175906
transform 1 0 10136 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _131_
timestamp 1698175906
transform 1 0 7000 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _132_
timestamp 1698175906
transform 1 0 7224 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _133_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8904 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _134_
timestamp 1698175906
transform 1 0 11088 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _135_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13440 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _136_
timestamp 1698175906
transform 1 0 13216 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _137_
timestamp 1698175906
transform 1 0 11592 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _138_
timestamp 1698175906
transform 1 0 13440 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _139_
timestamp 1698175906
transform 1 0 12992 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _140_
timestamp 1698175906
transform 1 0 7728 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _141_
timestamp 1698175906
transform 1 0 10976 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _142_
timestamp 1698175906
transform -1 0 8456 0 -1 10976
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _143_
timestamp 1698175906
transform -1 0 7728 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _144_
timestamp 1698175906
transform -1 0 7224 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _145_
timestamp 1698175906
transform -1 0 8512 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _146_
timestamp 1698175906
transform 1 0 8456 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _147_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9688 0 1 10192
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _148_
timestamp 1698175906
transform 1 0 7616 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _149_
timestamp 1698175906
transform 1 0 11312 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _150_
timestamp 1698175906
transform 1 0 11312 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _151_
timestamp 1698175906
transform -1 0 9184 0 -1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _152_
timestamp 1698175906
transform 1 0 9968 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _153_
timestamp 1698175906
transform 1 0 7392 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _154_
timestamp 1698175906
transform -1 0 8400 0 -1 10192
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _155_
timestamp 1698175906
transform 1 0 7896 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _156_
timestamp 1698175906
transform 1 0 7896 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _157_
timestamp 1698175906
transform -1 0 8960 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _158_
timestamp 1698175906
transform 1 0 7728 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _159_
timestamp 1698175906
transform 1 0 7504 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _160_
timestamp 1698175906
transform 1 0 7280 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _161_
timestamp 1698175906
transform -1 0 7168 0 1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _162_
timestamp 1698175906
transform 1 0 9912 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _163_
timestamp 1698175906
transform -1 0 8512 0 -1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _164_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8736 0 -1 12544
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nor4_2  _165_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9240 0 -1 12544
box -43 -43 1051 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _166_
timestamp 1698175906
transform -1 0 8400 0 1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _167_
timestamp 1698175906
transform 1 0 6664 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _168_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 6888 0 1 11760
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _169_
timestamp 1698175906
transform 1 0 9184 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _170_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11872 0 -1 10976
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _171_
timestamp 1698175906
transform 1 0 9296 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _172_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10864 0 -1 10976
box -43 -43 1051 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _173_
timestamp 1698175906
transform 1 0 11200 0 1 11760
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_4  _174_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8904 0 -1 9408
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _175_
timestamp 1698175906
transform 1 0 8288 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _176_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9240 0 1 7840
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _177_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10472 0 1 8624
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _178_
timestamp 1698175906
transform 1 0 10584 0 1 9408
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _179_
timestamp 1698175906
transform 1 0 8960 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _180_
timestamp 1698175906
transform 1 0 9128 0 -1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _181_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10024 0 1 9408
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _182_
timestamp 1698175906
transform 1 0 10024 0 -1 7840
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _183_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9296 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _184_
timestamp 1698175906
transform -1 0 13552 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _185_
timestamp 1698175906
transform 1 0 10584 0 1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_2  _186_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9184 0 1 9408
box -43 -43 883 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _187_
timestamp 1698175906
transform -1 0 13104 0 1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _188_
timestamp 1698175906
transform 1 0 12040 0 1 12544
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _189_
timestamp 1698175906
transform -1 0 13776 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _190_
timestamp 1698175906
transform 1 0 12656 0 -1 12544
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _191_
timestamp 1698175906
transform 1 0 10584 0 -1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _192_
timestamp 1698175906
transform -1 0 10528 0 -1 13328
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _193_
timestamp 1698175906
transform -1 0 10248 0 1 13328
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _194_
timestamp 1698175906
transform 1 0 9520 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _195_
timestamp 1698175906
transform -1 0 9912 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _196_
timestamp 1698175906
transform -1 0 10864 0 1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _197_
timestamp 1698175906
transform 1 0 9408 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _198_
timestamp 1698175906
transform 1 0 8624 0 -1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _199_
timestamp 1698175906
transform 1 0 13496 0 -1 10192
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _200_
timestamp 1698175906
transform 1 0 12824 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _201_
timestamp 1698175906
transform 1 0 11816 0 1 10192
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _202_
timestamp 1698175906
transform -1 0 13720 0 1 7840
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _203_
timestamp 1698175906
transform -1 0 13328 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _204_
timestamp 1698175906
transform -1 0 9576 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _205_
timestamp 1698175906
transform -1 0 9352 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _206_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9912 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _207_
timestamp 1698175906
transform -1 0 8512 0 -1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _208_
timestamp 1698175906
transform 1 0 10640 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _209_
timestamp 1698175906
transform 1 0 12712 0 1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _210_
timestamp 1698175906
transform -1 0 12880 0 -1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _211_
timestamp 1698175906
transform 1 0 8792 0 1 9408
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _212_
timestamp 1698175906
transform 1 0 9912 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _213_
timestamp 1698175906
transform 1 0 11144 0 -1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _214_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10472 0 1 7056
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _215_
timestamp 1698175906
transform -1 0 10920 0 1 6272
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _216_
timestamp 1698175906
transform 1 0 10472 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _217_
timestamp 1698175906
transform 1 0 11760 0 -1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _218_
timestamp 1698175906
transform -1 0 11088 0 1 7840
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _219_
timestamp 1698175906
transform -1 0 10304 0 -1 7056
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _220_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 10472 0 1 7840
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _221_
timestamp 1698175906
transform -1 0 10024 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _222_
timestamp 1698175906
transform 1 0 11144 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor3_1  _223_
timestamp 1698175906
transform -1 0 11144 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _224_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12768 0 -1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _225_
timestamp 1698175906
transform 1 0 12768 0 1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _226_
timestamp 1698175906
transform 1 0 12768 0 -1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _227_
timestamp 1698175906
transform 1 0 4928 0 1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _228_
timestamp 1698175906
transform 1 0 4928 0 1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _229_
timestamp 1698175906
transform 1 0 5992 0 -1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _230_
timestamp 1698175906
transform 1 0 5768 0 -1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _231_
timestamp 1698175906
transform -1 0 7504 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _232_
timestamp 1698175906
transform 1 0 6888 0 -1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _233_
timestamp 1698175906
transform -1 0 7000 0 -1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _234_
timestamp 1698175906
transform 1 0 10808 0 1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _235_
timestamp 1698175906
transform 1 0 6888 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _236_
timestamp 1698175906
transform 1 0 12544 0 -1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _237_
timestamp 1698175906
transform 1 0 12600 0 1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _238_
timestamp 1698175906
transform 1 0 9296 0 -1 14112
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _239_
timestamp 1698175906
transform 1 0 8288 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _240_
timestamp 1698175906
transform 1 0 12768 0 1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _241_
timestamp 1698175906
transform 1 0 12712 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _242_
timestamp 1698175906
transform 1 0 7336 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _243_
timestamp 1698175906
transform 1 0 11928 0 1 6272
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _244_
timestamp 1698175906
transform 1 0 10136 0 -1 6272
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _245_
timestamp 1698175906
transform 1 0 10696 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _246_
timestamp 1698175906
transform 1 0 8568 0 1 6272
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _247_
timestamp 1698175906
transform 1 0 10584 0 -1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _251_
timestamp 1698175906
transform 1 0 14168 0 -1 13328
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _252_
timestamp 1698175906
transform 1 0 14504 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _253_
timestamp 1698175906
transform -1 0 11256 0 -1 14112
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__160__A1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7840 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__200__A1
timestamp 1698175906
transform -1 0 12824 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__201__A1
timestamp 1698175906
transform -1 0 11984 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__224__CLK
timestamp 1698175906
transform -1 0 12768 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__225__CLK
timestamp 1698175906
transform 1 0 12656 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__226__CLK
timestamp 1698175906
transform 1 0 12656 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__227__CLK
timestamp 1698175906
transform -1 0 6776 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__227__D
timestamp 1698175906
transform 1 0 6552 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__228__CLK
timestamp 1698175906
transform 1 0 6776 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__229__CLK
timestamp 1698175906
transform 1 0 7728 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__230__CLK
timestamp 1698175906
transform -1 0 7616 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__231__CLK
timestamp 1698175906
transform 1 0 7616 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__232__CLK
timestamp 1698175906
transform 1 0 8736 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__233__CLK
timestamp 1698175906
transform 1 0 7112 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__234__CLK
timestamp 1698175906
transform 1 0 12544 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__235__CLK
timestamp 1698175906
transform 1 0 8736 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__236__CLK
timestamp 1698175906
transform 1 0 12432 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__237__CLK
timestamp 1698175906
transform 1 0 11928 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__238__CLK
timestamp 1698175906
transform -1 0 11480 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__239__CLK
timestamp 1698175906
transform 1 0 10360 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__240__CLK
timestamp 1698175906
transform 1 0 12656 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__241__CLK
timestamp 1698175906
transform 1 0 12320 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__242__CLK
timestamp 1698175906
transform 1 0 9072 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__243__CLK
timestamp 1698175906
transform 1 0 11816 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__244__CLK
timestamp 1698175906
transform 1 0 11872 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__245__CLK
timestamp 1698175906
transform 1 0 12432 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__246__CLK
timestamp 1698175906
transform 1 0 10304 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__247__CLK
timestamp 1698175906
transform 1 0 12320 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform 1 0 8848 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8960 0 -1 10192
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform 1 0 9408 0 -1 8624
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 9296 0 -1 11760
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_36 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 2688 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_44 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 3136 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_48 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 3360 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_0_53
timestamp 1698175906
transform 1 0 3640 0 1 1568
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_61
timestamp 1698175906
transform 1 0 4088 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_65 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 4312 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_67
timestamp 1698175906
transform 1 0 4424 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 4592 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 6496 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_138
timestamp 1698175906
transform 1 0 8400 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_142
timestamp 1698175906
transform 1 0 8624 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_198
timestamp 1698175906
transform 1 0 11760 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_202
timestamp 1698175906
transform 1 0 11984 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_232
timestamp 1698175906
transform 1 0 13664 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_236
timestamp 1698175906
transform 1 0 13888 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_266
timestamp 1698175906
transform 1 0 15568 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_270
timestamp 1698175906
transform 1 0 15792 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 16016 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 17920 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 19824 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 20048 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348
timestamp 1698175906
transform 1 0 20160 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 4368 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 4704 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 8288 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_142
timestamp 1698175906
transform 1 0 8624 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_144
timestamp 1698175906
transform 1 0 8736 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_171
timestamp 1698175906
transform 1 0 10248 0 -1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_203
timestamp 1698175906
transform 1 0 12040 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_207
timestamp 1698175906
transform 1 0 12264 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698175906
transform 1 0 12376 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_238
timestamp 1698175906
transform 1 0 14000 0 -1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_270
timestamp 1698175906
transform 1 0 15792 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_278
timestamp 1698175906
transform 1 0 16240 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 16464 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 20048 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 20160 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 784 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 2576 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 2744 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 6328 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 6664 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 10248 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698175906
transform 1 0 10584 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 14168 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 14504 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 18088 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 18424 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 784 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 4368 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 4704 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 8288 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 8624 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 12208 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 12544 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 16128 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 16464 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 20048 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 20160 0 -1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 784 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 2576 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 2744 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 6328 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 6664 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 10248 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 10584 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 14168 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 14504 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 18088 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 18424 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 784 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 4368 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 4704 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 8288 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 8624 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 12208 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 12544 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 16128 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 16464 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 20048 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 20160 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 784 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 2576 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 2744 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 6328 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 6664 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 10248 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 10584 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 14168 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 14504 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 18088 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 18424 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 784 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 4368 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 4704 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 8288 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 8624 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 12208 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 12544 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 16128 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 16464 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 20048 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 20160 0 -1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 784 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 2576 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 2744 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 6328 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 6664 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 10248 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 10584 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 14168 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 14504 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 18088 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 18424 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 784 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 4368 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 4704 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 8288 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 8624 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 12208 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 12544 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 16128 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 16464 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 20048 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 20160 0 -1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 784 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 2576 0 1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 2744 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 6328 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 6664 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 10248 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 10584 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 14168 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 14504 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 18088 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 18424 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 784 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 4368 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 4704 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 8288 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_11_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 -1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_158
timestamp 1698175906
transform 1 0 9520 0 -1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_166
timestamp 1698175906
transform 1 0 9968 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_168
timestamp 1698175906
transform 1 0 10080 0 -1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_198
timestamp 1698175906
transform 1 0 11760 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_11_202
timestamp 1698175906
transform 1 0 11984 0 -1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 12544 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 16128 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 16464 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 20048 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 20160 0 -1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 784 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 2576 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 2744 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 6328 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_107
timestamp 1698175906
transform 1 0 6664 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_139
timestamp 1698175906
transform 1 0 8456 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_170
timestamp 1698175906
transform 1 0 10192 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_174
timestamp 1698175906
transform 1 0 10416 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_183
timestamp 1698175906
transform 1 0 10920 0 1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_230
timestamp 1698175906
transform 1 0 13552 0 1 6272
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_238
timestamp 1698175906
transform 1 0 14000 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_242
timestamp 1698175906
transform 1 0 14224 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_244
timestamp 1698175906
transform 1 0 14336 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 14504 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 18088 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 18424 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 784 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 4368 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_72
timestamp 1698175906
transform 1 0 4704 0 -1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_104
timestamp 1698175906
transform 1 0 6496 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_120
timestamp 1698175906
transform 1 0 7392 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_128
timestamp 1698175906
transform 1 0 7840 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_132
timestamp 1698175906
transform 1 0 8064 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_142
timestamp 1698175906
transform 1 0 8624 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_146
timestamp 1698175906
transform 1 0 8848 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_155
timestamp 1698175906
transform 1 0 9352 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_172
timestamp 1698175906
transform 1 0 10304 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_180
timestamp 1698175906
transform 1 0 10752 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_184
timestamp 1698175906
transform 1 0 10976 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_186
timestamp 1698175906
transform 1 0 11088 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_193
timestamp 1698175906
transform 1 0 11480 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_209
timestamp 1698175906
transform 1 0 12376 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_218
timestamp 1698175906
transform 1 0 12880 0 -1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_250
timestamp 1698175906
transform 1 0 14672 0 -1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_266
timestamp 1698175906
transform 1 0 15568 0 -1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_274
timestamp 1698175906
transform 1 0 16016 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_278
timestamp 1698175906
transform 1 0 16240 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 16464 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 20048 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 20160 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 784 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 2576 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 2744 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 6328 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_107
timestamp 1698175906
transform 1 0 6664 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_115
timestamp 1698175906
transform 1 0 7112 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_148
timestamp 1698175906
transform 1 0 8960 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_152
timestamp 1698175906
transform 1 0 9184 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_160
timestamp 1698175906
transform 1 0 9632 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_164
timestamp 1698175906
transform 1 0 9856 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_177
timestamp 1698175906
transform 1 0 10584 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_208
timestamp 1698175906
transform 1 0 12320 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_212
timestamp 1698175906
transform 1 0 12544 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_214
timestamp 1698175906
transform 1 0 12656 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_221
timestamp 1698175906
transform 1 0 13048 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_237
timestamp 1698175906
transform 1 0 13944 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 14504 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 18088 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 18424 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 784 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 4368 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_72
timestamp 1698175906
transform 1 0 4704 0 -1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_104
timestamp 1698175906
transform 1 0 6496 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_108
timestamp 1698175906
transform 1 0 6720 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_110
timestamp 1698175906
transform 1 0 6832 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_142
timestamp 1698175906
transform 1 0 8624 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_154
timestamp 1698175906
transform 1 0 9296 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_156
timestamp 1698175906
transform 1 0 9408 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_165
timestamp 1698175906
transform 1 0 9912 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_174
timestamp 1698175906
transform 1 0 10416 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_190
timestamp 1698175906
transform 1 0 11312 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_204
timestamp 1698175906
transform 1 0 12096 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_212
timestamp 1698175906
transform 1 0 12544 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_214
timestamp 1698175906
transform 1 0 12656 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_244
timestamp 1698175906
transform 1 0 14336 0 -1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_276
timestamp 1698175906
transform 1 0 16128 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 16464 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698175906
transform 1 0 20048 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698175906
transform 1 0 20160 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 784 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 2576 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 2744 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 6328 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_107
timestamp 1698175906
transform 1 0 6664 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_139
timestamp 1698175906
transform 1 0 8456 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_159
timestamp 1698175906
transform 1 0 9576 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_163
timestamp 1698175906
transform 1 0 9800 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_165
timestamp 1698175906
transform 1 0 9912 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_186
timestamp 1698175906
transform 1 0 11088 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_226
timestamp 1698175906
transform 1 0 13328 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_233
timestamp 1698175906
transform 1 0 13720 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_241
timestamp 1698175906
transform 1 0 14168 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 14504 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 18088 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_317
timestamp 1698175906
transform 1 0 18424 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_321
timestamp 1698175906
transform 1 0 18648 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698175906
transform 1 0 784 0 -1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698175906
transform 1 0 4368 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_72
timestamp 1698175906
transform 1 0 4704 0 -1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_88
timestamp 1698175906
transform 1 0 5600 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_92
timestamp 1698175906
transform 1 0 5824 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_94
timestamp 1698175906
transform 1 0 5936 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_124
timestamp 1698175906
transform 1 0 7616 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_128
timestamp 1698175906
transform 1 0 7840 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_132
timestamp 1698175906
transform 1 0 8064 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_134
timestamp 1698175906
transform 1 0 8176 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_139
timestamp 1698175906
transform 1 0 8456 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_146
timestamp 1698175906
transform 1 0 8848 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_150
timestamp 1698175906
transform 1 0 9072 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_206
timestamp 1698175906
transform 1 0 12208 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_212
timestamp 1698175906
transform 1 0 12544 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_245
timestamp 1698175906
transform 1 0 14392 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_277
timestamp 1698175906
transform 1 0 16184 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_279
timestamp 1698175906
transform 1 0 16296 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_282
timestamp 1698175906
transform 1 0 16464 0 -1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_346
timestamp 1698175906
transform 1 0 20048 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_348
timestamp 1698175906
transform 1 0 20160 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698175906
transform 1 0 784 0 1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 2576 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698175906
transform 1 0 2744 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698175906
transform 1 0 6328 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_107
timestamp 1698175906
transform 1 0 6664 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_115
timestamp 1698175906
transform 1 0 7112 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_119
timestamp 1698175906
transform 1 0 7336 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_126
timestamp 1698175906
transform 1 0 7728 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_128
timestamp 1698175906
transform 1 0 7840 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_135
timestamp 1698175906
transform 1 0 8232 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_177
timestamp 1698175906
transform 1 0 10584 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_192
timestamp 1698175906
transform 1 0 11424 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_194
timestamp 1698175906
transform 1 0 11536 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_18_201
timestamp 1698175906
transform 1 0 11928 0 1 8624
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_217
timestamp 1698175906
transform 1 0 12824 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_219
timestamp 1698175906
transform 1 0 12936 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_236
timestamp 1698175906
transform 1 0 13888 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_244
timestamp 1698175906
transform 1 0 14336 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698175906
transform 1 0 14504 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698175906
transform 1 0 18088 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_317
timestamp 1698175906
transform 1 0 18424 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_321
timestamp 1698175906
transform 1 0 18648 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698175906
transform 1 0 784 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698175906
transform 1 0 4368 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_72
timestamp 1698175906
transform 1 0 4704 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_88
timestamp 1698175906
transform 1 0 5600 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_90
timestamp 1698175906
transform 1 0 5712 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_120
timestamp 1698175906
transform 1 0 7392 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_142
timestamp 1698175906
transform 1 0 8624 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_146
timestamp 1698175906
transform 1 0 8848 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_173
timestamp 1698175906
transform 1 0 10360 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_183
timestamp 1698175906
transform 1 0 10920 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_198
timestamp 1698175906
transform 1 0 11760 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_206
timestamp 1698175906
transform 1 0 12208 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_212
timestamp 1698175906
transform 1 0 12544 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_245
timestamp 1698175906
transform 1 0 14392 0 -1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_277
timestamp 1698175906
transform 1 0 16184 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_279
timestamp 1698175906
transform 1 0 16296 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_282
timestamp 1698175906
transform 1 0 16464 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_346
timestamp 1698175906
transform 1 0 20048 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_348
timestamp 1698175906
transform 1 0 20160 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 784 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 2576 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698175906
transform 1 0 2744 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698175906
transform 1 0 6328 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_107
timestamp 1698175906
transform 1 0 6664 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_123
timestamp 1698175906
transform 1 0 7560 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_125
timestamp 1698175906
transform 1 0 7672 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_140
timestamp 1698175906
transform 1 0 8512 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_144
timestamp 1698175906
transform 1 0 8736 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_174
timestamp 1698175906
transform 1 0 10416 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_205
timestamp 1698175906
transform 1 0 12152 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_207
timestamp 1698175906
transform 1 0 12264 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_214
timestamp 1698175906
transform 1 0 12656 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_226
timestamp 1698175906
transform 1 0 13328 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_235
timestamp 1698175906
transform 1 0 13832 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_243
timestamp 1698175906
transform 1 0 14280 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698175906
transform 1 0 14504 0 1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698175906
transform 1 0 18088 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_317
timestamp 1698175906
transform 1 0 18424 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_321
timestamp 1698175906
transform 1 0 18648 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698175906
transform 1 0 784 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698175906
transform 1 0 4368 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_72
timestamp 1698175906
transform 1 0 4704 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_104
timestamp 1698175906
transform 1 0 6496 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_106
timestamp 1698175906
transform 1 0 6608 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_109
timestamp 1698175906
transform 1 0 6776 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_117
timestamp 1698175906
transform 1 0 7224 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_119
timestamp 1698175906
transform 1 0 7336 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_138
timestamp 1698175906
transform 1 0 8400 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_198
timestamp 1698175906
transform 1 0 11760 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_202
timestamp 1698175906
transform 1 0 11984 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_212
timestamp 1698175906
transform 1 0 12544 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_214
timestamp 1698175906
transform 1 0 12656 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_225
timestamp 1698175906
transform 1 0 13272 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_236
timestamp 1698175906
transform 1 0 13888 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_268
timestamp 1698175906
transform 1 0 15680 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_276
timestamp 1698175906
transform 1 0 16128 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_282
timestamp 1698175906
transform 1 0 16464 0 -1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_346
timestamp 1698175906
transform 1 0 20048 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_348
timestamp 1698175906
transform 1 0 20160 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 784 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 2576 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_37
timestamp 1698175906
transform 1 0 2744 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_69
timestamp 1698175906
transform 1 0 4536 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_73
timestamp 1698175906
transform 1 0 4760 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_75
timestamp 1698175906
transform 1 0 4872 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_107
timestamp 1698175906
transform 1 0 6664 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_137
timestamp 1698175906
transform 1 0 8344 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_145
timestamp 1698175906
transform 1 0 8792 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_161
timestamp 1698175906
transform 1 0 9688 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_173
timestamp 1698175906
transform 1 0 10360 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_183
timestamp 1698175906
transform 1 0 10920 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_196
timestamp 1698175906
transform 1 0 11648 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_198
timestamp 1698175906
transform 1 0 11760 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_206
timestamp 1698175906
transform 1 0 12208 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_253
timestamp 1698175906
transform 1 0 14840 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_285
timestamp 1698175906
transform 1 0 16632 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_301
timestamp 1698175906
transform 1 0 17528 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_309
timestamp 1698175906
transform 1 0 17976 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_313
timestamp 1698175906
transform 1 0 18200 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_317
timestamp 1698175906
transform 1 0 18424 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_321
timestamp 1698175906
transform 1 0 18648 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698175906
transform 1 0 784 0 -1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698175906
transform 1 0 4368 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_72
timestamp 1698175906
transform 1 0 4704 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_104
timestamp 1698175906
transform 1 0 6496 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_107
timestamp 1698175906
transform 1 0 6664 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_111
timestamp 1698175906
transform 1 0 6888 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_117
timestamp 1698175906
transform 1 0 7224 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_119
timestamp 1698175906
transform 1 0 7336 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_126
timestamp 1698175906
transform 1 0 7728 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_128
timestamp 1698175906
transform 1 0 7840 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_139
timestamp 1698175906
transform 1 0 8456 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_166
timestamp 1698175906
transform 1 0 9968 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_168
timestamp 1698175906
transform 1 0 10080 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_175
timestamp 1698175906
transform 1 0 10472 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_212
timestamp 1698175906
transform 1 0 12544 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_216
timestamp 1698175906
transform 1 0 12768 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_232
timestamp 1698175906
transform 1 0 13664 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_264
timestamp 1698175906
transform 1 0 15456 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698175906
transform 1 0 16464 0 -1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_314
timestamp 1698175906
transform 1 0 18256 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_322
timestamp 1698175906
transform 1 0 18704 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698175906
transform 1 0 784 0 1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 2576 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_37
timestamp 1698175906
transform 1 0 2744 0 1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_69
timestamp 1698175906
transform 1 0 4536 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_73
timestamp 1698175906
transform 1 0 4760 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_75
timestamp 1698175906
transform 1 0 4872 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_107
timestamp 1698175906
transform 1 0 6664 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_123
timestamp 1698175906
transform 1 0 7560 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_155
timestamp 1698175906
transform 1 0 9352 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_165
timestamp 1698175906
transform 1 0 9912 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_174
timestamp 1698175906
transform 1 0 10416 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_177
timestamp 1698175906
transform 1 0 10584 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_210
timestamp 1698175906
transform 1 0 12432 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_214
timestamp 1698175906
transform 1 0 12656 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698175906
transform 1 0 14504 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 18088 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_317
timestamp 1698175906
transform 1 0 18424 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698175906
transform 1 0 18648 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2
timestamp 1698175906
transform 1 0 784 0 -1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_66
timestamp 1698175906
transform 1 0 4368 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_72
timestamp 1698175906
transform 1 0 4704 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_80
timestamp 1698175906
transform 1 0 5152 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_113
timestamp 1698175906
transform 1 0 7000 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_117
timestamp 1698175906
transform 1 0 7224 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_126
timestamp 1698175906
transform 1 0 7728 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_130
timestamp 1698175906
transform 1 0 7952 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_134
timestamp 1698175906
transform 1 0 8176 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_204
timestamp 1698175906
transform 1 0 12096 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_208
timestamp 1698175906
transform 1 0 12320 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_25_212
timestamp 1698175906
transform 1 0 12544 0 -1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_236
timestamp 1698175906
transform 1 0 13888 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_268
timestamp 1698175906
transform 1 0 15680 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_276
timestamp 1698175906
transform 1 0 16128 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_282
timestamp 1698175906
transform 1 0 16464 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_314
timestamp 1698175906
transform 1 0 18256 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_322
timestamp 1698175906
transform 1 0 18704 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_2
timestamp 1698175906
transform 1 0 784 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 2576 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698175906
transform 1 0 2744 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698175906
transform 1 0 6328 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_130
timestamp 1698175906
transform 1 0 7952 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_162
timestamp 1698175906
transform 1 0 9744 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_164
timestamp 1698175906
transform 1 0 9856 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_171
timestamp 1698175906
transform 1 0 10248 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_182
timestamp 1698175906
transform 1 0 10864 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_186
timestamp 1698175906
transform 1 0 11088 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_198
timestamp 1698175906
transform 1 0 11760 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_214
timestamp 1698175906
transform 1 0 12656 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_216
timestamp 1698175906
transform 1 0 12768 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_222
timestamp 1698175906
transform 1 0 13104 0 1 11760
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_238
timestamp 1698175906
transform 1 0 14000 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_242
timestamp 1698175906
transform 1 0 14224 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_244
timestamp 1698175906
transform 1 0 14336 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 14504 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 18088 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_317
timestamp 1698175906
transform 1 0 18424 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698175906
transform 1 0 784 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698175906
transform 1 0 4368 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_72
timestamp 1698175906
transform 1 0 4704 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_88
timestamp 1698175906
transform 1 0 5600 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_92
timestamp 1698175906
transform 1 0 5824 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_122
timestamp 1698175906
transform 1 0 7504 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_130
timestamp 1698175906
transform 1 0 7952 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_138
timestamp 1698175906
transform 1 0 8400 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_142
timestamp 1698175906
transform 1 0 8624 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_171
timestamp 1698175906
transform 1 0 10248 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_175
timestamp 1698175906
transform 1 0 10472 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_183
timestamp 1698175906
transform 1 0 10920 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_199
timestamp 1698175906
transform 1 0 11816 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_207
timestamp 1698175906
transform 1 0 12264 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_209
timestamp 1698175906
transform 1 0 12376 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_212
timestamp 1698175906
transform 1 0 12544 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_224
timestamp 1698175906
transform 1 0 13216 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_228
timestamp 1698175906
transform 1 0 13440 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_234
timestamp 1698175906
transform 1 0 13776 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_266
timestamp 1698175906
transform 1 0 15568 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_274
timestamp 1698175906
transform 1 0 16016 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_278
timestamp 1698175906
transform 1 0 16240 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_282
timestamp 1698175906
transform 1 0 16464 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_346
timestamp 1698175906
transform 1 0 20048 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_348
timestamp 1698175906
transform 1 0 20160 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_28
timestamp 1698175906
transform 1 0 2240 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_32
timestamp 1698175906
transform 1 0 2464 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 2576 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 2744 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 6328 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_107
timestamp 1698175906
transform 1 0 6664 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_109
timestamp 1698175906
transform 1 0 6776 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_116
timestamp 1698175906
transform 1 0 7168 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_138
timestamp 1698175906
transform 1 0 8400 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_170
timestamp 1698175906
transform 1 0 10192 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_174
timestamp 1698175906
transform 1 0 10416 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_177
timestamp 1698175906
transform 1 0 10584 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_195
timestamp 1698175906
transform 1 0 11592 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_199
timestamp 1698175906
transform 1 0 11816 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_242
timestamp 1698175906
transform 1 0 14224 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_244
timestamp 1698175906
transform 1 0 14336 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 14504 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 18088 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_317
timestamp 1698175906
transform 1 0 18424 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_321
timestamp 1698175906
transform 1 0 18648 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_28
timestamp 1698175906
transform 1 0 2240 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_60
timestamp 1698175906
transform 1 0 4032 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_68
timestamp 1698175906
transform 1 0 4480 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_72
timestamp 1698175906
transform 1 0 4704 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_104
timestamp 1698175906
transform 1 0 6496 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_108
timestamp 1698175906
transform 1 0 6720 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_110
timestamp 1698175906
transform 1 0 6832 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_142
timestamp 1698175906
transform 1 0 8624 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_146
timestamp 1698175906
transform 1 0 8848 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_154
timestamp 1698175906
transform 1 0 9296 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_164
timestamp 1698175906
transform 1 0 9856 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_166
timestamp 1698175906
transform 1 0 9968 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_176
timestamp 1698175906
transform 1 0 10528 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_206
timestamp 1698175906
transform 1 0 12208 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_247
timestamp 1698175906
transform 1 0 14504 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_279
timestamp 1698175906
transform 1 0 16296 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_282
timestamp 1698175906
transform 1 0 16464 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_314
timestamp 1698175906
transform 1 0 18256 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_322
timestamp 1698175906
transform 1 0 18704 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_2
timestamp 1698175906
transform 1 0 784 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 2576 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 2744 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 6328 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_107
timestamp 1698175906
transform 1 0 6664 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_123
timestamp 1698175906
transform 1 0 7560 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_131
timestamp 1698175906
transform 1 0 8008 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_135
timestamp 1698175906
transform 1 0 8232 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_171
timestamp 1698175906
transform 1 0 10248 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_182
timestamp 1698175906
transform 1 0 10864 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_198
timestamp 1698175906
transform 1 0 11760 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_206
timestamp 1698175906
transform 1 0 12208 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_212
timestamp 1698175906
transform 1 0 12544 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_220
timestamp 1698175906
transform 1 0 12992 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_224
timestamp 1698175906
transform 1 0 13216 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_230
timestamp 1698175906
transform 1 0 13552 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_238
timestamp 1698175906
transform 1 0 14000 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_242
timestamp 1698175906
transform 1 0 14224 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_244
timestamp 1698175906
transform 1 0 14336 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 14504 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 18088 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_317
timestamp 1698175906
transform 1 0 18424 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_321
timestamp 1698175906
transform 1 0 18648 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 784 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 4368 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_72
timestamp 1698175906
transform 1 0 4704 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_136
timestamp 1698175906
transform 1 0 8288 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_142
timestamp 1698175906
transform 1 0 8624 0 -1 14112
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_150
timestamp 1698175906
transform 1 0 9072 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_189
timestamp 1698175906
transform 1 0 11256 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_193
timestamp 1698175906
transform 1 0 11480 0 -1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_209
timestamp 1698175906
transform 1 0 12376 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698175906
transform 1 0 12544 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698175906
transform 1 0 16128 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 16464 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 20048 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 20160 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 784 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 2576 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 2744 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 6328 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_107
timestamp 1698175906
transform 1 0 6664 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_171
timestamp 1698175906
transform 1 0 10248 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698175906
transform 1 0 10584 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698175906
transform 1 0 14168 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 14504 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 18088 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 18424 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 784 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 4368 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 4704 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 8288 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 8624 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 12208 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 12544 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 16128 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 16464 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 20048 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 20160 0 -1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 784 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 2576 0 1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 2744 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 6328 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 6664 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 10248 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 10584 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 14168 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 14504 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 18088 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 18424 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 784 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 4368 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 4704 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 8288 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 8624 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 12208 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 12544 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 16128 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 16464 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 20048 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 20160 0 -1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 784 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 2576 0 1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 2744 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 6328 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 6664 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 10248 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 10584 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 14168 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 14504 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 18088 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 18424 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 784 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 4368 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 4704 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 8288 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 8624 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 12208 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 12544 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 16128 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 16464 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 20048 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 20160 0 -1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 784 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 2576 0 1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 2744 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 6328 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 6664 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 10248 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 10584 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 14168 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 14504 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 18088 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 18424 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 784 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 4368 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 4704 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 8288 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 8624 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 12208 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 12544 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 16128 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 16464 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 20048 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 20160 0 -1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 784 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 2576 0 1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 2744 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 6328 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 6664 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 10248 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 10584 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 14168 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 14504 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 18088 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_40_317
timestamp 1698175906
transform 1 0 18424 0 1 17248
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_40_333
timestamp 1698175906
transform 1 0 19320 0 1 17248
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_341
timestamp 1698175906
transform 1 0 19768 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 784 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 4368 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 4704 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 8288 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 8624 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 12208 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 12544 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 16128 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 16464 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 20048 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 20160 0 -1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 784 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 2576 0 1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 2744 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 6328 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698175906
transform 1 0 6664 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698175906
transform 1 0 10248 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698175906
transform 1 0 10584 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 14168 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 14504 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 18088 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 18424 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 784 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 4368 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 4704 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 8288 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_142
timestamp 1698175906
transform 1 0 8624 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_144
timestamp 1698175906
transform 1 0 8736 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_171
timestamp 1698175906
transform 1 0 10248 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_201
timestamp 1698175906
transform 1 0 11928 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 12376 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_212
timestamp 1698175906
transform 1 0 12544 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_276
timestamp 1698175906
transform 1 0 16128 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 16464 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 20048 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 20160 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 784 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 2688 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 4592 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 6496 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_138
timestamp 1698175906
transform 1 0 8400 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_142
timestamp 1698175906
transform 1 0 8624 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_172
timestamp 1698175906
transform 1 0 10304 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_232
timestamp 1698175906
transform 1 0 13664 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 13888 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_240
timestamp 1698175906
transform 1 0 14112 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 16016 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 17920 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 19824 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 20048 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 20160 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita25_24 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19992 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita25_25
timestamp 1698175906
transform 1 0 10416 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita25_26
timestamp 1698175906
transform -1 0 3640 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12544 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform 1 0 8792 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform 1 0 10304 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform 1 0 18760 0 1 12544
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform 1 0 10472 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform 1 0 18760 0 -1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform -1 0 10192 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform 1 0 12208 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform 1 0 18760 0 -1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform 1 0 18760 0 -1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform 1 0 18760 0 1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform -1 0 2240 0 1 12544
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform 1 0 8736 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform 1 0 14112 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform 1 0 8792 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform -1 0 2240 0 -1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform 1 0 18760 0 1 10192
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform 1 0 18760 0 1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform 1 0 10640 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform 1 0 18760 0 1 7840
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform 1 0 18760 0 1 9408
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform 1 0 18760 0 1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform 1 0 12208 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 20328 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 20328 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 20328 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 20328 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 20328 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 20328 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 20328 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 672 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 20328 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 672 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 20328 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 672 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 20328 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 672 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 20328 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 672 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 20328 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 672 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 20328 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 672 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 20328 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 672 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 20328 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 672 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 20328 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 672 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 20328 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 672 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 20328 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 672 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 20328 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 672 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 20328 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 672 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 20328 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 672 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 20328 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 672 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 20328 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 672 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 20328 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 672 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 20328 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 672 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 20328 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 672 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 20328 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 672 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 20328 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 672 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 20328 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 672 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 20328 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 672 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 20328 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 672 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 20328 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 672 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 20328 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 672 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 20328 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 672 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 20328 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 672 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 20328 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 672 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 20328 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 672 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 20328 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 672 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 20328 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 672 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 20328 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 672 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 20328 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 672 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 20328 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 672 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 20328 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 672 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 20328 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 672 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 20328 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 2576 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 4480 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 6384 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 8288 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 10192 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 12096 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 14000 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 15904 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 17808 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 19712 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 4592 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 8512 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 12432 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 16352 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 6552 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 10472 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 14392 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 18312 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 4592 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 8512 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 12432 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 16352 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 6552 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 10472 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 14392 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 18312 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 4592 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 8512 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 12432 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 16352 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 6552 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 10472 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 14392 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 18312 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 4592 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 8512 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 12432 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 16352 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 2632 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 6552 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 10472 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 14392 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 18312 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 4592 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 8512 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 12432 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 16352 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 2632 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 6552 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 10472 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 14392 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 18312 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 4592 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 8512 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 12432 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 16352 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 2632 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 6552 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 10472 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 14392 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 18312 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 4592 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 8512 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 12432 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 16352 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 2632 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 6552 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 10472 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 14392 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 18312 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 4592 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 8512 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 12432 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 16352 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 2632 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 6552 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 10472 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 14392 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 18312 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 4592 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 8512 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 12432 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 16352 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 2632 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 6552 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 10472 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 14392 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 18312 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 4592 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 8512 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 12432 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 16352 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 2632 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 6552 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 10472 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 14392 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 18312 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 4592 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 8512 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 12432 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 16352 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 2632 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 6552 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 10472 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 14392 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 18312 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 4592 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 8512 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 12432 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 16352 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 2632 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 6552 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 10472 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 14392 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 18312 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 4592 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 8512 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 12432 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 16352 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 2632 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 6552 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 10472 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 14392 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 18312 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 4592 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 8512 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 12432 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 16352 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 2632 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 6552 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 10472 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 14392 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 18312 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 4592 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 8512 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 12432 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 16352 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 2632 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 6552 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 10472 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 14392 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 18312 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 4592 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 8512 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 12432 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 16352 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 2632 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 6552 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 10472 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 14392 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 18312 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 4592 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 8512 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 12432 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 16352 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 2632 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 6552 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 10472 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 14392 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 18312 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 4592 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 8512 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 12432 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 16352 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 2632 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 6552 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 10472 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 14392 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 18312 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 4592 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 8512 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 12432 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 16352 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 2632 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 6552 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 10472 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 14392 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 18312 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 4592 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 8512 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 12432 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 16352 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 2632 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 6552 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 10472 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 14392 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 18312 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 4592 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 8512 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 12432 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 16352 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 2632 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 6552 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 10472 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 14392 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 18312 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 4592 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 8512 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 12432 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 16352 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 2576 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 4480 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 6384 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 8288 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 10192 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 12096 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 14000 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 15904 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 17808 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 19712 0 1 18816
box -43 -43 155 435
<< labels >>
flabel metal3 s 0 13776 400 13832 0 FreeSans 224 0 0 0 clk
port 0 nsew signal input
flabel metal3 s 20600 17136 21000 17192 0 FreeSans 224 0 0 0 segm[0]
port 1 nsew signal tristate
flabel metal2 s 12096 0 12152 400 0 FreeSans 224 90 0 0 segm[10]
port 2 nsew signal tristate
flabel metal2 s 8736 0 8792 400 0 FreeSans 224 90 0 0 segm[11]
port 3 nsew signal tristate
flabel metal2 s 10080 0 10136 400 0 FreeSans 224 90 0 0 segm[12]
port 4 nsew signal tristate
flabel metal3 s 20600 12432 21000 12488 0 FreeSans 224 0 0 0 segm[13]
port 5 nsew signal tristate
flabel metal2 s 11088 20600 11144 21000 0 FreeSans 224 90 0 0 segm[1]
port 6 nsew signal tristate
flabel metal2 s 10416 20600 10472 21000 0 FreeSans 224 90 0 0 segm[2]
port 7 nsew signal tristate
flabel metal3 s 20600 10416 21000 10472 0 FreeSans 224 0 0 0 segm[3]
port 8 nsew signal tristate
flabel metal2 s 3360 0 3416 400 0 FreeSans 224 90 0 0 segm[4]
port 9 nsew signal tristate
flabel metal2 s 9744 20600 9800 21000 0 FreeSans 224 90 0 0 segm[5]
port 10 nsew signal tristate
flabel metal2 s 11424 0 11480 400 0 FreeSans 224 90 0 0 segm[6]
port 11 nsew signal tristate
flabel metal3 s 20600 11424 21000 11480 0 FreeSans 224 0 0 0 segm[7]
port 12 nsew signal tristate
flabel metal3 s 20600 13440 21000 13496 0 FreeSans 224 0 0 0 segm[8]
port 13 nsew signal tristate
flabel metal3 s 20600 13104 21000 13160 0 FreeSans 224 0 0 0 segm[9]
port 14 nsew signal tristate
flabel metal3 s 0 12432 400 12488 0 FreeSans 224 0 0 0 sel[0]
port 15 nsew signal tristate
flabel metal2 s 9072 0 9128 400 0 FreeSans 224 90 0 0 sel[10]
port 16 nsew signal tristate
flabel metal2 s 13104 0 13160 400 0 FreeSans 224 90 0 0 sel[11]
port 17 nsew signal tristate
flabel metal2 s 8736 20600 8792 21000 0 FreeSans 224 90 0 0 sel[1]
port 18 nsew signal tristate
flabel metal3 s 0 12768 400 12824 0 FreeSans 224 0 0 0 sel[2]
port 19 nsew signal tristate
flabel metal3 s 20600 10080 21000 10136 0 FreeSans 224 0 0 0 sel[3]
port 20 nsew signal tristate
flabel metal3 s 20600 11088 21000 11144 0 FreeSans 224 0 0 0 sel[4]
port 21 nsew signal tristate
flabel metal2 s 10752 20600 10808 21000 0 FreeSans 224 90 0 0 sel[5]
port 22 nsew signal tristate
flabel metal3 s 20600 7728 21000 7784 0 FreeSans 224 0 0 0 sel[6]
port 23 nsew signal tristate
flabel metal3 s 20600 9408 21000 9464 0 FreeSans 224 0 0 0 sel[7]
port 24 nsew signal tristate
flabel metal3 s 20600 8736 21000 8792 0 FreeSans 224 0 0 0 sel[8]
port 25 nsew signal tristate
flabel metal2 s 12096 20600 12152 21000 0 FreeSans 224 90 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 2224 1538 2384 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 17584 1538 17744 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 9904 1538 10064 19238 0 FreeSans 640 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 10500 19208 10500 19208 0 vdd
rlabel metal1 10500 18816 10500 18816 0 vss
rlabel metal2 11312 11228 11312 11228 0 _000_
rlabel metal3 8148 7588 8148 7588 0 _001_
rlabel metal3 12768 12796 12768 12796 0 _002_
rlabel metal2 13132 12488 13132 12488 0 _003_
rlabel metal2 9996 13748 9996 13748 0 _004_
rlabel metal2 9548 13300 9548 13300 0 _005_
rlabel metal2 12964 10220 12964 10220 0 _006_
rlabel metal2 13188 7812 13188 7812 0 _007_
rlabel metal2 8260 7000 8260 7000 0 _008_
rlabel metal2 12404 6636 12404 6636 0 _009_
rlabel metal2 10612 6244 10612 6244 0 _010_
rlabel metal2 10808 7756 10808 7756 0 _011_
rlabel metal2 9044 6664 9044 6664 0 _012_
rlabel metal2 11004 12852 11004 12852 0 _013_
rlabel metal2 13244 9296 13244 9296 0 _014_
rlabel metal2 13356 11032 13356 11032 0 _015_
rlabel metal2 13216 8484 13216 8484 0 _016_
rlabel metal2 6580 10668 6580 10668 0 _017_
rlabel metal2 6972 11228 6972 11228 0 _018_
rlabel metal2 6468 8624 6468 8624 0 _019_
rlabel metal3 8848 9212 8848 9212 0 _020_
rlabel metal2 7028 12516 7028 12516 0 _021_
rlabel metal2 8148 12880 8148 12880 0 _022_
rlabel metal2 6524 11732 6524 11732 0 _023_
rlabel metal2 8260 12012 8260 12012 0 _024_
rlabel metal3 9184 12404 9184 12404 0 _025_
rlabel metal2 8316 12600 8316 12600 0 _026_
rlabel metal2 6860 11956 6860 11956 0 _027_
rlabel metal2 12068 10612 12068 10612 0 _028_
rlabel metal2 11452 11620 11452 11620 0 _029_
rlabel metal3 10304 10780 10304 10780 0 _030_
rlabel metal3 12292 11956 12292 11956 0 _031_
rlabel metal2 9716 9996 9716 9996 0 _032_
rlabel metal2 9100 9604 9100 9604 0 _033_
rlabel metal2 9100 7784 9100 7784 0 _034_
rlabel metal2 10444 9800 10444 9800 0 _035_
rlabel metal2 10696 9492 10696 9492 0 _036_
rlabel metal2 9492 11396 9492 11396 0 _037_
rlabel metal2 9408 8428 9408 8428 0 _038_
rlabel metal2 10276 8848 10276 8848 0 _039_
rlabel metal3 9660 7588 9660 7588 0 _040_
rlabel metal3 12824 13468 12824 13468 0 _041_
rlabel metal2 10808 12740 10808 12740 0 _042_
rlabel metal2 10332 12880 10332 12880 0 _043_
rlabel metal2 12964 12432 12964 12432 0 _044_
rlabel metal3 13244 12404 13244 12404 0 _045_
rlabel metal2 9996 13482 9996 13482 0 _046_
rlabel metal2 10220 13468 10220 13468 0 _047_
rlabel metal2 9856 10836 9856 10836 0 _048_
rlabel metal2 9688 13132 9688 13132 0 _049_
rlabel metal3 10052 13468 10052 13468 0 _050_
rlabel metal2 10108 10192 10108 10192 0 _051_
rlabel metal3 13538 9940 13538 9940 0 _052_
rlabel metal3 12628 8036 12628 8036 0 _053_
rlabel metal2 13384 8036 13384 8036 0 _054_
rlabel metal3 10220 8036 10220 8036 0 _055_
rlabel metal2 9156 6944 9156 6944 0 _056_
rlabel metal3 9044 6860 9044 6860 0 _057_
rlabel metal2 11060 8708 11060 8708 0 _058_
rlabel metal2 12824 6916 12824 6916 0 _059_
rlabel metal2 9156 10024 9156 10024 0 _060_
rlabel metal2 9940 7756 9940 7756 0 _061_
rlabel metal2 11284 7112 11284 7112 0 _062_
rlabel metal2 10780 6804 10780 6804 0 _063_
rlabel metal2 10640 8036 10640 8036 0 _064_
rlabel metal2 11900 7840 11900 7840 0 _065_
rlabel metal3 9912 6860 9912 6860 0 _066_
rlabel metal3 9884 7924 9884 7924 0 _067_
rlabel metal2 11284 12600 11284 12600 0 _068_
rlabel metal2 8428 9520 8428 9520 0 _069_
rlabel metal2 11676 9576 11676 9576 0 _070_
rlabel metal2 13748 8372 13748 8372 0 _071_
rlabel metal3 13356 9548 13356 9548 0 _072_
rlabel metal3 7224 10388 7224 10388 0 _073_
rlabel metal2 7420 10528 7420 10528 0 _074_
rlabel metal2 7756 10696 7756 10696 0 _075_
rlabel metal2 9044 8624 9044 8624 0 _076_
rlabel metal3 9156 8708 9156 8708 0 _077_
rlabel metal2 10108 12824 10108 12824 0 _078_
rlabel metal3 12516 9604 12516 9604 0 _079_
rlabel metal2 8764 9016 8764 9016 0 _080_
rlabel metal3 9380 8764 9380 8764 0 _081_
rlabel metal3 9632 9268 9632 9268 0 _082_
rlabel metal2 10388 9240 10388 9240 0 _083_
rlabel metal2 10836 11424 10836 11424 0 _084_
rlabel metal2 10668 12348 10668 12348 0 _085_
rlabel metal2 13496 10836 13496 10836 0 _086_
rlabel metal2 7252 10444 7252 10444 0 _087_
rlabel metal2 8036 10920 8036 10920 0 _088_
rlabel metal2 13328 10780 13328 10780 0 _089_
rlabel metal2 13720 11620 13720 11620 0 _090_
rlabel metal2 13580 11172 13580 11172 0 _091_
rlabel metal2 13524 8568 13524 8568 0 _092_
rlabel metal2 13468 8820 13468 8820 0 _093_
rlabel metal2 10220 10164 10220 10164 0 _094_
rlabel metal2 8316 10304 8316 10304 0 _095_
rlabel metal2 7476 10836 7476 10836 0 _096_
rlabel metal2 8148 9828 8148 9828 0 _097_
rlabel metal2 8820 11536 8820 11536 0 _098_
rlabel metal2 9492 10668 9492 10668 0 _099_
rlabel metal2 11620 10584 11620 10584 0 _100_
rlabel metal3 11088 11844 11088 11844 0 _101_
rlabel metal2 6972 12348 6972 12348 0 _102_
rlabel metal3 7924 9996 7924 9996 0 _103_
rlabel metal2 7364 11340 7364 11340 0 _104_
rlabel metal2 11228 10808 11228 10808 0 _105_
rlabel metal2 10108 9688 10108 9688 0 _106_
rlabel metal2 7308 11872 7308 11872 0 _107_
rlabel metal2 7868 12096 7868 12096 0 _108_
rlabel metal2 7644 11732 7644 11732 0 _109_
rlabel metal2 7392 11676 7392 11676 0 _110_
rlabel metal3 10696 13132 10696 13132 0 _111_
rlabel metal3 1239 13804 1239 13804 0 clk
rlabel metal3 9856 10052 9856 10052 0 clknet_0_clk
rlabel metal2 6076 8820 6076 8820 0 clknet_1_0__leaf_clk
rlabel metal2 10388 13720 10388 13720 0 clknet_1_1__leaf_clk
rlabel metal3 6664 10444 6664 10444 0 dut25.count\[0\]
rlabel metal2 7308 11200 7308 11200 0 dut25.count\[1\]
rlabel metal2 7532 8428 7532 8428 0 dut25.count\[2\]
rlabel metal2 7532 8736 7532 8736 0 dut25.count\[3\]
rlabel metal2 11956 7630 11956 7630 0 net1
rlabel metal3 15190 13188 15190 13188 0 net10
rlabel metal2 14252 13384 14252 13384 0 net11
rlabel metal2 5460 12124 5460 12124 0 net12
rlabel metal2 9100 4312 9100 4312 0 net13
rlabel metal3 13888 6524 13888 6524 0 net14
rlabel metal2 8400 13636 8400 13636 0 net15
rlabel metal2 5964 12712 5964 12712 0 net16
rlabel metal3 18844 10332 18844 10332 0 net17
rlabel metal2 14308 11200 14308 11200 0 net18
rlabel metal3 10864 13972 10864 13972 0 net19
rlabel metal2 8652 8036 8652 8036 0 net2
rlabel metal2 13580 7756 13580 7756 0 net20
rlabel metal2 14308 9380 14308 9380 0 net21
rlabel metal2 14308 8596 14308 8596 0 net22
rlabel metal2 12180 15960 12180 15960 0 net23
rlabel metal2 20132 17248 20132 17248 0 net24
rlabel metal3 10836 18956 10836 18956 0 net25
rlabel metal2 3388 1015 3388 1015 0 net26
rlabel metal2 10136 6524 10136 6524 0 net3
rlabel metal2 14140 12768 14140 12768 0 net4
rlabel metal3 11004 14028 11004 14028 0 net5
rlabel metal2 14644 10360 14644 10360 0 net6
rlabel metal2 10724 13524 10724 13524 0 net7
rlabel metal2 11676 5964 11676 5964 0 net8
rlabel metal2 18844 11424 18844 11424 0 net9
rlabel metal3 12628 2044 12628 2044 0 segm[10]
rlabel metal3 9072 2044 9072 2044 0 segm[11]
rlabel metal3 10500 1708 10500 1708 0 segm[12]
rlabel metal2 20020 12628 20020 12628 0 segm[13]
rlabel metal2 10444 19677 10444 19677 0 segm[2]
rlabel metal2 19964 10584 19964 10584 0 segm[3]
rlabel metal2 9772 19873 9772 19873 0 segm[5]
rlabel metal3 12124 1820 12124 1820 0 segm[6]
rlabel metal3 20321 11452 20321 11452 0 segm[7]
rlabel metal2 19964 13244 19964 13244 0 segm[8]
rlabel metal2 20020 13356 20020 13356 0 segm[9]
rlabel metal3 707 12460 707 12460 0 sel[0]
rlabel metal2 9100 1029 9100 1029 0 sel[10]
rlabel metal2 13132 1029 13132 1029 0 sel[11]
rlabel metal2 8764 19677 8764 19677 0 sel[1]
rlabel metal3 679 12796 679 12796 0 sel[2]
rlabel metal2 20020 10276 20020 10276 0 sel[3]
rlabel metal2 20020 11172 20020 11172 0 sel[4]
rlabel metal2 10780 19873 10780 19873 0 sel[5]
rlabel metal2 20020 7924 20020 7924 0 sel[6]
rlabel metal2 20020 9548 20020 9548 0 sel[7]
rlabel metal2 20020 8820 20020 8820 0 sel[8]
rlabel metal2 12124 19873 12124 19873 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 21000 21000
<< end >>
