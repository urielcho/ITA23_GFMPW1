magic
tech gf180mcuD
magscale 1 10
timestamp 1699641393
<< metal1 >>
rect 1344 38442 40656 38476
rect 1344 38390 4478 38442
rect 4530 38390 4582 38442
rect 4634 38390 4686 38442
rect 4738 38390 35198 38442
rect 35250 38390 35302 38442
rect 35354 38390 35406 38442
rect 35458 38390 40656 38442
rect 1344 38356 40656 38390
rect 14814 38274 14866 38286
rect 14814 38210 14866 38222
rect 18622 38274 18674 38286
rect 18622 38210 18674 38222
rect 25566 38274 25618 38286
rect 25566 38210 25618 38222
rect 21858 38110 21870 38162
rect 21922 38110 21934 38162
rect 14242 37998 14254 38050
rect 14306 37998 14318 38050
rect 17602 37998 17614 38050
rect 17666 37998 17678 38050
rect 20738 37998 20750 38050
rect 20802 37998 20814 38050
rect 24546 37998 24558 38050
rect 24610 37998 24622 38050
rect 1344 37658 40656 37692
rect 1344 37606 19838 37658
rect 19890 37606 19942 37658
rect 19994 37606 20046 37658
rect 20098 37606 40656 37658
rect 1344 37572 40656 37606
rect 15262 37490 15314 37502
rect 15262 37426 15314 37438
rect 22430 37490 22482 37502
rect 22430 37426 22482 37438
rect 26238 37490 26290 37502
rect 26238 37426 26290 37438
rect 14242 37214 14254 37266
rect 14306 37214 14318 37266
rect 25554 37214 25566 37266
rect 25618 37214 25630 37266
rect 1344 36874 40656 36908
rect 1344 36822 4478 36874
rect 4530 36822 4582 36874
rect 4634 36822 4686 36874
rect 4738 36822 35198 36874
rect 35250 36822 35302 36874
rect 35354 36822 35406 36874
rect 35458 36822 40656 36874
rect 1344 36788 40656 36822
rect 1344 36090 40656 36124
rect 1344 36038 19838 36090
rect 19890 36038 19942 36090
rect 19994 36038 20046 36090
rect 20098 36038 40656 36090
rect 1344 36004 40656 36038
rect 1344 35306 40656 35340
rect 1344 35254 4478 35306
rect 4530 35254 4582 35306
rect 4634 35254 4686 35306
rect 4738 35254 35198 35306
rect 35250 35254 35302 35306
rect 35354 35254 35406 35306
rect 35458 35254 40656 35306
rect 1344 35220 40656 35254
rect 1344 34522 40656 34556
rect 1344 34470 19838 34522
rect 19890 34470 19942 34522
rect 19994 34470 20046 34522
rect 20098 34470 40656 34522
rect 1344 34436 40656 34470
rect 1344 33738 40656 33772
rect 1344 33686 4478 33738
rect 4530 33686 4582 33738
rect 4634 33686 4686 33738
rect 4738 33686 35198 33738
rect 35250 33686 35302 33738
rect 35354 33686 35406 33738
rect 35458 33686 40656 33738
rect 1344 33652 40656 33686
rect 1344 32954 40656 32988
rect 1344 32902 19838 32954
rect 19890 32902 19942 32954
rect 19994 32902 20046 32954
rect 20098 32902 40656 32954
rect 1344 32868 40656 32902
rect 1344 32170 40656 32204
rect 1344 32118 4478 32170
rect 4530 32118 4582 32170
rect 4634 32118 4686 32170
rect 4738 32118 35198 32170
rect 35250 32118 35302 32170
rect 35354 32118 35406 32170
rect 35458 32118 40656 32170
rect 1344 32084 40656 32118
rect 1344 31386 40656 31420
rect 1344 31334 19838 31386
rect 19890 31334 19942 31386
rect 19994 31334 20046 31386
rect 20098 31334 40656 31386
rect 1344 31300 40656 31334
rect 1344 30602 40656 30636
rect 1344 30550 4478 30602
rect 4530 30550 4582 30602
rect 4634 30550 4686 30602
rect 4738 30550 35198 30602
rect 35250 30550 35302 30602
rect 35354 30550 35406 30602
rect 35458 30550 40656 30602
rect 1344 30516 40656 30550
rect 1344 29818 40656 29852
rect 1344 29766 19838 29818
rect 19890 29766 19942 29818
rect 19994 29766 20046 29818
rect 20098 29766 40656 29818
rect 1344 29732 40656 29766
rect 1344 29034 40656 29068
rect 1344 28982 4478 29034
rect 4530 28982 4582 29034
rect 4634 28982 4686 29034
rect 4738 28982 35198 29034
rect 35250 28982 35302 29034
rect 35354 28982 35406 29034
rect 35458 28982 40656 29034
rect 1344 28948 40656 28982
rect 19506 28702 19518 28754
rect 19570 28702 19582 28754
rect 19966 28642 20018 28654
rect 16706 28590 16718 28642
rect 16770 28590 16782 28642
rect 19966 28578 20018 28590
rect 17378 28478 17390 28530
rect 17442 28478 17454 28530
rect 13806 28418 13858 28430
rect 13806 28354 13858 28366
rect 1344 28250 40656 28284
rect 1344 28198 19838 28250
rect 19890 28198 19942 28250
rect 19994 28198 20046 28250
rect 20098 28198 40656 28250
rect 1344 28164 40656 28198
rect 17502 28082 17554 28094
rect 17502 28018 17554 28030
rect 17950 27970 18002 27982
rect 17950 27906 18002 27918
rect 18286 27858 18338 27870
rect 23550 27858 23602 27870
rect 10770 27806 10782 27858
rect 10834 27806 10846 27858
rect 14018 27806 14030 27858
rect 14082 27806 14094 27858
rect 20178 27806 20190 27858
rect 20242 27806 20254 27858
rect 18286 27794 18338 27806
rect 23550 27794 23602 27806
rect 11442 27694 11454 27746
rect 11506 27694 11518 27746
rect 13570 27694 13582 27746
rect 13634 27694 13646 27746
rect 14690 27694 14702 27746
rect 14754 27694 14766 27746
rect 16818 27694 16830 27746
rect 16882 27694 16894 27746
rect 20850 27694 20862 27746
rect 20914 27694 20926 27746
rect 22978 27694 22990 27746
rect 23042 27694 23054 27746
rect 1344 27466 40656 27500
rect 1344 27414 4478 27466
rect 4530 27414 4582 27466
rect 4634 27414 4686 27466
rect 4738 27414 35198 27466
rect 35250 27414 35302 27466
rect 35354 27414 35406 27466
rect 35458 27414 40656 27466
rect 1344 27380 40656 27414
rect 15150 27298 15202 27310
rect 15150 27234 15202 27246
rect 15934 27298 15986 27310
rect 15934 27234 15986 27246
rect 1934 27186 1986 27198
rect 1934 27122 1986 27134
rect 16046 27186 16098 27198
rect 21422 27186 21474 27198
rect 26014 27186 26066 27198
rect 16930 27134 16942 27186
rect 16994 27134 17006 27186
rect 25554 27134 25566 27186
rect 25618 27134 25630 27186
rect 16046 27122 16098 27134
rect 21422 27122 21474 27134
rect 26014 27122 26066 27134
rect 40014 27186 40066 27198
rect 40014 27122 40066 27134
rect 14702 27074 14754 27086
rect 4274 27022 4286 27074
rect 4338 27022 4350 27074
rect 14702 27010 14754 27022
rect 15038 27074 15090 27086
rect 16706 27022 16718 27074
rect 16770 27022 16782 27074
rect 22642 27022 22654 27074
rect 22706 27022 22718 27074
rect 37650 27022 37662 27074
rect 37714 27022 37726 27074
rect 15038 27010 15090 27022
rect 13806 26962 13858 26974
rect 13806 26898 13858 26910
rect 13918 26962 13970 26974
rect 13918 26898 13970 26910
rect 14142 26962 14194 26974
rect 16942 26962 16994 26974
rect 14354 26910 14366 26962
rect 14418 26910 14430 26962
rect 14142 26898 14194 26910
rect 16942 26898 16994 26910
rect 17166 26962 17218 26974
rect 17166 26898 17218 26910
rect 17390 26962 17442 26974
rect 17390 26898 17442 26910
rect 18958 26962 19010 26974
rect 18958 26898 19010 26910
rect 19294 26962 19346 26974
rect 19294 26898 19346 26910
rect 21310 26962 21362 26974
rect 21310 26898 21362 26910
rect 21758 26962 21810 26974
rect 27134 26962 27186 26974
rect 23426 26910 23438 26962
rect 23490 26910 23502 26962
rect 21758 26898 21810 26910
rect 27134 26898 27186 26910
rect 27582 26962 27634 26974
rect 27582 26898 27634 26910
rect 27694 26962 27746 26974
rect 27694 26898 27746 26910
rect 15150 26850 15202 26862
rect 15150 26786 15202 26798
rect 21534 26850 21586 26862
rect 21534 26786 21586 26798
rect 26798 26850 26850 26862
rect 26798 26786 26850 26798
rect 27022 26850 27074 26862
rect 27022 26786 27074 26798
rect 27358 26850 27410 26862
rect 27358 26786 27410 26798
rect 1344 26682 40656 26716
rect 1344 26630 19838 26682
rect 19890 26630 19942 26682
rect 19994 26630 20046 26682
rect 20098 26630 40656 26682
rect 1344 26596 40656 26630
rect 20750 26514 20802 26526
rect 20750 26450 20802 26462
rect 23774 26514 23826 26526
rect 23774 26450 23826 26462
rect 14814 26402 14866 26414
rect 14814 26338 14866 26350
rect 14926 26402 14978 26414
rect 14926 26338 14978 26350
rect 18622 26402 18674 26414
rect 18622 26338 18674 26350
rect 19742 26402 19794 26414
rect 19742 26338 19794 26350
rect 19854 26402 19906 26414
rect 19854 26338 19906 26350
rect 20078 26402 20130 26414
rect 20078 26338 20130 26350
rect 21982 26402 22034 26414
rect 21982 26338 22034 26350
rect 22878 26402 22930 26414
rect 22878 26338 22930 26350
rect 14590 26290 14642 26302
rect 14242 26238 14254 26290
rect 14306 26238 14318 26290
rect 14590 26226 14642 26238
rect 18958 26290 19010 26302
rect 18958 26226 19010 26238
rect 20190 26290 20242 26302
rect 20190 26226 20242 26238
rect 20638 26290 20690 26302
rect 20638 26226 20690 26238
rect 20974 26290 21026 26302
rect 20974 26226 21026 26238
rect 21198 26290 21250 26302
rect 21198 26226 21250 26238
rect 21422 26290 21474 26302
rect 22766 26290 22818 26302
rect 21746 26238 21758 26290
rect 21810 26238 21822 26290
rect 21422 26226 21474 26238
rect 22766 26226 22818 26238
rect 23102 26290 23154 26302
rect 23102 26226 23154 26238
rect 23214 26290 23266 26302
rect 23538 26238 23550 26290
rect 23602 26238 23614 26290
rect 25554 26238 25566 26290
rect 25618 26238 25630 26290
rect 37650 26238 37662 26290
rect 37714 26238 37726 26290
rect 23214 26226 23266 26238
rect 15374 26178 15426 26190
rect 11442 26126 11454 26178
rect 11506 26126 11518 26178
rect 13570 26126 13582 26178
rect 13634 26126 13646 26178
rect 15374 26114 15426 26126
rect 18174 26178 18226 26190
rect 18174 26114 18226 26126
rect 18734 26178 18786 26190
rect 28814 26178 28866 26190
rect 26226 26126 26238 26178
rect 26290 26126 26302 26178
rect 28354 26126 28366 26178
rect 28418 26126 28430 26178
rect 18734 26114 18786 26126
rect 28814 26114 28866 26126
rect 18286 26066 18338 26078
rect 18286 26002 18338 26014
rect 19182 26066 19234 26078
rect 19182 26002 19234 26014
rect 19294 26066 19346 26078
rect 19294 26002 19346 26014
rect 20750 26066 20802 26078
rect 20750 26002 20802 26014
rect 22094 26066 22146 26078
rect 22094 26002 22146 26014
rect 23438 26066 23490 26078
rect 23438 26002 23490 26014
rect 40014 26066 40066 26078
rect 40014 26002 40066 26014
rect 1344 25898 40656 25932
rect 1344 25846 4478 25898
rect 4530 25846 4582 25898
rect 4634 25846 4686 25898
rect 4738 25846 35198 25898
rect 35250 25846 35302 25898
rect 35354 25846 35406 25898
rect 35458 25846 40656 25898
rect 1344 25812 40656 25846
rect 21758 25730 21810 25742
rect 21758 25666 21810 25678
rect 13694 25618 13746 25630
rect 21534 25618 21586 25630
rect 29262 25618 29314 25630
rect 18834 25566 18846 25618
rect 18898 25566 18910 25618
rect 19282 25566 19294 25618
rect 19346 25566 19358 25618
rect 26450 25566 26462 25618
rect 26514 25566 26526 25618
rect 28578 25566 28590 25618
rect 28642 25566 28654 25618
rect 13694 25554 13746 25566
rect 21534 25554 21586 25566
rect 29262 25554 29314 25566
rect 13806 25506 13858 25518
rect 13806 25442 13858 25454
rect 14254 25506 14306 25518
rect 19630 25506 19682 25518
rect 19170 25454 19182 25506
rect 19234 25454 19246 25506
rect 14254 25442 14306 25454
rect 19630 25442 19682 25454
rect 22318 25506 22370 25518
rect 25666 25454 25678 25506
rect 25730 25454 25742 25506
rect 22318 25442 22370 25454
rect 13582 25394 13634 25406
rect 13582 25330 13634 25342
rect 17950 25394 18002 25406
rect 17950 25330 18002 25342
rect 18286 25394 18338 25406
rect 18286 25330 18338 25342
rect 18510 25394 18562 25406
rect 18510 25330 18562 25342
rect 19854 25394 19906 25406
rect 19854 25330 19906 25342
rect 21310 25394 21362 25406
rect 21970 25342 21982 25394
rect 22034 25342 22046 25394
rect 21310 25330 21362 25342
rect 18062 25282 18114 25294
rect 18062 25218 18114 25230
rect 18734 25282 18786 25294
rect 18734 25218 18786 25230
rect 19406 25282 19458 25294
rect 19406 25218 19458 25230
rect 20414 25282 20466 25294
rect 20738 25230 20750 25282
rect 20802 25230 20814 25282
rect 21858 25230 21870 25282
rect 21922 25230 21934 25282
rect 20414 25218 20466 25230
rect 1344 25114 40656 25148
rect 1344 25062 19838 25114
rect 19890 25062 19942 25114
rect 19994 25062 20046 25114
rect 20098 25062 40656 25114
rect 1344 25028 40656 25062
rect 26014 24946 26066 24958
rect 17378 24894 17390 24946
rect 17442 24894 17454 24946
rect 19394 24894 19406 24946
rect 19458 24894 19470 24946
rect 26014 24882 26066 24894
rect 26238 24946 26290 24958
rect 26238 24882 26290 24894
rect 27582 24946 27634 24958
rect 27582 24882 27634 24894
rect 27806 24946 27858 24958
rect 27806 24882 27858 24894
rect 18286 24834 18338 24846
rect 26350 24834 26402 24846
rect 20626 24782 20638 24834
rect 20690 24782 20702 24834
rect 18286 24770 18338 24782
rect 26350 24770 26402 24782
rect 18398 24722 18450 24734
rect 17602 24670 17614 24722
rect 17666 24670 17678 24722
rect 18398 24658 18450 24670
rect 19070 24722 19122 24734
rect 27918 24722 27970 24734
rect 20402 24670 20414 24722
rect 20466 24670 20478 24722
rect 19070 24658 19122 24670
rect 27918 24658 27970 24670
rect 18286 24498 18338 24510
rect 18286 24434 18338 24446
rect 1344 24330 40656 24364
rect 1344 24278 4478 24330
rect 4530 24278 4582 24330
rect 4634 24278 4686 24330
rect 4738 24278 35198 24330
rect 35250 24278 35302 24330
rect 35354 24278 35406 24330
rect 35458 24278 40656 24330
rect 1344 24244 40656 24278
rect 13694 24162 13746 24174
rect 13694 24098 13746 24110
rect 1934 24050 1986 24062
rect 1934 23986 1986 23998
rect 40014 24050 40066 24062
rect 40014 23986 40066 23998
rect 4274 23886 4286 23938
rect 4338 23886 4350 23938
rect 37650 23886 37662 23938
rect 37714 23886 37726 23938
rect 13694 23826 13746 23838
rect 13694 23762 13746 23774
rect 13806 23826 13858 23838
rect 13806 23762 13858 23774
rect 14254 23826 14306 23838
rect 14254 23762 14306 23774
rect 14366 23826 14418 23838
rect 14366 23762 14418 23774
rect 18174 23826 18226 23838
rect 18174 23762 18226 23774
rect 18510 23826 18562 23838
rect 18510 23762 18562 23774
rect 14030 23714 14082 23726
rect 14030 23650 14082 23662
rect 16606 23714 16658 23726
rect 16606 23650 16658 23662
rect 18398 23714 18450 23726
rect 18398 23650 18450 23662
rect 26126 23714 26178 23726
rect 37326 23714 37378 23726
rect 26450 23662 26462 23714
rect 26514 23662 26526 23714
rect 26126 23650 26178 23662
rect 37326 23650 37378 23662
rect 1344 23546 40656 23580
rect 1344 23494 19838 23546
rect 19890 23494 19942 23546
rect 19994 23494 20046 23546
rect 20098 23494 40656 23546
rect 1344 23460 40656 23494
rect 14366 23378 14418 23390
rect 14366 23314 14418 23326
rect 17614 23378 17666 23390
rect 19854 23378 19906 23390
rect 18498 23326 18510 23378
rect 18562 23326 18574 23378
rect 17614 23314 17666 23326
rect 19854 23314 19906 23326
rect 17726 23266 17778 23278
rect 19630 23266 19682 23278
rect 13122 23214 13134 23266
rect 13186 23214 13198 23266
rect 15586 23214 15598 23266
rect 15650 23214 15662 23266
rect 18834 23214 18846 23266
rect 18898 23214 18910 23266
rect 17726 23202 17778 23214
rect 19630 23202 19682 23214
rect 21198 23266 21250 23278
rect 21198 23202 21250 23214
rect 16046 23154 16098 23166
rect 19518 23154 19570 23166
rect 13906 23102 13918 23154
rect 13970 23102 13982 23154
rect 15362 23102 15374 23154
rect 15426 23102 15438 23154
rect 18274 23102 18286 23154
rect 18338 23102 18350 23154
rect 19058 23102 19070 23154
rect 19122 23102 19134 23154
rect 16046 23090 16098 23102
rect 19518 23090 19570 23102
rect 20190 23154 20242 23166
rect 20190 23090 20242 23102
rect 20526 23154 20578 23166
rect 20526 23090 20578 23102
rect 20638 23154 20690 23166
rect 21858 23102 21870 23154
rect 21922 23102 21934 23154
rect 37874 23102 37886 23154
rect 37938 23102 37950 23154
rect 20638 23090 20690 23102
rect 16718 23042 16770 23054
rect 10994 22990 11006 23042
rect 11058 22990 11070 23042
rect 16718 22978 16770 22990
rect 16830 23042 16882 23054
rect 16830 22978 16882 22990
rect 17502 23042 17554 23054
rect 17502 22978 17554 22990
rect 20302 23042 20354 23054
rect 25342 23042 25394 23054
rect 21074 22990 21086 23042
rect 21138 22990 21150 23042
rect 22530 22990 22542 23042
rect 22594 22990 22606 23042
rect 24658 22990 24670 23042
rect 24722 22990 24734 23042
rect 20302 22978 20354 22990
rect 25342 22978 25394 22990
rect 15934 22930 15986 22942
rect 15934 22866 15986 22878
rect 21422 22930 21474 22942
rect 21422 22866 21474 22878
rect 40014 22930 40066 22942
rect 40014 22866 40066 22878
rect 1344 22762 40656 22796
rect 1344 22710 4478 22762
rect 4530 22710 4582 22762
rect 4634 22710 4686 22762
rect 4738 22710 35198 22762
rect 35250 22710 35302 22762
rect 35354 22710 35406 22762
rect 35458 22710 40656 22762
rect 1344 22676 40656 22710
rect 17278 22594 17330 22606
rect 17278 22530 17330 22542
rect 17950 22594 18002 22606
rect 17950 22530 18002 22542
rect 18846 22594 18898 22606
rect 28254 22594 28306 22606
rect 20514 22542 20526 22594
rect 20578 22591 20590 22594
rect 20850 22591 20862 22594
rect 20578 22545 20862 22591
rect 20578 22542 20590 22545
rect 20850 22542 20862 22545
rect 20914 22542 20926 22594
rect 18846 22530 18898 22542
rect 28254 22530 28306 22542
rect 40014 22482 40066 22494
rect 16370 22430 16382 22482
rect 16434 22430 16446 22482
rect 22754 22430 22766 22482
rect 22818 22430 22830 22482
rect 26786 22430 26798 22482
rect 26850 22430 26862 22482
rect 40014 22418 40066 22430
rect 16942 22370 16994 22382
rect 20750 22370 20802 22382
rect 22318 22370 22370 22382
rect 27806 22370 27858 22382
rect 13570 22318 13582 22370
rect 13634 22318 13646 22370
rect 18386 22318 18398 22370
rect 18450 22318 18462 22370
rect 19618 22318 19630 22370
rect 19682 22318 19694 22370
rect 21522 22318 21534 22370
rect 21586 22318 21598 22370
rect 22530 22318 22542 22370
rect 22594 22318 22606 22370
rect 23986 22318 23998 22370
rect 24050 22318 24062 22370
rect 29362 22318 29374 22370
rect 29426 22318 29438 22370
rect 37650 22318 37662 22370
rect 37714 22318 37726 22370
rect 16942 22306 16994 22318
rect 20750 22306 20802 22318
rect 22318 22306 22370 22318
rect 27806 22306 27858 22318
rect 17614 22258 17666 22270
rect 14242 22206 14254 22258
rect 14306 22206 14318 22258
rect 17614 22194 17666 22206
rect 17838 22258 17890 22270
rect 21310 22258 21362 22270
rect 28142 22258 28194 22270
rect 18946 22206 18958 22258
rect 19010 22206 19022 22258
rect 19730 22206 19742 22258
rect 19794 22206 19806 22258
rect 24658 22206 24670 22258
rect 24722 22206 24734 22258
rect 17838 22194 17890 22206
rect 21310 22194 21362 22206
rect 28142 22194 28194 22206
rect 17166 22146 17218 22158
rect 27246 22146 27298 22158
rect 20178 22094 20190 22146
rect 20242 22094 20254 22146
rect 17166 22082 17218 22094
rect 27246 22082 27298 22094
rect 27470 22146 27522 22158
rect 27470 22082 27522 22094
rect 27694 22146 27746 22158
rect 27694 22082 27746 22094
rect 28254 22146 28306 22158
rect 29586 22094 29598 22146
rect 29650 22094 29662 22146
rect 28254 22082 28306 22094
rect 1344 21978 40656 22012
rect 1344 21926 19838 21978
rect 19890 21926 19942 21978
rect 19994 21926 20046 21978
rect 20098 21926 40656 21978
rect 1344 21892 40656 21926
rect 14590 21810 14642 21822
rect 25454 21810 25506 21822
rect 15250 21758 15262 21810
rect 15314 21758 15326 21810
rect 15922 21758 15934 21810
rect 15986 21758 15998 21810
rect 18386 21758 18398 21810
rect 18450 21758 18462 21810
rect 14590 21746 14642 21758
rect 25454 21746 25506 21758
rect 14926 21698 14978 21710
rect 25342 21698 25394 21710
rect 17938 21646 17950 21698
rect 18002 21646 18014 21698
rect 18162 21646 18174 21698
rect 18226 21646 18238 21698
rect 14926 21634 14978 21646
rect 25342 21634 25394 21646
rect 25566 21698 25618 21710
rect 27794 21646 27806 21698
rect 27858 21646 27870 21698
rect 25566 21634 25618 21646
rect 16830 21586 16882 21598
rect 11330 21534 11342 21586
rect 11394 21534 11406 21586
rect 12002 21534 12014 21586
rect 12066 21534 12078 21586
rect 15698 21534 15710 21586
rect 15762 21534 15774 21586
rect 16370 21534 16382 21586
rect 16434 21534 16446 21586
rect 16830 21522 16882 21534
rect 18622 21586 18674 21598
rect 25230 21586 25282 21598
rect 19058 21534 19070 21586
rect 19122 21534 19134 21586
rect 26002 21534 26014 21586
rect 26066 21534 26078 21586
rect 27010 21534 27022 21586
rect 27074 21534 27086 21586
rect 37650 21534 37662 21586
rect 37714 21534 37726 21586
rect 18622 21522 18674 21534
rect 25230 21522 25282 21534
rect 26686 21474 26738 21486
rect 40014 21474 40066 21486
rect 14130 21422 14142 21474
rect 14194 21422 14206 21474
rect 22866 21422 22878 21474
rect 22930 21422 22942 21474
rect 29922 21422 29934 21474
rect 29986 21422 29998 21474
rect 26686 21410 26738 21422
rect 40014 21410 40066 21422
rect 1344 21194 40656 21228
rect 1344 21142 4478 21194
rect 4530 21142 4582 21194
rect 4634 21142 4686 21194
rect 4738 21142 35198 21194
rect 35250 21142 35302 21194
rect 35354 21142 35406 21194
rect 35458 21142 40656 21194
rect 1344 21108 40656 21142
rect 22530 20862 22542 20914
rect 22594 20862 22606 20914
rect 27010 20862 27022 20914
rect 27074 20862 27086 20914
rect 14366 20802 14418 20814
rect 21758 20802 21810 20814
rect 20066 20750 20078 20802
rect 20130 20750 20142 20802
rect 22866 20750 22878 20802
rect 22930 20750 22942 20802
rect 14366 20738 14418 20750
rect 21758 20738 21810 20750
rect 14590 20690 14642 20702
rect 14590 20626 14642 20638
rect 14702 20690 14754 20702
rect 21982 20690 22034 20702
rect 15698 20638 15710 20690
rect 15762 20638 15774 20690
rect 14702 20626 14754 20638
rect 21982 20626 22034 20638
rect 22094 20690 22146 20702
rect 22306 20638 22318 20690
rect 22370 20638 22382 20690
rect 22094 20626 22146 20638
rect 21534 20578 21586 20590
rect 21534 20514 21586 20526
rect 1344 20410 40656 20444
rect 1344 20358 19838 20410
rect 19890 20358 19942 20410
rect 19994 20358 20046 20410
rect 20098 20358 40656 20410
rect 1344 20324 40656 20358
rect 18174 20242 18226 20254
rect 18174 20178 18226 20190
rect 18622 20242 18674 20254
rect 18622 20178 18674 20190
rect 18846 20242 18898 20254
rect 18846 20178 18898 20190
rect 20190 20242 20242 20254
rect 22542 20242 22594 20254
rect 21410 20190 21422 20242
rect 21474 20190 21486 20242
rect 20190 20178 20242 20190
rect 22542 20178 22594 20190
rect 25902 20242 25954 20254
rect 25902 20178 25954 20190
rect 26014 20242 26066 20254
rect 26014 20178 26066 20190
rect 19854 20130 19906 20142
rect 19854 20066 19906 20078
rect 19966 20130 20018 20142
rect 19966 20066 20018 20078
rect 20750 20130 20802 20142
rect 20750 20066 20802 20078
rect 21758 20130 21810 20142
rect 21758 20066 21810 20078
rect 22654 20130 22706 20142
rect 22654 20066 22706 20078
rect 22766 20130 22818 20142
rect 23662 20130 23714 20142
rect 22978 20078 22990 20130
rect 23042 20078 23054 20130
rect 22766 20066 22818 20078
rect 23662 20066 23714 20078
rect 18734 20018 18786 20030
rect 18050 19966 18062 20018
rect 18114 19966 18126 20018
rect 18734 19954 18786 19966
rect 19294 20018 19346 20030
rect 22430 20018 22482 20030
rect 20962 19966 20974 20018
rect 21026 19966 21038 20018
rect 19294 19954 19346 19966
rect 22430 19954 22482 19966
rect 23438 20018 23490 20030
rect 23438 19954 23490 19966
rect 23774 20018 23826 20030
rect 23774 19954 23826 19966
rect 25342 20018 25394 20030
rect 25666 19966 25678 20018
rect 25730 19966 25742 20018
rect 26338 19966 26350 20018
rect 26402 19966 26414 20018
rect 37650 19966 37662 20018
rect 37714 19966 37726 20018
rect 25342 19954 25394 19966
rect 17726 19906 17778 19918
rect 29598 19906 29650 19918
rect 27010 19854 27022 19906
rect 27074 19854 27086 19906
rect 29138 19854 29150 19906
rect 29202 19854 29214 19906
rect 17726 19842 17778 19854
rect 29598 19842 29650 19854
rect 20638 19794 20690 19806
rect 20638 19730 20690 19742
rect 40014 19794 40066 19806
rect 40014 19730 40066 19742
rect 1344 19626 40656 19660
rect 1344 19574 4478 19626
rect 4530 19574 4582 19626
rect 4634 19574 4686 19626
rect 4738 19574 35198 19626
rect 35250 19574 35302 19626
rect 35354 19574 35406 19626
rect 35458 19574 40656 19626
rect 1344 19540 40656 19574
rect 19406 19458 19458 19470
rect 19406 19394 19458 19406
rect 22206 19458 22258 19470
rect 22206 19394 22258 19406
rect 26798 19458 26850 19470
rect 26798 19394 26850 19406
rect 15262 19346 15314 19358
rect 15262 19282 15314 19294
rect 40014 19346 40066 19358
rect 40014 19282 40066 19294
rect 19742 19234 19794 19246
rect 21310 19234 21362 19246
rect 14690 19182 14702 19234
rect 14754 19182 14766 19234
rect 16930 19182 16942 19234
rect 16994 19182 17006 19234
rect 17490 19182 17502 19234
rect 17554 19182 17566 19234
rect 18386 19182 18398 19234
rect 18450 19182 18462 19234
rect 18722 19182 18734 19234
rect 18786 19182 18798 19234
rect 20514 19182 20526 19234
rect 20578 19182 20590 19234
rect 19742 19170 19794 19182
rect 21310 19170 21362 19182
rect 25342 19234 25394 19246
rect 25666 19182 25678 19234
rect 25730 19182 25742 19234
rect 37874 19182 37886 19234
rect 37938 19182 37950 19234
rect 25342 19170 25394 19182
rect 19294 19122 19346 19134
rect 22430 19122 22482 19134
rect 17154 19070 17166 19122
rect 17218 19070 17230 19122
rect 17602 19070 17614 19122
rect 17666 19070 17678 19122
rect 18946 19070 18958 19122
rect 19010 19070 19022 19122
rect 20066 19070 20078 19122
rect 20130 19070 20142 19122
rect 21634 19070 21646 19122
rect 21698 19070 21710 19122
rect 19294 19058 19346 19070
rect 22430 19058 22482 19070
rect 25118 19122 25170 19134
rect 25118 19058 25170 19070
rect 25902 19122 25954 19134
rect 25902 19058 25954 19070
rect 26014 19122 26066 19134
rect 26014 19058 26066 19070
rect 26238 19122 26290 19134
rect 26238 19058 26290 19070
rect 14478 19010 14530 19022
rect 22318 19010 22370 19022
rect 20738 18958 20750 19010
rect 20802 18958 20814 19010
rect 14478 18946 14530 18958
rect 22318 18946 22370 18958
rect 24894 19010 24946 19022
rect 24894 18946 24946 18958
rect 25006 19010 25058 19022
rect 25006 18946 25058 18958
rect 26462 19010 26514 19022
rect 26462 18946 26514 18958
rect 26686 19010 26738 19022
rect 26686 18946 26738 18958
rect 1344 18842 40656 18876
rect 1344 18790 19838 18842
rect 19890 18790 19942 18842
rect 19994 18790 20046 18842
rect 20098 18790 40656 18842
rect 1344 18756 40656 18790
rect 22990 18674 23042 18686
rect 15922 18622 15934 18674
rect 15986 18622 15998 18674
rect 16818 18622 16830 18674
rect 16882 18622 16894 18674
rect 17826 18622 17838 18674
rect 17890 18622 17902 18674
rect 18162 18622 18174 18674
rect 18226 18622 18238 18674
rect 21634 18622 21646 18674
rect 21698 18622 21710 18674
rect 22990 18610 23042 18622
rect 24110 18674 24162 18686
rect 24110 18610 24162 18622
rect 24558 18674 24610 18686
rect 24558 18610 24610 18622
rect 19070 18562 19122 18574
rect 19070 18498 19122 18510
rect 19182 18562 19234 18574
rect 19182 18498 19234 18510
rect 21982 18562 22034 18574
rect 21982 18498 22034 18510
rect 23886 18562 23938 18574
rect 23886 18498 23938 18510
rect 15374 18450 15426 18462
rect 12226 18398 12238 18450
rect 12290 18398 12302 18450
rect 15374 18386 15426 18398
rect 17502 18450 17554 18462
rect 17502 18386 17554 18398
rect 18510 18450 18562 18462
rect 18510 18386 18562 18398
rect 18734 18450 18786 18462
rect 18734 18386 18786 18398
rect 19406 18450 19458 18462
rect 19406 18386 19458 18398
rect 19854 18450 19906 18462
rect 22542 18450 22594 18462
rect 20178 18398 20190 18450
rect 20242 18398 20254 18450
rect 20738 18398 20750 18450
rect 20802 18398 20814 18450
rect 21186 18398 21198 18450
rect 21250 18398 21262 18450
rect 21746 18398 21758 18450
rect 21810 18398 21822 18450
rect 19854 18386 19906 18398
rect 22542 18386 22594 18398
rect 23214 18450 23266 18462
rect 23214 18386 23266 18398
rect 23550 18450 23602 18462
rect 23550 18386 23602 18398
rect 24446 18450 24498 18462
rect 24446 18386 24498 18398
rect 24782 18450 24834 18462
rect 28590 18450 28642 18462
rect 25330 18398 25342 18450
rect 25394 18398 25406 18450
rect 37650 18398 37662 18450
rect 37714 18398 37726 18450
rect 24782 18386 24834 18398
rect 28590 18386 28642 18398
rect 16270 18338 16322 18350
rect 12898 18286 12910 18338
rect 12962 18286 12974 18338
rect 15026 18286 15038 18338
rect 15090 18286 15102 18338
rect 16270 18274 16322 18286
rect 22766 18338 22818 18350
rect 23090 18286 23102 18338
rect 23154 18286 23166 18338
rect 26002 18286 26014 18338
rect 26066 18286 26078 18338
rect 28130 18286 28142 18338
rect 28194 18286 28206 18338
rect 22766 18274 22818 18286
rect 15598 18226 15650 18238
rect 15598 18162 15650 18174
rect 16494 18226 16546 18238
rect 22318 18226 22370 18238
rect 20178 18174 20190 18226
rect 20242 18174 20254 18226
rect 21410 18174 21422 18226
rect 21474 18174 21486 18226
rect 16494 18162 16546 18174
rect 22318 18162 22370 18174
rect 24222 18226 24274 18238
rect 24222 18162 24274 18174
rect 40014 18226 40066 18238
rect 40014 18162 40066 18174
rect 1344 18058 40656 18092
rect 1344 18006 4478 18058
rect 4530 18006 4582 18058
rect 4634 18006 4686 18058
rect 4738 18006 35198 18058
rect 35250 18006 35302 18058
rect 35354 18006 35406 18058
rect 35458 18006 40656 18058
rect 1344 17972 40656 18006
rect 18622 17890 18674 17902
rect 28018 17838 28030 17890
rect 28082 17838 28094 17890
rect 18622 17826 18674 17838
rect 14254 17778 14306 17790
rect 22754 17726 22766 17778
rect 22818 17726 22830 17778
rect 24882 17726 24894 17778
rect 24946 17726 24958 17778
rect 14254 17714 14306 17726
rect 15150 17666 15202 17678
rect 14914 17614 14926 17666
rect 14978 17614 14990 17666
rect 15150 17602 15202 17614
rect 15598 17666 15650 17678
rect 15598 17602 15650 17614
rect 16718 17666 16770 17678
rect 19294 17666 19346 17678
rect 17602 17614 17614 17666
rect 17666 17614 17678 17666
rect 16718 17602 16770 17614
rect 19294 17602 19346 17614
rect 19406 17666 19458 17678
rect 25454 17666 25506 17678
rect 27022 17666 27074 17678
rect 20066 17614 20078 17666
rect 20130 17614 20142 17666
rect 21970 17614 21982 17666
rect 22034 17614 22046 17666
rect 25778 17614 25790 17666
rect 25842 17614 25854 17666
rect 26562 17614 26574 17666
rect 26626 17614 26638 17666
rect 19406 17602 19458 17614
rect 25454 17602 25506 17614
rect 27022 17602 27074 17614
rect 18510 17554 18562 17566
rect 15922 17502 15934 17554
rect 15986 17502 15998 17554
rect 17042 17502 17054 17554
rect 17106 17502 17118 17554
rect 18510 17490 18562 17502
rect 18958 17554 19010 17566
rect 25230 17554 25282 17566
rect 20290 17502 20302 17554
rect 20354 17502 20366 17554
rect 18958 17490 19010 17502
rect 25230 17490 25282 17502
rect 19070 17442 19122 17454
rect 17378 17390 17390 17442
rect 17442 17390 17454 17442
rect 19070 17378 19122 17390
rect 25342 17442 25394 17454
rect 25342 17378 25394 17390
rect 26798 17442 26850 17454
rect 26798 17378 26850 17390
rect 26910 17442 26962 17454
rect 26910 17378 26962 17390
rect 27134 17442 27186 17454
rect 27906 17390 27918 17442
rect 27970 17439 27982 17442
rect 28033 17439 28079 17838
rect 40014 17778 40066 17790
rect 40014 17714 40066 17726
rect 28366 17666 28418 17678
rect 28366 17602 28418 17614
rect 28478 17666 28530 17678
rect 37650 17614 37662 17666
rect 37714 17614 37726 17666
rect 28478 17602 28530 17614
rect 27970 17393 28079 17439
rect 27970 17390 27982 17393
rect 27134 17378 27186 17390
rect 1344 17274 40656 17308
rect 1344 17222 19838 17274
rect 19890 17222 19942 17274
rect 19994 17222 20046 17274
rect 20098 17222 40656 17274
rect 1344 17188 40656 17222
rect 15486 17106 15538 17118
rect 15486 17042 15538 17054
rect 23998 17106 24050 17118
rect 23998 17042 24050 17054
rect 25342 17106 25394 17118
rect 25342 17042 25394 17054
rect 26238 17106 26290 17118
rect 26238 17042 26290 17054
rect 24110 16994 24162 17006
rect 12898 16942 12910 16994
rect 12962 16942 12974 16994
rect 27346 16942 27358 16994
rect 27410 16942 27422 16994
rect 24110 16930 24162 16942
rect 12226 16830 12238 16882
rect 12290 16830 12302 16882
rect 26562 16830 26574 16882
rect 26626 16830 26638 16882
rect 15026 16718 15038 16770
rect 15090 16718 15102 16770
rect 29474 16718 29486 16770
rect 29538 16718 29550 16770
rect 1344 16490 40656 16524
rect 1344 16438 4478 16490
rect 4530 16438 4582 16490
rect 4634 16438 4686 16490
rect 4738 16438 35198 16490
rect 35250 16438 35302 16490
rect 35354 16438 35406 16490
rect 35458 16438 40656 16490
rect 1344 16404 40656 16438
rect 1344 15706 40656 15740
rect 1344 15654 19838 15706
rect 19890 15654 19942 15706
rect 19994 15654 20046 15706
rect 20098 15654 40656 15706
rect 1344 15620 40656 15654
rect 25678 15538 25730 15550
rect 25678 15474 25730 15486
rect 26126 15538 26178 15550
rect 26126 15474 26178 15486
rect 15486 15426 15538 15438
rect 15486 15362 15538 15374
rect 15710 15426 15762 15438
rect 15710 15362 15762 15374
rect 18174 15426 18226 15438
rect 18174 15362 18226 15374
rect 18734 15426 18786 15438
rect 18734 15362 18786 15374
rect 19294 15426 19346 15438
rect 19294 15362 19346 15374
rect 19630 15426 19682 15438
rect 19630 15362 19682 15374
rect 21870 15426 21922 15438
rect 22194 15374 22206 15426
rect 22258 15374 22270 15426
rect 21870 15362 21922 15374
rect 18846 15314 18898 15326
rect 16482 15262 16494 15314
rect 16546 15262 16558 15314
rect 18846 15250 18898 15262
rect 19070 15314 19122 15326
rect 25902 15314 25954 15326
rect 22418 15262 22430 15314
rect 22482 15262 22494 15314
rect 37650 15262 37662 15314
rect 37714 15262 37726 15314
rect 19070 15250 19122 15262
rect 25902 15250 25954 15262
rect 16158 15202 16210 15214
rect 15810 15150 15822 15202
rect 15874 15150 15886 15202
rect 16158 15138 16210 15150
rect 16270 15202 16322 15214
rect 16270 15138 16322 15150
rect 18398 15202 18450 15214
rect 18398 15138 18450 15150
rect 19854 15202 19906 15214
rect 19854 15138 19906 15150
rect 26014 15202 26066 15214
rect 26014 15138 26066 15150
rect 40014 15202 40066 15214
rect 40014 15138 40066 15150
rect 18062 15090 18114 15102
rect 18062 15026 18114 15038
rect 20190 15090 20242 15102
rect 20190 15026 20242 15038
rect 21758 15090 21810 15102
rect 21758 15026 21810 15038
rect 1344 14922 40656 14956
rect 1344 14870 4478 14922
rect 4530 14870 4582 14922
rect 4634 14870 4686 14922
rect 4738 14870 35198 14922
rect 35250 14870 35302 14922
rect 35354 14870 35406 14922
rect 35458 14870 40656 14922
rect 1344 14836 40656 14870
rect 23326 14642 23378 14654
rect 28254 14642 28306 14654
rect 17042 14590 17054 14642
rect 17106 14590 17118 14642
rect 19170 14590 19182 14642
rect 19234 14590 19246 14642
rect 25666 14590 25678 14642
rect 25730 14590 25742 14642
rect 27794 14590 27806 14642
rect 27858 14590 27870 14642
rect 23326 14578 23378 14590
rect 28254 14578 28306 14590
rect 19630 14530 19682 14542
rect 16258 14478 16270 14530
rect 16322 14478 16334 14530
rect 19630 14466 19682 14478
rect 19854 14530 19906 14542
rect 21870 14530 21922 14542
rect 20178 14478 20190 14530
rect 20242 14478 20254 14530
rect 21298 14478 21310 14530
rect 21362 14478 21374 14530
rect 19854 14466 19906 14478
rect 21870 14466 21922 14478
rect 22206 14530 22258 14542
rect 22206 14466 22258 14478
rect 22654 14530 22706 14542
rect 22654 14466 22706 14478
rect 22878 14530 22930 14542
rect 22878 14466 22930 14478
rect 23662 14530 23714 14542
rect 24994 14478 25006 14530
rect 25058 14478 25070 14530
rect 23662 14466 23714 14478
rect 19966 14418 20018 14430
rect 19966 14354 20018 14366
rect 23214 14418 23266 14430
rect 23214 14354 23266 14366
rect 23550 14418 23602 14430
rect 23550 14354 23602 14366
rect 19742 14306 19794 14318
rect 19742 14242 19794 14254
rect 20638 14306 20690 14318
rect 20638 14242 20690 14254
rect 21534 14306 21586 14318
rect 21534 14242 21586 14254
rect 21646 14306 21698 14318
rect 21646 14242 21698 14254
rect 21758 14306 21810 14318
rect 21758 14242 21810 14254
rect 22542 14306 22594 14318
rect 22542 14242 22594 14254
rect 1344 14138 40656 14172
rect 1344 14086 19838 14138
rect 19890 14086 19942 14138
rect 19994 14086 20046 14138
rect 20098 14086 40656 14138
rect 1344 14052 40656 14086
rect 16830 13970 16882 13982
rect 16830 13906 16882 13918
rect 21534 13970 21586 13982
rect 21534 13906 21586 13918
rect 26910 13970 26962 13982
rect 26910 13906 26962 13918
rect 21310 13858 21362 13870
rect 27022 13858 27074 13870
rect 13906 13806 13918 13858
rect 13970 13806 13982 13858
rect 18274 13806 18286 13858
rect 18338 13806 18350 13858
rect 22530 13806 22542 13858
rect 22594 13806 22606 13858
rect 25554 13806 25566 13858
rect 25618 13806 25630 13858
rect 21310 13794 21362 13806
rect 27022 13794 27074 13806
rect 21198 13746 21250 13758
rect 25230 13746 25282 13758
rect 13234 13694 13246 13746
rect 13298 13694 13310 13746
rect 17602 13694 17614 13746
rect 17666 13694 17678 13746
rect 21858 13694 21870 13746
rect 21922 13694 21934 13746
rect 21198 13682 21250 13694
rect 25230 13682 25282 13694
rect 16034 13582 16046 13634
rect 16098 13582 16110 13634
rect 20402 13582 20414 13634
rect 20466 13582 20478 13634
rect 24658 13582 24670 13634
rect 24722 13582 24734 13634
rect 1344 13354 40656 13388
rect 1344 13302 4478 13354
rect 4530 13302 4582 13354
rect 4634 13302 4686 13354
rect 4738 13302 35198 13354
rect 35250 13302 35302 13354
rect 35354 13302 35406 13354
rect 35458 13302 40656 13354
rect 1344 13268 40656 13302
rect 20526 13186 20578 13198
rect 20526 13122 20578 13134
rect 16382 13074 16434 13086
rect 25006 13074 25058 13086
rect 22082 13022 22094 13074
rect 22146 13022 22158 13074
rect 24210 13022 24222 13074
rect 24274 13022 24286 13074
rect 16382 13010 16434 13022
rect 25006 13010 25058 13022
rect 25454 13074 25506 13086
rect 25454 13010 25506 13022
rect 20638 12962 20690 12974
rect 21410 12910 21422 12962
rect 21474 12910 21486 12962
rect 20638 12898 20690 12910
rect 20526 12738 20578 12750
rect 20526 12674 20578 12686
rect 1344 12570 40656 12604
rect 1344 12518 19838 12570
rect 19890 12518 19942 12570
rect 19994 12518 20046 12570
rect 20098 12518 40656 12570
rect 1344 12484 40656 12518
rect 1344 11786 40656 11820
rect 1344 11734 4478 11786
rect 4530 11734 4582 11786
rect 4634 11734 4686 11786
rect 4738 11734 35198 11786
rect 35250 11734 35302 11786
rect 35354 11734 35406 11786
rect 35458 11734 40656 11786
rect 1344 11700 40656 11734
rect 1344 11002 40656 11036
rect 1344 10950 19838 11002
rect 19890 10950 19942 11002
rect 19994 10950 20046 11002
rect 20098 10950 40656 11002
rect 1344 10916 40656 10950
rect 1344 10218 40656 10252
rect 1344 10166 4478 10218
rect 4530 10166 4582 10218
rect 4634 10166 4686 10218
rect 4738 10166 35198 10218
rect 35250 10166 35302 10218
rect 35354 10166 35406 10218
rect 35458 10166 40656 10218
rect 1344 10132 40656 10166
rect 1344 9434 40656 9468
rect 1344 9382 19838 9434
rect 19890 9382 19942 9434
rect 19994 9382 20046 9434
rect 20098 9382 40656 9434
rect 1344 9348 40656 9382
rect 1344 8650 40656 8684
rect 1344 8598 4478 8650
rect 4530 8598 4582 8650
rect 4634 8598 4686 8650
rect 4738 8598 35198 8650
rect 35250 8598 35302 8650
rect 35354 8598 35406 8650
rect 35458 8598 40656 8650
rect 1344 8564 40656 8598
rect 1344 7866 40656 7900
rect 1344 7814 19838 7866
rect 19890 7814 19942 7866
rect 19994 7814 20046 7866
rect 20098 7814 40656 7866
rect 1344 7780 40656 7814
rect 1344 7082 40656 7116
rect 1344 7030 4478 7082
rect 4530 7030 4582 7082
rect 4634 7030 4686 7082
rect 4738 7030 35198 7082
rect 35250 7030 35302 7082
rect 35354 7030 35406 7082
rect 35458 7030 40656 7082
rect 1344 6996 40656 7030
rect 1344 6298 40656 6332
rect 1344 6246 19838 6298
rect 19890 6246 19942 6298
rect 19994 6246 20046 6298
rect 20098 6246 40656 6298
rect 1344 6212 40656 6246
rect 1344 5514 40656 5548
rect 1344 5462 4478 5514
rect 4530 5462 4582 5514
rect 4634 5462 4686 5514
rect 4738 5462 35198 5514
rect 35250 5462 35302 5514
rect 35354 5462 35406 5514
rect 35458 5462 40656 5514
rect 1344 5428 40656 5462
rect 1344 4730 40656 4764
rect 1344 4678 19838 4730
rect 19890 4678 19942 4730
rect 19994 4678 20046 4730
rect 20098 4678 40656 4730
rect 1344 4644 40656 4678
rect 17378 4286 17390 4338
rect 17442 4286 17454 4338
rect 20402 4286 20414 4338
rect 20466 4286 20478 4338
rect 25330 4286 25342 4338
rect 25394 4286 25406 4338
rect 18498 4174 18510 4226
rect 18562 4174 18574 4226
rect 21422 4114 21474 4126
rect 21422 4050 21474 4062
rect 26238 4114 26290 4126
rect 26238 4050 26290 4062
rect 1344 3946 40656 3980
rect 1344 3894 4478 3946
rect 4530 3894 4582 3946
rect 4634 3894 4686 3946
rect 4738 3894 35198 3946
rect 35250 3894 35302 3946
rect 35354 3894 35406 3946
rect 35458 3894 40656 3946
rect 1344 3860 40656 3894
rect 25566 3666 25618 3678
rect 25566 3602 25618 3614
rect 18050 3502 18062 3554
rect 18114 3502 18126 3554
rect 23538 3502 23550 3554
rect 23602 3502 23614 3554
rect 24546 3502 24558 3554
rect 24610 3502 24622 3554
rect 19394 3390 19406 3442
rect 19458 3390 19470 3442
rect 22194 3390 22206 3442
rect 22258 3390 22270 3442
rect 1344 3162 40656 3196
rect 1344 3110 19838 3162
rect 19890 3110 19942 3162
rect 19994 3110 20046 3162
rect 20098 3110 40656 3162
rect 1344 3076 40656 3110
<< via1 >>
rect 4478 38390 4530 38442
rect 4582 38390 4634 38442
rect 4686 38390 4738 38442
rect 35198 38390 35250 38442
rect 35302 38390 35354 38442
rect 35406 38390 35458 38442
rect 14814 38222 14866 38274
rect 18622 38222 18674 38274
rect 25566 38222 25618 38274
rect 21870 38110 21922 38162
rect 14254 37998 14306 38050
rect 17614 37998 17666 38050
rect 20750 37998 20802 38050
rect 24558 37998 24610 38050
rect 19838 37606 19890 37658
rect 19942 37606 19994 37658
rect 20046 37606 20098 37658
rect 15262 37438 15314 37490
rect 22430 37438 22482 37490
rect 26238 37438 26290 37490
rect 14254 37214 14306 37266
rect 25566 37214 25618 37266
rect 4478 36822 4530 36874
rect 4582 36822 4634 36874
rect 4686 36822 4738 36874
rect 35198 36822 35250 36874
rect 35302 36822 35354 36874
rect 35406 36822 35458 36874
rect 19838 36038 19890 36090
rect 19942 36038 19994 36090
rect 20046 36038 20098 36090
rect 4478 35254 4530 35306
rect 4582 35254 4634 35306
rect 4686 35254 4738 35306
rect 35198 35254 35250 35306
rect 35302 35254 35354 35306
rect 35406 35254 35458 35306
rect 19838 34470 19890 34522
rect 19942 34470 19994 34522
rect 20046 34470 20098 34522
rect 4478 33686 4530 33738
rect 4582 33686 4634 33738
rect 4686 33686 4738 33738
rect 35198 33686 35250 33738
rect 35302 33686 35354 33738
rect 35406 33686 35458 33738
rect 19838 32902 19890 32954
rect 19942 32902 19994 32954
rect 20046 32902 20098 32954
rect 4478 32118 4530 32170
rect 4582 32118 4634 32170
rect 4686 32118 4738 32170
rect 35198 32118 35250 32170
rect 35302 32118 35354 32170
rect 35406 32118 35458 32170
rect 19838 31334 19890 31386
rect 19942 31334 19994 31386
rect 20046 31334 20098 31386
rect 4478 30550 4530 30602
rect 4582 30550 4634 30602
rect 4686 30550 4738 30602
rect 35198 30550 35250 30602
rect 35302 30550 35354 30602
rect 35406 30550 35458 30602
rect 19838 29766 19890 29818
rect 19942 29766 19994 29818
rect 20046 29766 20098 29818
rect 4478 28982 4530 29034
rect 4582 28982 4634 29034
rect 4686 28982 4738 29034
rect 35198 28982 35250 29034
rect 35302 28982 35354 29034
rect 35406 28982 35458 29034
rect 19518 28702 19570 28754
rect 16718 28590 16770 28642
rect 19966 28590 20018 28642
rect 17390 28478 17442 28530
rect 13806 28366 13858 28418
rect 19838 28198 19890 28250
rect 19942 28198 19994 28250
rect 20046 28198 20098 28250
rect 17502 28030 17554 28082
rect 17950 27918 18002 27970
rect 10782 27806 10834 27858
rect 14030 27806 14082 27858
rect 18286 27806 18338 27858
rect 20190 27806 20242 27858
rect 23550 27806 23602 27858
rect 11454 27694 11506 27746
rect 13582 27694 13634 27746
rect 14702 27694 14754 27746
rect 16830 27694 16882 27746
rect 20862 27694 20914 27746
rect 22990 27694 23042 27746
rect 4478 27414 4530 27466
rect 4582 27414 4634 27466
rect 4686 27414 4738 27466
rect 35198 27414 35250 27466
rect 35302 27414 35354 27466
rect 35406 27414 35458 27466
rect 15150 27246 15202 27298
rect 15934 27246 15986 27298
rect 1934 27134 1986 27186
rect 16046 27134 16098 27186
rect 16942 27134 16994 27186
rect 21422 27134 21474 27186
rect 25566 27134 25618 27186
rect 26014 27134 26066 27186
rect 40014 27134 40066 27186
rect 4286 27022 4338 27074
rect 14702 27022 14754 27074
rect 15038 27022 15090 27074
rect 16718 27022 16770 27074
rect 22654 27022 22706 27074
rect 37662 27022 37714 27074
rect 13806 26910 13858 26962
rect 13918 26910 13970 26962
rect 14142 26910 14194 26962
rect 14366 26910 14418 26962
rect 16942 26910 16994 26962
rect 17166 26910 17218 26962
rect 17390 26910 17442 26962
rect 18958 26910 19010 26962
rect 19294 26910 19346 26962
rect 21310 26910 21362 26962
rect 21758 26910 21810 26962
rect 23438 26910 23490 26962
rect 27134 26910 27186 26962
rect 27582 26910 27634 26962
rect 27694 26910 27746 26962
rect 15150 26798 15202 26850
rect 21534 26798 21586 26850
rect 26798 26798 26850 26850
rect 27022 26798 27074 26850
rect 27358 26798 27410 26850
rect 19838 26630 19890 26682
rect 19942 26630 19994 26682
rect 20046 26630 20098 26682
rect 20750 26462 20802 26514
rect 23774 26462 23826 26514
rect 14814 26350 14866 26402
rect 14926 26350 14978 26402
rect 18622 26350 18674 26402
rect 19742 26350 19794 26402
rect 19854 26350 19906 26402
rect 20078 26350 20130 26402
rect 21982 26350 22034 26402
rect 22878 26350 22930 26402
rect 14254 26238 14306 26290
rect 14590 26238 14642 26290
rect 18958 26238 19010 26290
rect 20190 26238 20242 26290
rect 20638 26238 20690 26290
rect 20974 26238 21026 26290
rect 21198 26238 21250 26290
rect 21422 26238 21474 26290
rect 21758 26238 21810 26290
rect 22766 26238 22818 26290
rect 23102 26238 23154 26290
rect 23214 26238 23266 26290
rect 23550 26238 23602 26290
rect 25566 26238 25618 26290
rect 37662 26238 37714 26290
rect 11454 26126 11506 26178
rect 13582 26126 13634 26178
rect 15374 26126 15426 26178
rect 18174 26126 18226 26178
rect 18734 26126 18786 26178
rect 26238 26126 26290 26178
rect 28366 26126 28418 26178
rect 28814 26126 28866 26178
rect 18286 26014 18338 26066
rect 19182 26014 19234 26066
rect 19294 26014 19346 26066
rect 20750 26014 20802 26066
rect 22094 26014 22146 26066
rect 23438 26014 23490 26066
rect 40014 26014 40066 26066
rect 4478 25846 4530 25898
rect 4582 25846 4634 25898
rect 4686 25846 4738 25898
rect 35198 25846 35250 25898
rect 35302 25846 35354 25898
rect 35406 25846 35458 25898
rect 21758 25678 21810 25730
rect 13694 25566 13746 25618
rect 18846 25566 18898 25618
rect 19294 25566 19346 25618
rect 21534 25566 21586 25618
rect 26462 25566 26514 25618
rect 28590 25566 28642 25618
rect 29262 25566 29314 25618
rect 13806 25454 13858 25506
rect 14254 25454 14306 25506
rect 19182 25454 19234 25506
rect 19630 25454 19682 25506
rect 22318 25454 22370 25506
rect 25678 25454 25730 25506
rect 13582 25342 13634 25394
rect 17950 25342 18002 25394
rect 18286 25342 18338 25394
rect 18510 25342 18562 25394
rect 19854 25342 19906 25394
rect 21310 25342 21362 25394
rect 21982 25342 22034 25394
rect 18062 25230 18114 25282
rect 18734 25230 18786 25282
rect 19406 25230 19458 25282
rect 20414 25230 20466 25282
rect 20750 25230 20802 25282
rect 21870 25230 21922 25282
rect 19838 25062 19890 25114
rect 19942 25062 19994 25114
rect 20046 25062 20098 25114
rect 17390 24894 17442 24946
rect 19406 24894 19458 24946
rect 26014 24894 26066 24946
rect 26238 24894 26290 24946
rect 27582 24894 27634 24946
rect 27806 24894 27858 24946
rect 18286 24782 18338 24834
rect 20638 24782 20690 24834
rect 26350 24782 26402 24834
rect 17614 24670 17666 24722
rect 18398 24670 18450 24722
rect 19070 24670 19122 24722
rect 20414 24670 20466 24722
rect 27918 24670 27970 24722
rect 18286 24446 18338 24498
rect 4478 24278 4530 24330
rect 4582 24278 4634 24330
rect 4686 24278 4738 24330
rect 35198 24278 35250 24330
rect 35302 24278 35354 24330
rect 35406 24278 35458 24330
rect 13694 24110 13746 24162
rect 1934 23998 1986 24050
rect 40014 23998 40066 24050
rect 4286 23886 4338 23938
rect 37662 23886 37714 23938
rect 13694 23774 13746 23826
rect 13806 23774 13858 23826
rect 14254 23774 14306 23826
rect 14366 23774 14418 23826
rect 18174 23774 18226 23826
rect 18510 23774 18562 23826
rect 14030 23662 14082 23714
rect 16606 23662 16658 23714
rect 18398 23662 18450 23714
rect 26126 23662 26178 23714
rect 26462 23662 26514 23714
rect 37326 23662 37378 23714
rect 19838 23494 19890 23546
rect 19942 23494 19994 23546
rect 20046 23494 20098 23546
rect 14366 23326 14418 23378
rect 17614 23326 17666 23378
rect 18510 23326 18562 23378
rect 19854 23326 19906 23378
rect 13134 23214 13186 23266
rect 15598 23214 15650 23266
rect 17726 23214 17778 23266
rect 18846 23214 18898 23266
rect 19630 23214 19682 23266
rect 21198 23214 21250 23266
rect 13918 23102 13970 23154
rect 15374 23102 15426 23154
rect 16046 23102 16098 23154
rect 18286 23102 18338 23154
rect 19070 23102 19122 23154
rect 19518 23102 19570 23154
rect 20190 23102 20242 23154
rect 20526 23102 20578 23154
rect 20638 23102 20690 23154
rect 21870 23102 21922 23154
rect 37886 23102 37938 23154
rect 11006 22990 11058 23042
rect 16718 22990 16770 23042
rect 16830 22990 16882 23042
rect 17502 22990 17554 23042
rect 20302 22990 20354 23042
rect 21086 22990 21138 23042
rect 22542 22990 22594 23042
rect 24670 22990 24722 23042
rect 25342 22990 25394 23042
rect 15934 22878 15986 22930
rect 21422 22878 21474 22930
rect 40014 22878 40066 22930
rect 4478 22710 4530 22762
rect 4582 22710 4634 22762
rect 4686 22710 4738 22762
rect 35198 22710 35250 22762
rect 35302 22710 35354 22762
rect 35406 22710 35458 22762
rect 17278 22542 17330 22594
rect 17950 22542 18002 22594
rect 18846 22542 18898 22594
rect 20526 22542 20578 22594
rect 20862 22542 20914 22594
rect 28254 22542 28306 22594
rect 16382 22430 16434 22482
rect 22766 22430 22818 22482
rect 26798 22430 26850 22482
rect 40014 22430 40066 22482
rect 13582 22318 13634 22370
rect 16942 22318 16994 22370
rect 18398 22318 18450 22370
rect 19630 22318 19682 22370
rect 20750 22318 20802 22370
rect 21534 22318 21586 22370
rect 22318 22318 22370 22370
rect 22542 22318 22594 22370
rect 23998 22318 24050 22370
rect 27806 22318 27858 22370
rect 29374 22318 29426 22370
rect 37662 22318 37714 22370
rect 14254 22206 14306 22258
rect 17614 22206 17666 22258
rect 17838 22206 17890 22258
rect 18958 22206 19010 22258
rect 19742 22206 19794 22258
rect 21310 22206 21362 22258
rect 24670 22206 24722 22258
rect 28142 22206 28194 22258
rect 17166 22094 17218 22146
rect 20190 22094 20242 22146
rect 27246 22094 27298 22146
rect 27470 22094 27522 22146
rect 27694 22094 27746 22146
rect 28254 22094 28306 22146
rect 29598 22094 29650 22146
rect 19838 21926 19890 21978
rect 19942 21926 19994 21978
rect 20046 21926 20098 21978
rect 14590 21758 14642 21810
rect 15262 21758 15314 21810
rect 15934 21758 15986 21810
rect 18398 21758 18450 21810
rect 25454 21758 25506 21810
rect 14926 21646 14978 21698
rect 17950 21646 18002 21698
rect 18174 21646 18226 21698
rect 25342 21646 25394 21698
rect 25566 21646 25618 21698
rect 27806 21646 27858 21698
rect 11342 21534 11394 21586
rect 12014 21534 12066 21586
rect 15710 21534 15762 21586
rect 16382 21534 16434 21586
rect 16830 21534 16882 21586
rect 18622 21534 18674 21586
rect 19070 21534 19122 21586
rect 25230 21534 25282 21586
rect 26014 21534 26066 21586
rect 27022 21534 27074 21586
rect 37662 21534 37714 21586
rect 14142 21422 14194 21474
rect 22878 21422 22930 21474
rect 26686 21422 26738 21474
rect 29934 21422 29986 21474
rect 40014 21422 40066 21474
rect 4478 21142 4530 21194
rect 4582 21142 4634 21194
rect 4686 21142 4738 21194
rect 35198 21142 35250 21194
rect 35302 21142 35354 21194
rect 35406 21142 35458 21194
rect 22542 20862 22594 20914
rect 27022 20862 27074 20914
rect 14366 20750 14418 20802
rect 20078 20750 20130 20802
rect 21758 20750 21810 20802
rect 22878 20750 22930 20802
rect 14590 20638 14642 20690
rect 14702 20638 14754 20690
rect 15710 20638 15762 20690
rect 21982 20638 22034 20690
rect 22094 20638 22146 20690
rect 22318 20638 22370 20690
rect 21534 20526 21586 20578
rect 19838 20358 19890 20410
rect 19942 20358 19994 20410
rect 20046 20358 20098 20410
rect 18174 20190 18226 20242
rect 18622 20190 18674 20242
rect 18846 20190 18898 20242
rect 20190 20190 20242 20242
rect 21422 20190 21474 20242
rect 22542 20190 22594 20242
rect 25902 20190 25954 20242
rect 26014 20190 26066 20242
rect 19854 20078 19906 20130
rect 19966 20078 20018 20130
rect 20750 20078 20802 20130
rect 21758 20078 21810 20130
rect 22654 20078 22706 20130
rect 22766 20078 22818 20130
rect 22990 20078 23042 20130
rect 23662 20078 23714 20130
rect 18062 19966 18114 20018
rect 18734 19966 18786 20018
rect 19294 19966 19346 20018
rect 20974 19966 21026 20018
rect 22430 19966 22482 20018
rect 23438 19966 23490 20018
rect 23774 19966 23826 20018
rect 25342 19966 25394 20018
rect 25678 19966 25730 20018
rect 26350 19966 26402 20018
rect 37662 19966 37714 20018
rect 17726 19854 17778 19906
rect 27022 19854 27074 19906
rect 29150 19854 29202 19906
rect 29598 19854 29650 19906
rect 20638 19742 20690 19794
rect 40014 19742 40066 19794
rect 4478 19574 4530 19626
rect 4582 19574 4634 19626
rect 4686 19574 4738 19626
rect 35198 19574 35250 19626
rect 35302 19574 35354 19626
rect 35406 19574 35458 19626
rect 19406 19406 19458 19458
rect 22206 19406 22258 19458
rect 26798 19406 26850 19458
rect 15262 19294 15314 19346
rect 40014 19294 40066 19346
rect 14702 19182 14754 19234
rect 16942 19182 16994 19234
rect 17502 19182 17554 19234
rect 18398 19182 18450 19234
rect 18734 19182 18786 19234
rect 19742 19182 19794 19234
rect 20526 19182 20578 19234
rect 21310 19182 21362 19234
rect 25342 19182 25394 19234
rect 25678 19182 25730 19234
rect 37886 19182 37938 19234
rect 17166 19070 17218 19122
rect 17614 19070 17666 19122
rect 18958 19070 19010 19122
rect 19294 19070 19346 19122
rect 20078 19070 20130 19122
rect 21646 19070 21698 19122
rect 22430 19070 22482 19122
rect 25118 19070 25170 19122
rect 25902 19070 25954 19122
rect 26014 19070 26066 19122
rect 26238 19070 26290 19122
rect 14478 18958 14530 19010
rect 20750 18958 20802 19010
rect 22318 18958 22370 19010
rect 24894 18958 24946 19010
rect 25006 18958 25058 19010
rect 26462 18958 26514 19010
rect 26686 18958 26738 19010
rect 19838 18790 19890 18842
rect 19942 18790 19994 18842
rect 20046 18790 20098 18842
rect 15934 18622 15986 18674
rect 16830 18622 16882 18674
rect 17838 18622 17890 18674
rect 18174 18622 18226 18674
rect 21646 18622 21698 18674
rect 22990 18622 23042 18674
rect 24110 18622 24162 18674
rect 24558 18622 24610 18674
rect 19070 18510 19122 18562
rect 19182 18510 19234 18562
rect 21982 18510 22034 18562
rect 23886 18510 23938 18562
rect 12238 18398 12290 18450
rect 15374 18398 15426 18450
rect 17502 18398 17554 18450
rect 18510 18398 18562 18450
rect 18734 18398 18786 18450
rect 19406 18398 19458 18450
rect 19854 18398 19906 18450
rect 20190 18398 20242 18450
rect 20750 18398 20802 18450
rect 21198 18398 21250 18450
rect 21758 18398 21810 18450
rect 22542 18398 22594 18450
rect 23214 18398 23266 18450
rect 23550 18398 23602 18450
rect 24446 18398 24498 18450
rect 24782 18398 24834 18450
rect 25342 18398 25394 18450
rect 28590 18398 28642 18450
rect 37662 18398 37714 18450
rect 12910 18286 12962 18338
rect 15038 18286 15090 18338
rect 16270 18286 16322 18338
rect 22766 18286 22818 18338
rect 23102 18286 23154 18338
rect 26014 18286 26066 18338
rect 28142 18286 28194 18338
rect 15598 18174 15650 18226
rect 16494 18174 16546 18226
rect 20190 18174 20242 18226
rect 21422 18174 21474 18226
rect 22318 18174 22370 18226
rect 24222 18174 24274 18226
rect 40014 18174 40066 18226
rect 4478 18006 4530 18058
rect 4582 18006 4634 18058
rect 4686 18006 4738 18058
rect 35198 18006 35250 18058
rect 35302 18006 35354 18058
rect 35406 18006 35458 18058
rect 18622 17838 18674 17890
rect 28030 17838 28082 17890
rect 14254 17726 14306 17778
rect 22766 17726 22818 17778
rect 24894 17726 24946 17778
rect 14926 17614 14978 17666
rect 15150 17614 15202 17666
rect 15598 17614 15650 17666
rect 16718 17614 16770 17666
rect 17614 17614 17666 17666
rect 19294 17614 19346 17666
rect 19406 17614 19458 17666
rect 20078 17614 20130 17666
rect 21982 17614 22034 17666
rect 25454 17614 25506 17666
rect 25790 17614 25842 17666
rect 26574 17614 26626 17666
rect 27022 17614 27074 17666
rect 15934 17502 15986 17554
rect 17054 17502 17106 17554
rect 18510 17502 18562 17554
rect 18958 17502 19010 17554
rect 20302 17502 20354 17554
rect 25230 17502 25282 17554
rect 17390 17390 17442 17442
rect 19070 17390 19122 17442
rect 25342 17390 25394 17442
rect 26798 17390 26850 17442
rect 26910 17390 26962 17442
rect 27134 17390 27186 17442
rect 27918 17390 27970 17442
rect 40014 17726 40066 17778
rect 28366 17614 28418 17666
rect 28478 17614 28530 17666
rect 37662 17614 37714 17666
rect 19838 17222 19890 17274
rect 19942 17222 19994 17274
rect 20046 17222 20098 17274
rect 15486 17054 15538 17106
rect 23998 17054 24050 17106
rect 25342 17054 25394 17106
rect 26238 17054 26290 17106
rect 12910 16942 12962 16994
rect 24110 16942 24162 16994
rect 27358 16942 27410 16994
rect 12238 16830 12290 16882
rect 26574 16830 26626 16882
rect 15038 16718 15090 16770
rect 29486 16718 29538 16770
rect 4478 16438 4530 16490
rect 4582 16438 4634 16490
rect 4686 16438 4738 16490
rect 35198 16438 35250 16490
rect 35302 16438 35354 16490
rect 35406 16438 35458 16490
rect 19838 15654 19890 15706
rect 19942 15654 19994 15706
rect 20046 15654 20098 15706
rect 25678 15486 25730 15538
rect 26126 15486 26178 15538
rect 15486 15374 15538 15426
rect 15710 15374 15762 15426
rect 18174 15374 18226 15426
rect 18734 15374 18786 15426
rect 19294 15374 19346 15426
rect 19630 15374 19682 15426
rect 21870 15374 21922 15426
rect 22206 15374 22258 15426
rect 16494 15262 16546 15314
rect 18846 15262 18898 15314
rect 19070 15262 19122 15314
rect 22430 15262 22482 15314
rect 25902 15262 25954 15314
rect 37662 15262 37714 15314
rect 15822 15150 15874 15202
rect 16158 15150 16210 15202
rect 16270 15150 16322 15202
rect 18398 15150 18450 15202
rect 19854 15150 19906 15202
rect 26014 15150 26066 15202
rect 40014 15150 40066 15202
rect 18062 15038 18114 15090
rect 20190 15038 20242 15090
rect 21758 15038 21810 15090
rect 4478 14870 4530 14922
rect 4582 14870 4634 14922
rect 4686 14870 4738 14922
rect 35198 14870 35250 14922
rect 35302 14870 35354 14922
rect 35406 14870 35458 14922
rect 17054 14590 17106 14642
rect 19182 14590 19234 14642
rect 23326 14590 23378 14642
rect 25678 14590 25730 14642
rect 27806 14590 27858 14642
rect 28254 14590 28306 14642
rect 16270 14478 16322 14530
rect 19630 14478 19682 14530
rect 19854 14478 19906 14530
rect 20190 14478 20242 14530
rect 21310 14478 21362 14530
rect 21870 14478 21922 14530
rect 22206 14478 22258 14530
rect 22654 14478 22706 14530
rect 22878 14478 22930 14530
rect 23662 14478 23714 14530
rect 25006 14478 25058 14530
rect 19966 14366 20018 14418
rect 23214 14366 23266 14418
rect 23550 14366 23602 14418
rect 19742 14254 19794 14306
rect 20638 14254 20690 14306
rect 21534 14254 21586 14306
rect 21646 14254 21698 14306
rect 21758 14254 21810 14306
rect 22542 14254 22594 14306
rect 19838 14086 19890 14138
rect 19942 14086 19994 14138
rect 20046 14086 20098 14138
rect 16830 13918 16882 13970
rect 21534 13918 21586 13970
rect 26910 13918 26962 13970
rect 13918 13806 13970 13858
rect 18286 13806 18338 13858
rect 21310 13806 21362 13858
rect 22542 13806 22594 13858
rect 25566 13806 25618 13858
rect 27022 13806 27074 13858
rect 13246 13694 13298 13746
rect 17614 13694 17666 13746
rect 21198 13694 21250 13746
rect 21870 13694 21922 13746
rect 25230 13694 25282 13746
rect 16046 13582 16098 13634
rect 20414 13582 20466 13634
rect 24670 13582 24722 13634
rect 4478 13302 4530 13354
rect 4582 13302 4634 13354
rect 4686 13302 4738 13354
rect 35198 13302 35250 13354
rect 35302 13302 35354 13354
rect 35406 13302 35458 13354
rect 20526 13134 20578 13186
rect 16382 13022 16434 13074
rect 22094 13022 22146 13074
rect 24222 13022 24274 13074
rect 25006 13022 25058 13074
rect 25454 13022 25506 13074
rect 20638 12910 20690 12962
rect 21422 12910 21474 12962
rect 20526 12686 20578 12738
rect 19838 12518 19890 12570
rect 19942 12518 19994 12570
rect 20046 12518 20098 12570
rect 4478 11734 4530 11786
rect 4582 11734 4634 11786
rect 4686 11734 4738 11786
rect 35198 11734 35250 11786
rect 35302 11734 35354 11786
rect 35406 11734 35458 11786
rect 19838 10950 19890 11002
rect 19942 10950 19994 11002
rect 20046 10950 20098 11002
rect 4478 10166 4530 10218
rect 4582 10166 4634 10218
rect 4686 10166 4738 10218
rect 35198 10166 35250 10218
rect 35302 10166 35354 10218
rect 35406 10166 35458 10218
rect 19838 9382 19890 9434
rect 19942 9382 19994 9434
rect 20046 9382 20098 9434
rect 4478 8598 4530 8650
rect 4582 8598 4634 8650
rect 4686 8598 4738 8650
rect 35198 8598 35250 8650
rect 35302 8598 35354 8650
rect 35406 8598 35458 8650
rect 19838 7814 19890 7866
rect 19942 7814 19994 7866
rect 20046 7814 20098 7866
rect 4478 7030 4530 7082
rect 4582 7030 4634 7082
rect 4686 7030 4738 7082
rect 35198 7030 35250 7082
rect 35302 7030 35354 7082
rect 35406 7030 35458 7082
rect 19838 6246 19890 6298
rect 19942 6246 19994 6298
rect 20046 6246 20098 6298
rect 4478 5462 4530 5514
rect 4582 5462 4634 5514
rect 4686 5462 4738 5514
rect 35198 5462 35250 5514
rect 35302 5462 35354 5514
rect 35406 5462 35458 5514
rect 19838 4678 19890 4730
rect 19942 4678 19994 4730
rect 20046 4678 20098 4730
rect 17390 4286 17442 4338
rect 20414 4286 20466 4338
rect 25342 4286 25394 4338
rect 18510 4174 18562 4226
rect 21422 4062 21474 4114
rect 26238 4062 26290 4114
rect 4478 3894 4530 3946
rect 4582 3894 4634 3946
rect 4686 3894 4738 3946
rect 35198 3894 35250 3946
rect 35302 3894 35354 3946
rect 35406 3894 35458 3946
rect 25566 3614 25618 3666
rect 18062 3502 18114 3554
rect 23550 3502 23602 3554
rect 24558 3502 24610 3554
rect 19406 3390 19458 3442
rect 22206 3390 22258 3442
rect 19838 3110 19890 3162
rect 19942 3110 19994 3162
rect 20046 3110 20098 3162
<< metal2 >>
rect 14112 41200 14224 42000
rect 14784 41200 14896 42000
rect 17472 41200 17584 42000
rect 19488 41200 19600 42000
rect 22176 41200 22288 42000
rect 22848 41200 22960 42000
rect 24864 41200 24976 42000
rect 4476 38444 4740 38454
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4476 38378 4740 38388
rect 14140 37492 14196 41200
rect 14812 38274 14868 41200
rect 14812 38222 14814 38274
rect 14866 38222 14868 38274
rect 14812 38210 14868 38222
rect 17500 38276 17556 41200
rect 17500 38210 17556 38220
rect 18620 38276 18676 38286
rect 18620 38182 18676 38220
rect 19516 38164 19572 41200
rect 19516 38098 19572 38108
rect 21868 38164 21924 38174
rect 21868 38070 21924 38108
rect 14252 38052 14308 38062
rect 14252 38050 14420 38052
rect 14252 37998 14254 38050
rect 14306 37998 14420 38050
rect 14252 37996 14420 37998
rect 14252 37986 14308 37996
rect 14140 37426 14196 37436
rect 14252 37266 14308 37278
rect 14252 37214 14254 37266
rect 14306 37214 14308 37266
rect 4476 36876 4740 36886
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4476 36810 4740 36820
rect 4476 35308 4740 35318
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4476 35242 4740 35252
rect 4476 33740 4740 33750
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4476 33674 4740 33684
rect 4476 32172 4740 32182
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4476 32106 4740 32116
rect 14252 31948 14308 37214
rect 13580 31892 14308 31948
rect 4476 30604 4740 30614
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4476 30538 4740 30548
rect 4476 29036 4740 29046
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4476 28970 4740 28980
rect 10780 27860 10836 27870
rect 10780 27766 10836 27804
rect 11452 27746 11508 27758
rect 11452 27694 11454 27746
rect 11506 27694 11508 27746
rect 4172 27636 4228 27646
rect 1932 27186 1988 27198
rect 1932 27134 1934 27186
rect 1986 27134 1988 27186
rect 1932 26292 1988 27134
rect 1932 26226 1988 26236
rect 1932 24050 1988 24062
rect 1932 23998 1934 24050
rect 1986 23998 1988 24050
rect 1932 23604 1988 23998
rect 1932 23538 1988 23548
rect 4172 22932 4228 27580
rect 4476 27468 4740 27478
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4476 27402 4740 27412
rect 11452 27300 11508 27694
rect 13580 27748 13636 31892
rect 14028 28644 14084 28654
rect 13804 28420 13860 28430
rect 14028 28420 14084 28588
rect 13804 28418 14084 28420
rect 13804 28366 13806 28418
rect 13858 28366 14084 28418
rect 13804 28364 14084 28366
rect 13804 28354 13860 28364
rect 14028 27860 14084 28364
rect 13580 27746 13972 27748
rect 13580 27694 13582 27746
rect 13634 27694 13972 27746
rect 13580 27692 13972 27694
rect 13580 27682 13636 27692
rect 11452 27234 11508 27244
rect 13804 27188 13860 27198
rect 4284 27074 4340 27086
rect 4284 27022 4286 27074
rect 4338 27022 4340 27074
rect 4284 26180 4340 27022
rect 13804 26962 13860 27132
rect 13804 26910 13806 26962
rect 13858 26910 13860 26962
rect 13804 26404 13860 26910
rect 13916 27076 13972 27692
rect 13916 26962 13972 27020
rect 13916 26910 13918 26962
rect 13970 26910 13972 26962
rect 13916 26898 13972 26910
rect 13468 26348 13860 26404
rect 4284 26114 4340 26124
rect 11452 26180 11508 26190
rect 11452 26086 11508 26124
rect 4476 25900 4740 25910
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4476 25834 4740 25844
rect 13468 24948 13524 26348
rect 14028 26292 14084 27804
rect 14140 26964 14196 26974
rect 14140 26870 14196 26908
rect 14364 26962 14420 37996
rect 17612 38050 17668 38062
rect 17612 37998 17614 38050
rect 17666 37998 17668 38050
rect 15260 37492 15316 37502
rect 15260 37398 15316 37436
rect 17612 31948 17668 37998
rect 19628 38052 19684 38062
rect 19628 35308 19684 37996
rect 20748 38052 20804 38062
rect 20748 37958 20804 37996
rect 19836 37660 20100 37670
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 19836 37594 20100 37604
rect 22204 37492 22260 41200
rect 22876 38276 22932 41200
rect 22876 38210 22932 38220
rect 24556 38050 24612 38062
rect 24556 37998 24558 38050
rect 24610 37998 24612 38050
rect 22428 37492 22484 37502
rect 22204 37490 22484 37492
rect 22204 37438 22430 37490
rect 22482 37438 22484 37490
rect 22204 37436 22484 37438
rect 22428 37426 22484 37436
rect 19836 36092 20100 36102
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 19836 36026 20100 36036
rect 16828 31892 17668 31948
rect 19516 35252 19684 35308
rect 16716 28644 16772 28654
rect 16716 28550 16772 28588
rect 14700 27748 14756 27758
rect 14700 27654 14756 27692
rect 15932 27748 15988 27758
rect 15148 27300 15204 27310
rect 15148 27206 15204 27244
rect 15932 27298 15988 27692
rect 15932 27246 15934 27298
rect 15986 27246 15988 27298
rect 15932 27234 15988 27246
rect 16828 27746 16884 31892
rect 19516 28754 19572 35252
rect 19836 34524 20100 34534
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 19836 34458 20100 34468
rect 19836 32956 20100 32966
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 19836 32890 20100 32900
rect 19836 31388 20100 31398
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 19836 31322 20100 31332
rect 19836 29820 20100 29830
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 19836 29754 20100 29764
rect 19516 28702 19518 28754
rect 19570 28702 19572 28754
rect 17500 28644 17556 28654
rect 17388 28530 17444 28542
rect 17388 28478 17390 28530
rect 17442 28478 17444 28530
rect 17388 27860 17444 28478
rect 17500 28082 17556 28588
rect 17500 28030 17502 28082
rect 17554 28030 17556 28082
rect 17500 28018 17556 28030
rect 17948 27970 18004 27982
rect 17948 27918 17950 27970
rect 18002 27918 18004 27970
rect 17948 27860 18004 27918
rect 17388 27804 18004 27860
rect 18284 27858 18340 27870
rect 18284 27806 18286 27858
rect 18338 27806 18340 27858
rect 16828 27694 16830 27746
rect 16882 27694 16884 27746
rect 14812 27188 14868 27198
rect 14476 27076 14532 27086
rect 14700 27076 14756 27086
rect 14532 27074 14756 27076
rect 14532 27022 14702 27074
rect 14754 27022 14756 27074
rect 14532 27020 14756 27022
rect 14476 27010 14532 27020
rect 14700 27010 14756 27020
rect 14364 26910 14366 26962
rect 14418 26910 14420 26962
rect 14364 26898 14420 26910
rect 14812 26628 14868 27132
rect 16044 27188 16100 27198
rect 16044 27094 16100 27132
rect 15036 27074 15092 27086
rect 15036 27022 15038 27074
rect 15090 27022 15092 27074
rect 14924 26964 14980 26974
rect 15036 26964 15092 27022
rect 16716 27076 16772 27114
rect 16716 27010 16772 27020
rect 14980 26908 15092 26964
rect 16828 26964 16884 27694
rect 16940 27188 16996 27198
rect 16940 27094 16996 27132
rect 16940 26964 16996 26974
rect 16828 26962 16996 26964
rect 16828 26910 16942 26962
rect 16994 26910 16996 26962
rect 16828 26908 16996 26910
rect 14924 26898 14980 26908
rect 16940 26898 16996 26908
rect 17164 26964 17220 26974
rect 17164 26870 17220 26908
rect 17388 26964 17444 26974
rect 17388 26962 18004 26964
rect 17388 26910 17390 26962
rect 17442 26910 18004 26962
rect 17388 26908 18004 26910
rect 17388 26898 17444 26908
rect 15148 26852 15204 26862
rect 15148 26758 15204 26796
rect 14812 26572 14980 26628
rect 14812 26402 14868 26414
rect 14812 26350 14814 26402
rect 14866 26350 14868 26402
rect 14252 26292 14308 26302
rect 14588 26292 14644 26302
rect 14028 26236 14252 26292
rect 14252 26198 14308 26236
rect 14364 26290 14644 26292
rect 14364 26238 14590 26290
rect 14642 26238 14644 26290
rect 14364 26236 14644 26238
rect 13580 26178 13636 26190
rect 13580 26126 13582 26178
rect 13634 26126 13636 26178
rect 13580 25620 13636 26126
rect 13692 25620 13748 25630
rect 13580 25618 13748 25620
rect 13580 25566 13694 25618
rect 13746 25566 13748 25618
rect 13580 25564 13748 25566
rect 13692 25554 13748 25564
rect 13804 25508 13860 25518
rect 13804 25414 13860 25452
rect 14252 25508 14308 25518
rect 14364 25508 14420 26236
rect 14588 26226 14644 26236
rect 14812 26180 14868 26350
rect 14924 26402 14980 26572
rect 14924 26350 14926 26402
rect 14978 26350 14980 26402
rect 14924 26338 14980 26350
rect 14812 26114 14868 26124
rect 15372 26180 15428 26190
rect 14252 25506 14420 25508
rect 14252 25454 14254 25506
rect 14306 25454 14420 25506
rect 14252 25452 14420 25454
rect 14252 25442 14308 25452
rect 13580 25396 13636 25406
rect 13580 25302 13636 25340
rect 4476 24332 4740 24342
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4476 24266 4740 24276
rect 4284 23940 4340 23950
rect 4284 23846 4340 23884
rect 11004 23940 11060 23950
rect 11004 23042 11060 23884
rect 13132 23716 13188 23726
rect 13132 23266 13188 23660
rect 13468 23604 13524 24892
rect 13692 24164 13748 24174
rect 13692 24162 13860 24164
rect 13692 24110 13694 24162
rect 13746 24110 13860 24162
rect 13692 24108 13860 24110
rect 13692 24098 13748 24108
rect 13804 24052 13860 24108
rect 13804 23996 14308 24052
rect 13692 23940 13748 23950
rect 13692 23826 13748 23884
rect 13692 23774 13694 23826
rect 13746 23774 13748 23826
rect 13692 23762 13748 23774
rect 13804 23826 13860 23838
rect 13804 23774 13806 23826
rect 13858 23774 13860 23826
rect 13804 23604 13860 23774
rect 14252 23826 14308 23996
rect 14252 23774 14254 23826
rect 14306 23774 14308 23826
rect 14252 23762 14308 23774
rect 14364 23828 14420 23838
rect 14364 23734 14420 23772
rect 14700 23828 14756 23838
rect 14028 23716 14084 23726
rect 14028 23622 14084 23660
rect 13468 23548 13860 23604
rect 14364 23604 14420 23614
rect 14364 23380 14420 23548
rect 13132 23214 13134 23266
rect 13186 23214 13188 23266
rect 13132 23202 13188 23214
rect 13916 23378 14644 23380
rect 13916 23326 14366 23378
rect 14418 23326 14644 23378
rect 13916 23324 14644 23326
rect 13916 23156 13972 23324
rect 14364 23314 14420 23324
rect 11004 22990 11006 23042
rect 11058 22990 11060 23042
rect 11004 22978 11060 22990
rect 13580 23154 13972 23156
rect 13580 23102 13918 23154
rect 13970 23102 13972 23154
rect 13580 23100 13972 23102
rect 4172 22866 4228 22876
rect 4476 22764 4740 22774
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4476 22698 4740 22708
rect 13580 22370 13636 23100
rect 13916 23090 13972 23100
rect 14140 23156 14196 23166
rect 13580 22318 13582 22370
rect 13634 22318 13636 22370
rect 13580 22306 13636 22318
rect 11340 21812 11396 21822
rect 11340 21586 11396 21756
rect 11340 21534 11342 21586
rect 11394 21534 11396 21586
rect 11340 21522 11396 21534
rect 12012 21588 12068 21598
rect 12012 21494 12068 21532
rect 14140 21474 14196 23100
rect 14252 22260 14308 22270
rect 14252 22258 14420 22260
rect 14252 22206 14254 22258
rect 14306 22206 14420 22258
rect 14252 22204 14420 22206
rect 14252 22194 14308 22204
rect 14140 21422 14142 21474
rect 14194 21422 14196 21474
rect 14140 21410 14196 21422
rect 4476 21196 4740 21206
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4476 21130 4740 21140
rect 14364 20802 14420 22204
rect 14588 21812 14644 23324
rect 14588 21718 14644 21756
rect 14700 21588 14756 23772
rect 15372 23716 15428 26124
rect 17948 25394 18004 26908
rect 18284 26908 18340 27806
rect 18956 26964 19012 26974
rect 19292 26962 19348 26974
rect 19292 26910 19294 26962
rect 19346 26910 19348 26962
rect 19292 26908 19348 26910
rect 18284 26852 18676 26908
rect 18620 26402 18676 26852
rect 18620 26350 18622 26402
rect 18674 26350 18676 26402
rect 18620 26338 18676 26350
rect 18956 26292 19012 26908
rect 18956 26198 19012 26236
rect 19068 26852 19348 26908
rect 19068 26404 19124 26852
rect 19516 26516 19572 28702
rect 19964 28644 20020 28654
rect 19964 28550 20020 28588
rect 19836 28252 20100 28262
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 19836 28186 20100 28196
rect 20188 27860 20244 27870
rect 20188 27766 20244 27804
rect 22652 27860 22708 27870
rect 20860 27748 20916 27758
rect 20748 27746 20916 27748
rect 20748 27694 20862 27746
rect 20914 27694 20916 27746
rect 20748 27692 20916 27694
rect 19836 26684 20100 26694
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 19836 26618 20100 26628
rect 19516 26450 19572 26460
rect 19964 26516 20020 26526
rect 17948 25342 17950 25394
rect 18002 25342 18004 25394
rect 17388 24948 17444 24958
rect 17948 24948 18004 25342
rect 18172 26178 18228 26190
rect 18172 26126 18174 26178
rect 18226 26126 18228 26178
rect 17388 24854 17444 24892
rect 17500 24892 18004 24948
rect 18060 25282 18116 25294
rect 18060 25230 18062 25282
rect 18114 25230 18116 25282
rect 17500 24724 17556 24892
rect 17388 24668 17556 24724
rect 17612 24722 17668 24734
rect 17612 24670 17614 24722
rect 17666 24670 17668 24722
rect 15372 23650 15428 23660
rect 16604 23716 16660 23726
rect 16604 23622 16660 23660
rect 15596 23268 15652 23278
rect 15596 23174 15652 23212
rect 15372 23156 15428 23166
rect 15372 23062 15428 23100
rect 16044 23156 16100 23166
rect 16044 23062 16100 23100
rect 16716 23042 16772 23054
rect 16716 22990 16718 23042
rect 16770 22990 16772 23042
rect 15932 22932 15988 22942
rect 15708 22930 15988 22932
rect 15708 22878 15934 22930
rect 15986 22878 15988 22930
rect 15708 22876 15988 22878
rect 15260 22708 15316 22718
rect 15260 21812 15316 22652
rect 15148 21810 15316 21812
rect 15148 21758 15262 21810
rect 15314 21758 15316 21810
rect 15148 21756 15316 21758
rect 14924 21700 14980 21710
rect 14924 21606 14980 21644
rect 14364 20750 14366 20802
rect 14418 20750 14420 20802
rect 14364 20738 14420 20750
rect 14588 21532 14756 21588
rect 14588 20690 14644 21532
rect 14588 20638 14590 20690
rect 14642 20638 14644 20690
rect 14588 20626 14644 20638
rect 14700 20690 14756 20702
rect 14700 20638 14702 20690
rect 14754 20638 14756 20690
rect 4476 19628 4740 19638
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4476 19562 4740 19572
rect 14700 19460 14756 20638
rect 14700 19394 14756 19404
rect 14700 19236 14756 19246
rect 14252 19234 14756 19236
rect 14252 19182 14702 19234
rect 14754 19182 14756 19234
rect 14252 19180 14756 19182
rect 12236 18450 12292 18462
rect 12236 18398 12238 18450
rect 12290 18398 12292 18450
rect 4476 18060 4740 18070
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4476 17994 4740 18004
rect 12236 16884 12292 18398
rect 12908 18338 12964 18350
rect 12908 18286 12910 18338
rect 12962 18286 12964 18338
rect 12908 17780 12964 18286
rect 12908 17714 12964 17724
rect 14252 17778 14308 19180
rect 14700 19170 14756 19180
rect 14252 17726 14254 17778
rect 14306 17726 14308 17778
rect 14252 17714 14308 17726
rect 14476 19010 14532 19022
rect 14476 18958 14478 19010
rect 14530 18958 14532 19010
rect 14476 18228 14532 18958
rect 15148 18452 15204 21756
rect 15260 21746 15316 21756
rect 15372 21812 15428 21822
rect 15372 20692 15428 21756
rect 15708 21700 15764 22876
rect 15932 22866 15988 22876
rect 16380 22482 16436 22494
rect 16380 22430 16382 22482
rect 16434 22430 16436 22482
rect 16380 22372 16436 22430
rect 16716 22372 16772 22990
rect 16828 23044 16884 23054
rect 16828 22950 16884 22988
rect 17276 22596 17332 22606
rect 17276 22502 17332 22540
rect 16940 22372 16996 22382
rect 16380 22370 16996 22372
rect 16380 22318 16942 22370
rect 16994 22318 16996 22370
rect 16380 22316 16996 22318
rect 15932 21812 15988 21822
rect 15932 21718 15988 21756
rect 15708 21586 15764 21644
rect 15708 21534 15710 21586
rect 15762 21534 15764 21586
rect 15708 21522 15764 21534
rect 16380 21586 16436 22316
rect 16940 22260 16996 22316
rect 16940 22194 16996 22204
rect 17164 22146 17220 22158
rect 17164 22094 17166 22146
rect 17218 22094 17220 22146
rect 17164 21812 17220 22094
rect 17164 21746 17220 21756
rect 16380 21534 16382 21586
rect 16434 21534 16436 21586
rect 16380 21522 16436 21534
rect 16828 21700 16884 21710
rect 16828 21586 16884 21644
rect 16828 21534 16830 21586
rect 16882 21534 16884 21586
rect 16828 21522 16884 21534
rect 17388 21476 17444 24668
rect 17612 23716 17668 24670
rect 17612 23378 17668 23660
rect 17612 23326 17614 23378
rect 17666 23326 17668 23378
rect 17612 23314 17668 23326
rect 17948 24724 18004 24734
rect 18060 24724 18116 25230
rect 18004 24668 18116 24724
rect 18172 25284 18228 26126
rect 18732 26180 18788 26190
rect 18732 26086 18788 26124
rect 18284 26068 18340 26078
rect 18284 25974 18340 26012
rect 18732 25956 18788 25966
rect 18620 25844 18676 25854
rect 18284 25396 18340 25406
rect 18284 25302 18340 25340
rect 18508 25394 18564 25406
rect 18508 25342 18510 25394
rect 18562 25342 18564 25394
rect 17724 23266 17780 23278
rect 17724 23214 17726 23266
rect 17778 23214 17780 23266
rect 17500 23044 17556 23054
rect 17500 22950 17556 22988
rect 17612 22260 17668 22270
rect 17612 22166 17668 22204
rect 17724 21812 17780 23214
rect 17836 23268 17892 23278
rect 17836 22260 17892 23212
rect 17948 22594 18004 24668
rect 18172 24500 18228 25228
rect 18508 24948 18564 25342
rect 18284 24892 18564 24948
rect 18284 24836 18340 24892
rect 18284 24742 18340 24780
rect 18396 24724 18452 24734
rect 18396 24630 18452 24668
rect 18284 24500 18340 24510
rect 18620 24500 18676 25788
rect 18732 25508 18788 25900
rect 19068 25844 19124 26348
rect 19740 26402 19796 26414
rect 19740 26350 19742 26402
rect 19794 26350 19796 26402
rect 19740 26292 19796 26350
rect 19852 26404 19908 26414
rect 19852 26310 19908 26348
rect 19628 26236 19796 26292
rect 19180 26068 19236 26078
rect 19180 25974 19236 26012
rect 19292 26066 19348 26078
rect 19292 26014 19294 26066
rect 19346 26014 19348 26066
rect 19068 25778 19124 25788
rect 18732 25284 18788 25452
rect 18844 25618 18900 25630
rect 18844 25566 18846 25618
rect 18898 25566 18900 25618
rect 18844 25284 18900 25566
rect 19292 25618 19348 26014
rect 19628 26068 19684 26236
rect 19628 26002 19684 26012
rect 19292 25566 19294 25618
rect 19346 25566 19348 25618
rect 19292 25554 19348 25566
rect 19180 25508 19236 25546
rect 19180 25442 19236 25452
rect 19628 25506 19684 25518
rect 19964 25508 20020 26460
rect 20748 26514 20804 27692
rect 20860 27682 20916 27692
rect 21756 27748 21812 27758
rect 21420 27188 21476 27198
rect 20748 26462 20750 26514
rect 20802 26462 20804 26514
rect 20748 26450 20804 26462
rect 20860 27186 21476 27188
rect 20860 27134 21422 27186
rect 21474 27134 21476 27186
rect 20860 27132 21476 27134
rect 20076 26404 20132 26414
rect 20076 26402 20244 26404
rect 20076 26350 20078 26402
rect 20130 26350 20244 26402
rect 20076 26348 20244 26350
rect 20076 26338 20132 26348
rect 20188 26290 20244 26348
rect 20188 26238 20190 26290
rect 20242 26238 20244 26290
rect 20188 26226 20244 26238
rect 20636 26292 20692 26302
rect 20860 26292 20916 27132
rect 21420 27122 21476 27132
rect 21308 26962 21364 26974
rect 21308 26910 21310 26962
rect 21362 26910 21364 26962
rect 21308 26908 21364 26910
rect 20972 26852 21364 26908
rect 21756 26962 21812 27692
rect 22652 27074 22708 27804
rect 23548 27860 23604 27870
rect 23548 27766 23604 27804
rect 22988 27748 23044 27758
rect 22988 27654 23044 27692
rect 24556 27748 24612 37998
rect 24892 37492 24948 41200
rect 35196 38444 35460 38454
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35196 38378 35460 38388
rect 25564 38276 25620 38286
rect 25564 38182 25620 38220
rect 24892 37426 24948 37436
rect 26236 37492 26292 37502
rect 26236 37398 26292 37436
rect 25564 37266 25620 37278
rect 25564 37214 25566 37266
rect 25618 37214 25620 37266
rect 24556 27682 24612 27692
rect 25452 27860 25508 27870
rect 22652 27022 22654 27074
rect 22706 27022 22708 27074
rect 22652 27010 22708 27022
rect 21756 26910 21758 26962
rect 21810 26910 21812 26962
rect 21756 26898 21812 26910
rect 23436 26962 23492 26974
rect 23436 26910 23438 26962
rect 23490 26910 23492 26962
rect 20972 26786 21028 26796
rect 21532 26850 21588 26862
rect 21532 26798 21534 26850
rect 21586 26798 21588 26850
rect 21532 26740 21588 26798
rect 21084 26684 21588 26740
rect 22540 26852 22596 26862
rect 20636 26290 20916 26292
rect 20636 26238 20638 26290
rect 20690 26238 20916 26290
rect 20636 26236 20916 26238
rect 20972 26292 21028 26302
rect 20636 26226 20692 26236
rect 20972 26198 21028 26236
rect 20524 26180 20580 26190
rect 20524 26068 20580 26124
rect 20748 26068 20804 26078
rect 20524 26066 20804 26068
rect 20524 26014 20750 26066
rect 20802 26014 20804 26066
rect 20524 26012 20804 26014
rect 20524 25732 20580 26012
rect 20748 26002 20804 26012
rect 21084 25844 21140 26684
rect 21420 26404 21476 26414
rect 20524 25666 20580 25676
rect 20636 25788 21140 25844
rect 21196 26290 21252 26302
rect 21196 26238 21198 26290
rect 21250 26238 21252 26290
rect 21196 26068 21252 26238
rect 21420 26290 21476 26348
rect 21980 26402 22036 26414
rect 21980 26350 21982 26402
rect 22034 26350 22036 26402
rect 21420 26238 21422 26290
rect 21474 26238 21476 26290
rect 21420 26226 21476 26238
rect 21756 26290 21812 26302
rect 21756 26238 21758 26290
rect 21810 26238 21812 26290
rect 21756 26068 21812 26238
rect 21196 26012 21812 26068
rect 19628 25454 19630 25506
rect 19682 25454 19684 25506
rect 19628 25396 19684 25454
rect 19628 25330 19684 25340
rect 19852 25452 20020 25508
rect 19852 25394 19908 25452
rect 19852 25342 19854 25394
rect 19906 25342 19908 25394
rect 19852 25330 19908 25342
rect 19068 25284 19124 25294
rect 18844 25228 19068 25284
rect 18732 25190 18788 25228
rect 19068 25218 19124 25228
rect 19404 25284 19460 25322
rect 19404 25218 19460 25228
rect 20412 25284 20468 25294
rect 20636 25284 20692 25788
rect 21084 25620 21140 25630
rect 20412 25282 20692 25284
rect 20412 25230 20414 25282
rect 20466 25230 20692 25282
rect 20412 25228 20692 25230
rect 20748 25284 20804 25294
rect 19836 25116 20100 25126
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20412 25060 20468 25228
rect 19836 25050 20100 25060
rect 20188 25004 20468 25060
rect 19404 24948 19460 24958
rect 19404 24854 19460 24892
rect 19068 24724 19124 24734
rect 19068 24630 19124 24668
rect 18172 24498 18340 24500
rect 18172 24446 18286 24498
rect 18338 24446 18340 24498
rect 18172 24444 18340 24446
rect 18284 24052 18340 24444
rect 17948 22542 17950 22594
rect 18002 22542 18004 22594
rect 17948 22530 18004 22542
rect 18060 23996 18340 24052
rect 18396 24444 18676 24500
rect 17836 22166 17892 22204
rect 17724 21746 17780 21756
rect 17948 21700 18004 21710
rect 17948 21606 18004 21644
rect 17388 21410 17444 21420
rect 18060 21252 18116 23996
rect 18172 23828 18228 23838
rect 18172 23734 18228 23772
rect 18396 23714 18452 24444
rect 18508 23828 18564 23838
rect 18508 23826 18788 23828
rect 18508 23774 18510 23826
rect 18562 23774 18788 23826
rect 18508 23772 18788 23774
rect 18508 23762 18564 23772
rect 18396 23662 18398 23714
rect 18450 23662 18452 23714
rect 18396 23604 18452 23662
rect 18396 23548 18564 23604
rect 18508 23378 18564 23548
rect 18508 23326 18510 23378
rect 18562 23326 18564 23378
rect 18508 23314 18564 23326
rect 18284 23154 18340 23166
rect 18284 23102 18286 23154
rect 18338 23102 18340 23154
rect 18284 22596 18340 23102
rect 18732 23156 18788 23772
rect 19836 23548 20100 23558
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 19836 23482 20100 23492
rect 19852 23380 19908 23390
rect 20188 23380 20244 25004
rect 20636 24834 20692 24846
rect 20636 24782 20638 24834
rect 20690 24782 20692 24834
rect 19852 23378 20244 23380
rect 19852 23326 19854 23378
rect 19906 23326 20244 23378
rect 19852 23324 20244 23326
rect 20412 24724 20468 24734
rect 19852 23314 19908 23324
rect 18732 23090 18788 23100
rect 18844 23266 18900 23278
rect 18844 23214 18846 23266
rect 18898 23214 18900 23266
rect 18844 22932 18900 23214
rect 19628 23266 19684 23278
rect 19628 23214 19630 23266
rect 19682 23214 19684 23266
rect 19068 23156 19124 23166
rect 19516 23156 19572 23166
rect 19068 23154 19572 23156
rect 19068 23102 19070 23154
rect 19122 23102 19518 23154
rect 19570 23102 19572 23154
rect 19068 23100 19572 23102
rect 19068 23044 19124 23100
rect 19516 23090 19572 23100
rect 19068 22978 19124 22988
rect 18844 22866 18900 22876
rect 19180 22932 19236 22942
rect 18284 22372 18340 22540
rect 18844 22596 18900 22606
rect 18844 22502 18900 22540
rect 18396 22372 18452 22382
rect 18284 22370 18452 22372
rect 18284 22318 18398 22370
rect 18450 22318 18452 22370
rect 18284 22316 18452 22318
rect 18396 22306 18452 22316
rect 19068 22372 19124 22382
rect 18844 22260 18900 22270
rect 18172 21812 18228 21822
rect 18172 21698 18228 21756
rect 18172 21646 18174 21698
rect 18226 21646 18228 21698
rect 18172 21634 18228 21646
rect 18396 21810 18452 21822
rect 18396 21758 18398 21810
rect 18450 21758 18452 21810
rect 17500 21196 18116 21252
rect 18172 21476 18228 21486
rect 15708 20692 15764 20702
rect 15260 20690 15764 20692
rect 15260 20638 15710 20690
rect 15762 20638 15764 20690
rect 15260 20636 15764 20638
rect 15260 19348 15316 20636
rect 15708 20626 15764 20636
rect 17164 19796 17220 19806
rect 15260 19346 15540 19348
rect 15260 19294 15262 19346
rect 15314 19294 15540 19346
rect 15260 19292 15540 19294
rect 15260 19282 15316 19292
rect 15372 18452 15428 18462
rect 15148 18450 15428 18452
rect 15148 18398 15374 18450
rect 15426 18398 15428 18450
rect 15148 18396 15428 18398
rect 15036 18340 15092 18350
rect 12908 16996 12964 17006
rect 12908 16902 12964 16940
rect 14476 16996 14532 18172
rect 14924 18284 15036 18340
rect 14924 17666 14980 18284
rect 15036 18246 15092 18284
rect 15148 17668 15204 17678
rect 14924 17614 14926 17666
rect 14978 17614 14980 17666
rect 14924 17602 14980 17614
rect 15036 17612 15148 17668
rect 14476 16930 14532 16940
rect 12236 16790 12292 16828
rect 15036 16770 15092 17612
rect 15148 17574 15204 17612
rect 15036 16718 15038 16770
rect 15090 16718 15092 16770
rect 15036 16706 15092 16718
rect 15372 17444 15428 18396
rect 4476 16492 4740 16502
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4476 16426 4740 16436
rect 15372 15428 15428 17388
rect 15484 17106 15540 19292
rect 16940 19236 16996 19246
rect 15932 19124 15988 19134
rect 15932 18674 15988 19068
rect 15932 18622 15934 18674
rect 15986 18622 15988 18674
rect 15932 18610 15988 18622
rect 16828 18676 16884 18686
rect 16940 18676 16996 19180
rect 17164 19122 17220 19740
rect 17500 19234 17556 21196
rect 18172 20242 18228 21420
rect 18172 20190 18174 20242
rect 18226 20190 18228 20242
rect 18172 20178 18228 20190
rect 18396 20244 18452 21758
rect 18620 21586 18676 21598
rect 18620 21534 18622 21586
rect 18674 21534 18676 21586
rect 18620 21476 18676 21534
rect 18620 21410 18676 21420
rect 18060 20020 18116 20030
rect 17724 19906 17780 19918
rect 17724 19854 17726 19906
rect 17778 19854 17780 19906
rect 17500 19182 17502 19234
rect 17554 19182 17556 19234
rect 17500 19170 17556 19182
rect 17612 19460 17668 19470
rect 17164 19070 17166 19122
rect 17218 19070 17220 19122
rect 17164 19058 17220 19070
rect 17612 19122 17668 19404
rect 17612 19070 17614 19122
rect 17666 19070 17668 19122
rect 16828 18674 16996 18676
rect 16828 18622 16830 18674
rect 16882 18622 16996 18674
rect 16828 18620 16996 18622
rect 16828 18610 16884 18620
rect 16492 18452 16548 18462
rect 16268 18340 16324 18350
rect 16268 18246 16324 18284
rect 15596 18228 15652 18238
rect 15596 18134 15652 18172
rect 16492 18226 16548 18396
rect 17500 18452 17556 18462
rect 17500 18358 17556 18396
rect 16492 18174 16494 18226
rect 16546 18174 16548 18226
rect 15596 17668 15652 17678
rect 15596 17574 15652 17612
rect 15932 17556 15988 17566
rect 16492 17556 16548 18174
rect 16716 18340 16772 18350
rect 16716 17666 16772 18284
rect 16716 17614 16718 17666
rect 16770 17614 16772 17666
rect 16716 17602 16772 17614
rect 17612 17666 17668 19070
rect 17724 19012 17780 19854
rect 17724 18452 17780 18956
rect 17836 18676 17892 18686
rect 17836 18582 17892 18620
rect 17724 18386 17780 18396
rect 17612 17614 17614 17666
rect 17666 17614 17668 17666
rect 17612 17602 17668 17614
rect 15932 17554 16548 17556
rect 15932 17502 15934 17554
rect 15986 17502 16548 17554
rect 15932 17500 16548 17502
rect 17052 17556 17108 17566
rect 15932 17490 15988 17500
rect 17052 17462 17108 17500
rect 18060 17556 18116 19964
rect 18172 19348 18228 19358
rect 18172 18674 18228 19292
rect 18396 19234 18452 20188
rect 18620 20242 18676 20254
rect 18620 20190 18622 20242
rect 18674 20190 18676 20242
rect 18620 20132 18676 20190
rect 18844 20244 18900 22204
rect 18956 22258 19012 22270
rect 18956 22206 18958 22258
rect 19010 22206 19012 22258
rect 18956 20468 19012 22206
rect 19068 21586 19124 22316
rect 19068 21534 19070 21586
rect 19122 21534 19124 21586
rect 19068 21522 19124 21534
rect 18956 20402 19012 20412
rect 18844 20242 19124 20244
rect 18844 20190 18846 20242
rect 18898 20190 19124 20242
rect 18844 20188 19124 20190
rect 18844 20178 18900 20188
rect 18396 19182 18398 19234
rect 18450 19182 18452 19234
rect 18396 19170 18452 19182
rect 18508 20076 18676 20132
rect 19068 20132 19124 20188
rect 18508 19236 18564 20076
rect 19068 20066 19124 20076
rect 18732 20020 18788 20030
rect 18620 20018 18788 20020
rect 18620 19966 18734 20018
rect 18786 19966 18788 20018
rect 18620 19964 18788 19966
rect 18620 19460 18676 19964
rect 18732 19954 18788 19964
rect 19180 19796 19236 22876
rect 19628 22708 19684 23214
rect 19628 22642 19684 22652
rect 20188 23154 20244 23166
rect 20188 23102 20190 23154
rect 20242 23102 20244 23154
rect 20188 22708 20244 23102
rect 20188 22642 20244 22652
rect 20300 23042 20356 23054
rect 20300 22990 20302 23042
rect 20354 22990 20356 23042
rect 19628 22370 19684 22382
rect 19628 22318 19630 22370
rect 19682 22318 19684 22370
rect 19628 22260 19684 22318
rect 19292 22204 19684 22260
rect 19740 22258 19796 22270
rect 19740 22206 19742 22258
rect 19794 22206 19796 22258
rect 19292 21700 19348 22204
rect 19740 22148 19796 22206
rect 19628 22092 19796 22148
rect 20188 22146 20244 22158
rect 20188 22094 20190 22146
rect 20242 22094 20244 22146
rect 19628 21924 19684 22092
rect 20188 22036 20244 22094
rect 19836 21980 20100 21990
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20188 21970 20244 21980
rect 19836 21914 20100 21924
rect 19628 21858 19684 21868
rect 19292 20018 19348 21644
rect 20188 21812 20244 21822
rect 20076 20804 20132 20814
rect 20076 20710 20132 20748
rect 19292 19966 19294 20018
rect 19346 19966 19348 20018
rect 19292 19908 19348 19966
rect 19292 19842 19348 19852
rect 19404 20468 19460 20478
rect 19460 20412 19684 20468
rect 18620 19394 18676 19404
rect 18844 19740 19236 19796
rect 18172 18622 18174 18674
rect 18226 18622 18228 18674
rect 18172 18564 18228 18622
rect 18172 18498 18228 18508
rect 18508 18450 18564 19180
rect 18732 19234 18788 19246
rect 18732 19182 18734 19234
rect 18786 19182 18788 19234
rect 18732 19124 18788 19182
rect 18732 19058 18788 19068
rect 18508 18398 18510 18450
rect 18562 18398 18564 18450
rect 18508 18386 18564 18398
rect 18620 18452 18676 18462
rect 18620 17890 18676 18396
rect 18732 18452 18788 18462
rect 18844 18452 18900 19740
rect 19404 19460 19460 20412
rect 19628 20132 19684 20412
rect 19836 20412 20100 20422
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 19836 20346 20100 20356
rect 20188 20242 20244 21756
rect 20300 21588 20356 22990
rect 20300 21522 20356 21532
rect 20188 20190 20190 20242
rect 20242 20190 20244 20242
rect 20188 20178 20244 20190
rect 19852 20132 19908 20142
rect 19628 20130 19908 20132
rect 19628 20078 19854 20130
rect 19906 20078 19908 20130
rect 19628 20076 19908 20078
rect 19068 19458 19460 19460
rect 19068 19406 19406 19458
rect 19458 19406 19460 19458
rect 19068 19404 19460 19406
rect 18732 18450 18900 18452
rect 18732 18398 18734 18450
rect 18786 18398 18900 18450
rect 18732 18396 18900 18398
rect 18732 18386 18788 18396
rect 18620 17838 18622 17890
rect 18674 17838 18676 17890
rect 18620 17826 18676 17838
rect 18844 17668 18900 18396
rect 18956 19122 19012 19134
rect 18956 19070 18958 19122
rect 19010 19070 19012 19122
rect 18956 17780 19012 19070
rect 19068 18562 19124 19404
rect 19404 19394 19460 19404
rect 19740 19234 19796 20076
rect 19852 20066 19908 20076
rect 19964 20130 20020 20142
rect 19964 20078 19966 20130
rect 20018 20078 20020 20130
rect 19964 20020 20020 20078
rect 19964 19954 20020 19964
rect 19740 19182 19742 19234
rect 19794 19182 19796 19234
rect 19740 19170 19796 19182
rect 19292 19122 19348 19134
rect 19292 19070 19294 19122
rect 19346 19070 19348 19122
rect 19292 19012 19348 19070
rect 19292 18946 19348 18956
rect 19404 19124 19460 19134
rect 19404 18788 19460 19068
rect 20076 19124 20132 19134
rect 20076 19030 20132 19068
rect 19292 18732 19460 18788
rect 19836 18844 20100 18854
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 19836 18778 20100 18788
rect 19068 18510 19070 18562
rect 19122 18510 19124 18562
rect 19068 18498 19124 18510
rect 19180 18562 19236 18574
rect 19180 18510 19182 18562
rect 19234 18510 19236 18562
rect 19180 18452 19236 18510
rect 19180 18386 19236 18396
rect 18956 17724 19236 17780
rect 18844 17602 18900 17612
rect 18060 17490 18116 17500
rect 18508 17556 18564 17566
rect 18508 17462 18564 17500
rect 18956 17554 19012 17566
rect 18956 17502 18958 17554
rect 19010 17502 19012 17554
rect 15484 17054 15486 17106
rect 15538 17054 15540 17106
rect 15484 16884 15540 17054
rect 17388 17442 17444 17454
rect 17388 17390 17390 17442
rect 17442 17390 17444 17442
rect 15540 16828 15652 16884
rect 15484 16818 15540 16828
rect 15484 15428 15540 15438
rect 15372 15426 15540 15428
rect 15372 15374 15486 15426
rect 15538 15374 15540 15426
rect 15372 15372 15540 15374
rect 15484 15362 15540 15372
rect 13916 15204 13972 15214
rect 4476 14924 4740 14934
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4476 14858 4740 14868
rect 13356 14308 13412 14318
rect 13244 14252 13356 14308
rect 13244 13746 13300 14252
rect 13356 14242 13412 14252
rect 13916 13858 13972 15148
rect 15484 14308 15540 14318
rect 15596 14308 15652 16828
rect 15540 14252 15652 14308
rect 15708 15426 15764 15438
rect 15708 15374 15710 15426
rect 15762 15374 15764 15426
rect 15484 14242 15540 14252
rect 13916 13806 13918 13858
rect 13970 13806 13972 13858
rect 13916 13794 13972 13806
rect 13244 13694 13246 13746
rect 13298 13694 13300 13746
rect 13244 13682 13300 13694
rect 15708 13636 15764 15374
rect 16492 15428 16548 15438
rect 16492 15314 16548 15372
rect 17388 15428 17444 17390
rect 18956 17444 19012 17502
rect 18956 17378 19012 17388
rect 19068 17442 19124 17454
rect 19068 17390 19070 17442
rect 19122 17390 19124 17442
rect 19068 16324 19124 17390
rect 18732 16268 19124 16324
rect 17388 15362 17444 15372
rect 18172 15426 18228 15438
rect 18172 15374 18174 15426
rect 18226 15374 18228 15426
rect 16492 15262 16494 15314
rect 16546 15262 16548 15314
rect 16492 15250 16548 15262
rect 18172 15316 18228 15374
rect 18732 15426 18788 16268
rect 18732 15374 18734 15426
rect 18786 15374 18788 15426
rect 18732 15362 18788 15374
rect 18172 15250 18228 15260
rect 18844 15316 18900 15326
rect 15820 15204 15876 15214
rect 16156 15204 16212 15214
rect 15820 15202 16212 15204
rect 15820 15150 15822 15202
rect 15874 15150 16158 15202
rect 16210 15150 16212 15202
rect 15820 15148 16212 15150
rect 15820 15138 15876 15148
rect 16156 15138 16212 15148
rect 16268 15204 16324 15242
rect 16268 15138 16324 15148
rect 18396 15204 18452 15242
rect 18844 15222 18900 15260
rect 19068 15314 19124 15326
rect 19068 15262 19070 15314
rect 19122 15262 19124 15314
rect 18396 15138 18452 15148
rect 18060 15092 18116 15102
rect 17052 15090 18116 15092
rect 17052 15038 18062 15090
rect 18114 15038 18116 15090
rect 17052 15036 18116 15038
rect 17052 14642 17108 15036
rect 18060 15026 18116 15036
rect 17052 14590 17054 14642
rect 17106 14590 17108 14642
rect 17052 14578 17108 14590
rect 19068 14644 19124 15262
rect 19180 15148 19236 17724
rect 19292 17666 19348 18732
rect 19852 18676 19908 18686
rect 19404 18450 19460 18462
rect 19404 18398 19406 18450
rect 19458 18398 19460 18450
rect 19404 18340 19460 18398
rect 19852 18450 19908 18620
rect 20300 18676 20356 18686
rect 20412 18676 20468 24668
rect 20636 23492 20692 24782
rect 20636 23426 20692 23436
rect 20524 23156 20580 23166
rect 20524 22594 20580 23100
rect 20524 22542 20526 22594
rect 20578 22542 20580 22594
rect 20524 22530 20580 22542
rect 20636 23154 20692 23166
rect 20636 23102 20638 23154
rect 20690 23102 20692 23154
rect 20636 20132 20692 23102
rect 20748 22708 20804 25228
rect 21084 23042 21140 25564
rect 21196 25396 21252 26012
rect 21980 25956 22036 26350
rect 22540 26292 22596 26796
rect 23436 26628 23492 26910
rect 23100 26572 23492 26628
rect 22876 26402 22932 26414
rect 22876 26350 22878 26402
rect 22930 26350 22932 26402
rect 22428 26236 22540 26292
rect 21980 25890 22036 25900
rect 22092 26066 22148 26078
rect 22092 26014 22094 26066
rect 22146 26014 22148 26066
rect 21532 25844 21588 25854
rect 21532 25618 21588 25788
rect 21756 25732 21812 25742
rect 21756 25638 21812 25676
rect 21532 25566 21534 25618
rect 21586 25566 21588 25618
rect 21532 25554 21588 25566
rect 21644 25620 21700 25630
rect 21308 25396 21364 25406
rect 21196 25394 21364 25396
rect 21196 25342 21310 25394
rect 21362 25342 21364 25394
rect 21196 25340 21364 25342
rect 21308 23492 21364 25340
rect 21644 25284 21700 25564
rect 21980 25394 22036 25406
rect 21980 25342 21982 25394
rect 22034 25342 22036 25394
rect 21644 25218 21700 25228
rect 21868 25284 21924 25294
rect 21868 25190 21924 25228
rect 21980 23604 22036 25342
rect 22092 24948 22148 26014
rect 22316 25508 22372 25518
rect 22316 25414 22372 25452
rect 22092 24882 22148 24892
rect 21308 23426 21364 23436
rect 21756 23548 22036 23604
rect 21196 23268 21252 23278
rect 21196 23266 21588 23268
rect 21196 23214 21198 23266
rect 21250 23214 21588 23266
rect 21196 23212 21588 23214
rect 21196 23202 21252 23212
rect 21084 22990 21086 23042
rect 21138 22990 21140 23042
rect 21084 22978 21140 22990
rect 21420 22932 21476 22942
rect 20748 22642 20804 22652
rect 21308 22708 21364 22718
rect 20860 22594 20916 22606
rect 20860 22542 20862 22594
rect 20914 22542 20916 22594
rect 20748 22372 20804 22382
rect 20748 22278 20804 22316
rect 20748 20132 20804 20142
rect 20636 20130 20804 20132
rect 20636 20078 20750 20130
rect 20802 20078 20804 20130
rect 20636 20076 20804 20078
rect 20748 20066 20804 20076
rect 20524 20020 20580 20030
rect 20524 19234 20580 19964
rect 20636 19796 20692 19806
rect 20860 19796 20916 22542
rect 21308 22258 21364 22652
rect 21420 22372 21476 22876
rect 21420 22306 21476 22316
rect 21532 22372 21588 23212
rect 21644 22708 21700 22718
rect 21756 22708 21812 23548
rect 21980 23380 22036 23390
rect 21700 22652 21812 22708
rect 21868 23154 21924 23166
rect 21868 23102 21870 23154
rect 21922 23102 21924 23154
rect 21644 22642 21700 22652
rect 21532 22370 21812 22372
rect 21532 22318 21534 22370
rect 21586 22318 21812 22370
rect 21532 22316 21812 22318
rect 21532 22306 21588 22316
rect 21308 22206 21310 22258
rect 21362 22206 21364 22258
rect 21308 21812 21364 22206
rect 21308 21746 21364 21756
rect 21756 20804 21812 22316
rect 21868 21924 21924 23102
rect 21868 21858 21924 21868
rect 21420 20802 21812 20804
rect 21420 20750 21758 20802
rect 21810 20750 21812 20802
rect 21420 20748 21812 20750
rect 21420 20242 21476 20748
rect 21756 20738 21812 20748
rect 21980 20690 22036 23324
rect 22428 23156 22484 26236
rect 22540 26226 22596 26236
rect 22764 26290 22820 26302
rect 22764 26238 22766 26290
rect 22818 26238 22820 26290
rect 22764 25284 22820 26238
rect 22876 26068 22932 26350
rect 23100 26290 23156 26572
rect 23772 26516 23828 26526
rect 23772 26422 23828 26460
rect 23100 26238 23102 26290
rect 23154 26238 23156 26290
rect 23100 26226 23156 26238
rect 23212 26292 23268 26302
rect 23212 26198 23268 26236
rect 23548 26290 23604 26302
rect 23548 26238 23550 26290
rect 23602 26238 23604 26290
rect 23436 26068 23492 26078
rect 22876 26066 23492 26068
rect 22876 26014 23438 26066
rect 23490 26014 23492 26066
rect 22876 26012 23492 26014
rect 23436 26002 23492 26012
rect 23548 25620 23604 26238
rect 25452 26292 25508 27804
rect 25564 27186 25620 37214
rect 35196 36876 35460 36886
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35196 36810 35460 36820
rect 35196 35308 35460 35318
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35196 35242 35460 35252
rect 35196 33740 35460 33750
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35196 33674 35460 33684
rect 35196 32172 35460 32182
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35196 32106 35460 32116
rect 35196 30604 35460 30614
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35196 30538 35460 30548
rect 35196 29036 35460 29046
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35196 28970 35460 28980
rect 25564 27134 25566 27186
rect 25618 27134 25620 27186
rect 25564 26516 25620 27134
rect 26012 27860 26068 27870
rect 26012 27186 26068 27804
rect 35196 27468 35460 27478
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35196 27402 35460 27412
rect 26012 27134 26014 27186
rect 26066 27134 26068 27186
rect 26012 27122 26068 27134
rect 40012 27186 40068 27198
rect 40012 27134 40014 27186
rect 40066 27134 40068 27186
rect 27580 27076 27636 27086
rect 27132 26964 27188 26974
rect 27132 26962 27300 26964
rect 27132 26910 27134 26962
rect 27186 26910 27300 26962
rect 27132 26908 27300 26910
rect 27132 26898 27188 26908
rect 25564 26450 25620 26460
rect 26348 26852 26404 26862
rect 25564 26292 25620 26302
rect 25452 26290 25732 26292
rect 25452 26238 25566 26290
rect 25618 26238 25732 26290
rect 25452 26236 25732 26238
rect 25564 26226 25620 26236
rect 23548 25554 23604 25564
rect 25676 26180 25732 26236
rect 26236 26180 26292 26190
rect 23436 25508 23492 25518
rect 23436 25284 23492 25452
rect 25676 25506 25732 26124
rect 25676 25454 25678 25506
rect 25730 25454 25732 25506
rect 23436 25228 23604 25284
rect 22764 25218 22820 25228
rect 22316 23100 22484 23156
rect 22316 22596 22372 23100
rect 22540 23044 22596 23054
rect 22316 22370 22372 22540
rect 22316 22318 22318 22370
rect 22370 22318 22372 22370
rect 22316 22306 22372 22318
rect 22428 23042 22596 23044
rect 22428 22990 22542 23042
rect 22594 22990 22596 23042
rect 22428 22988 22596 22990
rect 22316 22036 22372 22046
rect 22204 21980 22316 22036
rect 21980 20638 21982 20690
rect 22034 20638 22036 20690
rect 21980 20626 22036 20638
rect 22092 20690 22148 20702
rect 22092 20638 22094 20690
rect 22146 20638 22148 20690
rect 21532 20580 21588 20590
rect 21532 20486 21588 20524
rect 21420 20190 21422 20242
rect 21474 20190 21476 20242
rect 20972 20020 21028 20030
rect 20972 19926 21028 19964
rect 21420 20020 21476 20190
rect 21756 20132 21812 20142
rect 21756 20038 21812 20076
rect 21420 19954 21476 19964
rect 22092 20020 22148 20638
rect 21308 19908 21364 19918
rect 20692 19740 20916 19796
rect 21196 19796 21252 19806
rect 20636 19702 20692 19740
rect 20524 19182 20526 19234
rect 20578 19182 20580 19234
rect 20524 19170 20580 19182
rect 20748 19012 20804 19022
rect 20748 19010 20916 19012
rect 20748 18958 20750 19010
rect 20802 18958 20916 19010
rect 20748 18956 20916 18958
rect 20748 18946 20804 18956
rect 20356 18620 20468 18676
rect 20748 18788 20804 18798
rect 20300 18610 20356 18620
rect 19852 18398 19854 18450
rect 19906 18398 19908 18450
rect 19852 18386 19908 18398
rect 20076 18452 20132 18462
rect 20188 18452 20244 18462
rect 20132 18450 20244 18452
rect 20132 18398 20190 18450
rect 20242 18398 20244 18450
rect 20132 18396 20244 18398
rect 19404 18274 19460 18284
rect 19628 18228 19684 18238
rect 19292 17614 19294 17666
rect 19346 17614 19348 17666
rect 19292 17602 19348 17614
rect 19404 17668 19460 17678
rect 19404 17574 19460 17612
rect 19292 15428 19348 15438
rect 19628 15428 19684 18172
rect 20076 17666 20132 18396
rect 20188 18386 20244 18396
rect 20748 18450 20804 18732
rect 20748 18398 20750 18450
rect 20802 18398 20804 18450
rect 20748 18386 20804 18398
rect 20860 18452 20916 18956
rect 20860 18386 20916 18396
rect 21196 18450 21252 19740
rect 21308 19234 21364 19852
rect 21308 19182 21310 19234
rect 21362 19182 21364 19234
rect 21308 19170 21364 19182
rect 21644 19124 21700 19134
rect 22092 19124 22148 19964
rect 21644 19122 22148 19124
rect 21644 19070 21646 19122
rect 21698 19070 22148 19122
rect 21644 19068 22148 19070
rect 22204 20356 22260 21980
rect 22316 21970 22372 21980
rect 22316 21812 22372 21822
rect 22316 20690 22372 21756
rect 22316 20638 22318 20690
rect 22370 20638 22372 20690
rect 22316 20580 22372 20638
rect 22316 20514 22372 20524
rect 22204 20300 22372 20356
rect 22204 19458 22260 20300
rect 22316 20020 22372 20300
rect 22428 20244 22484 22988
rect 22540 22978 22596 22988
rect 22764 22484 22820 22494
rect 22764 22482 23044 22484
rect 22764 22430 22766 22482
rect 22818 22430 23044 22482
rect 22764 22428 23044 22430
rect 22764 22418 22820 22428
rect 22540 22372 22596 22382
rect 22540 22278 22596 22316
rect 22988 21588 23044 22428
rect 22876 21474 22932 21486
rect 22876 21422 22878 21474
rect 22930 21422 22932 21474
rect 22540 20916 22596 20926
rect 22540 20914 22820 20916
rect 22540 20862 22542 20914
rect 22594 20862 22820 20914
rect 22540 20860 22820 20862
rect 22540 20850 22596 20860
rect 22540 20244 22596 20254
rect 22428 20242 22596 20244
rect 22428 20190 22542 20242
rect 22594 20190 22596 20242
rect 22428 20188 22596 20190
rect 22540 20178 22596 20188
rect 22652 20130 22708 20142
rect 22652 20078 22654 20130
rect 22706 20078 22708 20130
rect 22428 20020 22484 20030
rect 22316 20018 22484 20020
rect 22316 19966 22430 20018
rect 22482 19966 22484 20018
rect 22316 19964 22484 19966
rect 22428 19954 22484 19964
rect 22204 19406 22206 19458
rect 22258 19406 22260 19458
rect 21644 19058 21700 19068
rect 21756 18900 21812 18910
rect 21196 18398 21198 18450
rect 21250 18398 21252 18450
rect 21196 18386 21252 18398
rect 21644 18674 21700 18686
rect 21644 18622 21646 18674
rect 21698 18622 21700 18674
rect 20188 18228 20244 18238
rect 20188 18134 20244 18172
rect 21420 18228 21476 18238
rect 21420 18134 21476 18172
rect 21644 18116 21700 18622
rect 21756 18450 21812 18844
rect 22204 18788 22260 19406
rect 22428 19124 22484 19134
rect 22652 19124 22708 20078
rect 22764 20130 22820 20860
rect 22876 20804 22932 21422
rect 22876 20710 22932 20748
rect 22764 20078 22766 20130
rect 22818 20078 22820 20130
rect 22764 20066 22820 20078
rect 22988 20130 23044 21532
rect 22988 20078 22990 20130
rect 23042 20078 23044 20130
rect 22988 20066 23044 20078
rect 23436 20020 23492 20030
rect 22484 19068 22708 19124
rect 23212 20018 23492 20020
rect 23212 19966 23438 20018
rect 23490 19966 23492 20018
rect 23212 19964 23492 19966
rect 22428 19030 22484 19068
rect 22204 18722 22260 18732
rect 22316 19010 22372 19022
rect 22316 18958 22318 19010
rect 22370 18958 22372 19010
rect 22092 18676 22148 18686
rect 21756 18398 21758 18450
rect 21810 18398 21812 18450
rect 21756 18386 21812 18398
rect 21980 18562 22036 18574
rect 21980 18510 21982 18562
rect 22034 18510 22036 18562
rect 21980 18340 22036 18510
rect 21980 18274 22036 18284
rect 22092 18228 22148 18620
rect 22316 18452 22372 18958
rect 22316 18396 22484 18452
rect 22316 18228 22372 18238
rect 22092 18226 22372 18228
rect 22092 18174 22318 18226
rect 22370 18174 22372 18226
rect 22092 18172 22372 18174
rect 22316 18162 22372 18172
rect 21756 18116 21812 18126
rect 21644 18060 21756 18116
rect 21756 18050 21812 18060
rect 20076 17614 20078 17666
rect 20130 17614 20132 17666
rect 20076 17602 20132 17614
rect 20300 17780 20356 17790
rect 20300 17554 20356 17724
rect 20300 17502 20302 17554
rect 20354 17502 20356 17554
rect 20300 17490 20356 17502
rect 21980 17666 22036 17678
rect 21980 17614 21982 17666
rect 22034 17614 22036 17666
rect 19836 17276 20100 17286
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 19836 17210 20100 17220
rect 21980 17108 22036 17614
rect 19836 15708 20100 15718
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 19836 15642 20100 15652
rect 19292 15426 19684 15428
rect 19292 15374 19294 15426
rect 19346 15374 19630 15426
rect 19682 15374 19684 15426
rect 19292 15372 19684 15374
rect 19292 15362 19348 15372
rect 19628 15362 19684 15372
rect 21868 15428 21924 15438
rect 21868 15334 21924 15372
rect 19852 15202 19908 15214
rect 19852 15150 19854 15202
rect 19906 15150 19908 15202
rect 19852 15148 19908 15150
rect 19180 15092 19908 15148
rect 19964 15204 20020 15214
rect 19180 14644 19236 14654
rect 19068 14642 19236 14644
rect 19068 14590 19182 14642
rect 19234 14590 19236 14642
rect 19068 14588 19236 14590
rect 16268 14530 16324 14542
rect 16268 14478 16270 14530
rect 16322 14478 16324 14530
rect 16268 14308 16324 14478
rect 18284 14532 18340 14542
rect 16828 14308 16884 14318
rect 16324 14252 16436 14308
rect 16268 14242 16324 14252
rect 16044 13636 16100 13646
rect 15708 13634 16100 13636
rect 15708 13582 16046 13634
rect 16098 13582 16100 13634
rect 15708 13580 16100 13582
rect 4476 13356 4740 13366
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4476 13290 4740 13300
rect 16044 12516 16100 13580
rect 16380 13074 16436 14252
rect 16828 13970 16884 14252
rect 16828 13918 16830 13970
rect 16882 13918 16884 13970
rect 16828 13906 16884 13918
rect 17612 14308 17668 14318
rect 17612 13746 17668 14252
rect 18284 13858 18340 14476
rect 18284 13806 18286 13858
rect 18338 13806 18340 13858
rect 18284 13794 18340 13806
rect 17612 13694 17614 13746
rect 17666 13694 17668 13746
rect 17612 13682 17668 13694
rect 16380 13022 16382 13074
rect 16434 13022 16436 13074
rect 16380 13010 16436 13022
rect 16044 12450 16100 12460
rect 17388 12516 17444 12526
rect 4476 11788 4740 11798
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4476 11722 4740 11732
rect 4476 10220 4740 10230
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4476 10154 4740 10164
rect 4476 8652 4740 8662
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4476 8586 4740 8596
rect 4476 7084 4740 7094
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4476 7018 4740 7028
rect 4476 5516 4740 5526
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4476 5450 4740 5460
rect 17388 4338 17444 12460
rect 17388 4286 17390 4338
rect 17442 4286 17444 4338
rect 17388 4274 17444 4286
rect 16156 4228 16212 4238
rect 4476 3948 4740 3958
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4476 3882 4740 3892
rect 16156 800 16212 4172
rect 18508 4228 18564 4238
rect 18508 4134 18564 4172
rect 18060 3556 18116 3566
rect 18060 3462 18116 3500
rect 19180 3556 19236 14588
rect 19628 14532 19684 14542
rect 19740 14532 19796 15092
rect 19964 14868 20020 15148
rect 20188 15092 20244 15102
rect 20188 15090 21364 15092
rect 20188 15038 20190 15090
rect 20242 15038 21364 15090
rect 20188 15036 21364 15038
rect 20188 15026 20244 15036
rect 19964 14812 20244 14868
rect 19628 14530 19796 14532
rect 19628 14478 19630 14530
rect 19682 14478 19796 14530
rect 19628 14476 19796 14478
rect 19852 14532 19908 14542
rect 19628 14466 19684 14476
rect 19852 14438 19908 14476
rect 20188 14532 20244 14812
rect 20188 14438 20244 14476
rect 21308 14530 21364 15036
rect 21756 15090 21812 15102
rect 21756 15038 21758 15090
rect 21810 15038 21812 15090
rect 21756 14532 21812 15038
rect 21308 14478 21310 14530
rect 21362 14478 21364 14530
rect 21308 14466 21364 14478
rect 21420 14476 21812 14532
rect 21868 14532 21924 14542
rect 19964 14420 20020 14430
rect 19964 14326 20020 14364
rect 21420 14420 21476 14476
rect 21868 14438 21924 14476
rect 19740 14308 19796 14318
rect 19628 14306 19796 14308
rect 19628 14254 19742 14306
rect 19794 14254 19796 14306
rect 19628 14252 19796 14254
rect 19628 13188 19684 14252
rect 19740 14242 19796 14252
rect 20636 14308 20692 14318
rect 21420 14308 21476 14364
rect 20636 14214 20692 14252
rect 21196 14252 21476 14308
rect 21532 14306 21588 14318
rect 21532 14254 21534 14306
rect 21586 14254 21588 14306
rect 19836 14140 20100 14150
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 19836 14074 20100 14084
rect 21196 13746 21252 14252
rect 21532 13970 21588 14254
rect 21532 13918 21534 13970
rect 21586 13918 21588 13970
rect 21532 13906 21588 13918
rect 21644 14306 21700 14318
rect 21644 14254 21646 14306
rect 21698 14254 21700 14306
rect 21308 13860 21364 13870
rect 21308 13766 21364 13804
rect 21196 13694 21198 13746
rect 21250 13694 21252 13746
rect 19628 13122 19684 13132
rect 20412 13634 20468 13646
rect 20412 13582 20414 13634
rect 20466 13582 20468 13634
rect 20412 12740 20468 13582
rect 20524 13188 20580 13198
rect 20524 13094 20580 13132
rect 20636 12964 20692 12974
rect 21196 12964 21252 13694
rect 21644 13524 21700 14254
rect 21756 14308 21812 14318
rect 21756 14214 21812 14252
rect 21868 13748 21924 13758
rect 21980 13748 22036 17052
rect 22204 15426 22260 15438
rect 22204 15374 22206 15426
rect 22258 15374 22260 15426
rect 22204 14532 22260 15374
rect 22204 14438 22260 14476
rect 22428 15314 22484 18396
rect 22540 18450 22596 19068
rect 22988 18676 23044 18686
rect 23212 18676 23268 19964
rect 23436 19954 23492 19964
rect 23548 18900 23604 25228
rect 24668 23044 24724 23054
rect 24556 22988 24668 23044
rect 23996 22370 24052 22382
rect 23996 22318 23998 22370
rect 24050 22318 24052 22370
rect 23996 21924 24052 22318
rect 23996 21858 24052 21868
rect 24556 21812 24612 22988
rect 24668 22950 24724 22988
rect 25340 23044 25396 23054
rect 25676 23044 25732 25454
rect 26012 26178 26292 26180
rect 26012 26126 26238 26178
rect 26290 26126 26292 26178
rect 26012 26124 26292 26126
rect 26012 24946 26068 26124
rect 26236 26114 26292 26124
rect 26012 24894 26014 24946
rect 26066 24894 26068 24946
rect 26012 24882 26068 24894
rect 26236 24948 26292 24958
rect 26236 24854 26292 24892
rect 26348 24834 26404 26796
rect 26796 26850 26852 26862
rect 26796 26798 26798 26850
rect 26850 26798 26852 26850
rect 26460 25620 26516 25630
rect 26796 25620 26852 26798
rect 26460 25618 26852 25620
rect 26460 25566 26462 25618
rect 26514 25566 26852 25618
rect 26460 25564 26852 25566
rect 27020 26850 27076 26862
rect 27020 26798 27022 26850
rect 27074 26798 27076 26850
rect 26460 25554 26516 25564
rect 27020 25508 27076 26798
rect 27244 25732 27300 26908
rect 27580 26962 27636 27020
rect 28364 27076 28420 27086
rect 27580 26910 27582 26962
rect 27634 26910 27636 26962
rect 27580 26898 27636 26910
rect 27692 26962 27748 26974
rect 27692 26910 27694 26962
rect 27746 26910 27748 26962
rect 27356 26852 27412 26862
rect 27356 26758 27412 26796
rect 27244 25676 27636 25732
rect 27020 25442 27076 25452
rect 27580 24946 27636 25676
rect 27580 24894 27582 24946
rect 27634 24894 27636 24946
rect 27580 24882 27636 24894
rect 26348 24782 26350 24834
rect 26402 24782 26404 24834
rect 26348 24770 26404 24782
rect 27692 24724 27748 26910
rect 28364 26178 28420 27020
rect 37660 27076 37716 27086
rect 37660 26982 37716 27020
rect 37660 26290 37716 26302
rect 37660 26238 37662 26290
rect 37714 26238 37716 26290
rect 28364 26126 28366 26178
rect 28418 26126 28420 26178
rect 28364 26114 28420 26126
rect 28812 26180 28868 26190
rect 28868 26124 29316 26180
rect 28812 26086 28868 26124
rect 27804 25620 27860 25630
rect 27804 24946 27860 25564
rect 28588 25620 28644 25630
rect 28588 25526 28644 25564
rect 29260 25618 29316 26124
rect 35196 25900 35460 25910
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35196 25834 35460 25844
rect 29260 25566 29262 25618
rect 29314 25566 29316 25618
rect 29260 25554 29316 25566
rect 37660 25620 37716 26238
rect 40012 26292 40068 27134
rect 40012 26226 40068 26236
rect 37660 25554 37716 25564
rect 40012 26066 40068 26078
rect 40012 26014 40014 26066
rect 40066 26014 40068 26066
rect 40012 25620 40068 26014
rect 40012 25554 40068 25564
rect 27804 24894 27806 24946
rect 27858 24894 27860 24946
rect 27804 24882 27860 24894
rect 27916 24724 27972 24734
rect 27692 24722 27972 24724
rect 27692 24670 27918 24722
rect 27970 24670 27972 24722
rect 27692 24668 27972 24670
rect 26124 23716 26180 23726
rect 26124 23622 26180 23660
rect 26460 23716 26516 23726
rect 26460 23622 26516 23660
rect 27916 23716 27972 24668
rect 35196 24332 35460 24342
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35196 24266 35460 24276
rect 40012 24050 40068 24062
rect 40012 23998 40014 24050
rect 40066 23998 40068 24050
rect 37660 23938 37716 23950
rect 37660 23886 37662 23938
rect 37714 23886 37716 23938
rect 27916 23650 27972 23660
rect 28364 23716 28420 23726
rect 25340 23042 25732 23044
rect 25340 22990 25342 23042
rect 25394 22990 25732 23042
rect 25340 22988 25732 22990
rect 24556 21746 24612 21756
rect 24668 22258 24724 22270
rect 24668 22206 24670 22258
rect 24722 22206 24724 22258
rect 24668 21700 24724 22206
rect 25340 21924 25396 22988
rect 28252 22596 28308 22606
rect 28028 22594 28308 22596
rect 28028 22542 28254 22594
rect 28306 22542 28308 22594
rect 28028 22540 28308 22542
rect 26796 22484 26852 22494
rect 26572 22482 26852 22484
rect 26572 22430 26798 22482
rect 26850 22430 26852 22482
rect 26572 22428 26852 22430
rect 25340 21858 25396 21868
rect 25452 22036 25508 22046
rect 25452 21810 25508 21980
rect 25452 21758 25454 21810
rect 25506 21758 25508 21810
rect 25452 21746 25508 21758
rect 25900 21812 25956 21822
rect 24668 21634 24724 21644
rect 25340 21700 25396 21710
rect 25340 21606 25396 21644
rect 25564 21698 25620 21710
rect 25564 21646 25566 21698
rect 25618 21646 25620 21698
rect 25228 21586 25284 21598
rect 25228 21534 25230 21586
rect 25282 21534 25284 21586
rect 25228 21476 25284 21534
rect 25564 21588 25620 21646
rect 25564 21522 25620 21532
rect 25228 21410 25284 21420
rect 25340 21364 25396 21374
rect 25340 20244 25396 21308
rect 23660 20132 23716 20142
rect 23660 20038 23716 20076
rect 23772 20020 23828 20030
rect 23772 19926 23828 19964
rect 25340 20018 25396 20188
rect 25900 20242 25956 21756
rect 26572 21812 26628 22428
rect 26796 22418 26852 22428
rect 27804 22372 27860 22382
rect 28028 22372 28084 22540
rect 28252 22530 28308 22540
rect 28364 22372 28420 23660
rect 37324 23716 37380 23726
rect 37660 23716 37716 23886
rect 37324 23714 37716 23716
rect 37324 23662 37326 23714
rect 37378 23662 37716 23714
rect 37324 23660 37716 23662
rect 37324 23044 37380 23660
rect 40012 23604 40068 23998
rect 40012 23538 40068 23548
rect 37324 22978 37380 22988
rect 37884 23154 37940 23166
rect 37884 23102 37886 23154
rect 37938 23102 37940 23154
rect 35196 22764 35460 22774
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35196 22698 35460 22708
rect 27804 22370 28084 22372
rect 27804 22318 27806 22370
rect 27858 22318 28084 22370
rect 27804 22316 28084 22318
rect 28140 22316 28420 22372
rect 29372 22370 29428 22382
rect 29372 22318 29374 22370
rect 29426 22318 29428 22370
rect 27804 22306 27860 22316
rect 28140 22258 28196 22316
rect 28140 22206 28142 22258
rect 28194 22206 28196 22258
rect 27244 22146 27300 22158
rect 27244 22094 27246 22146
rect 27298 22094 27300 22146
rect 26572 21746 26628 21756
rect 26684 21924 26740 21934
rect 26684 21812 26740 21868
rect 27244 21812 27300 22094
rect 27468 22148 27524 22158
rect 27692 22148 27748 22158
rect 27468 22146 27636 22148
rect 27468 22094 27470 22146
rect 27522 22094 27636 22146
rect 27468 22092 27636 22094
rect 27468 22082 27524 22092
rect 26684 21756 27300 21812
rect 27580 21812 27636 22092
rect 27692 22146 27972 22148
rect 27692 22094 27694 22146
rect 27746 22094 27972 22146
rect 27692 22092 27972 22094
rect 27692 22082 27748 22092
rect 27580 21756 27860 21812
rect 25900 20190 25902 20242
rect 25954 20190 25956 20242
rect 25900 20178 25956 20190
rect 26012 21586 26068 21598
rect 26012 21534 26014 21586
rect 26066 21534 26068 21586
rect 26012 20242 26068 21534
rect 26012 20190 26014 20242
rect 26066 20190 26068 20242
rect 26012 20178 26068 20190
rect 26684 21474 26740 21756
rect 26684 21422 26686 21474
rect 26738 21422 26740 21474
rect 25340 19966 25342 20018
rect 25394 19966 25396 20018
rect 25340 19234 25396 19966
rect 25340 19182 25342 19234
rect 25394 19182 25396 19234
rect 25340 19170 25396 19182
rect 25676 20020 25732 20030
rect 25676 19234 25732 19964
rect 25676 19182 25678 19234
rect 25730 19182 25732 19234
rect 25676 19170 25732 19182
rect 26348 20020 26404 20030
rect 26684 20020 26740 21422
rect 27020 21586 27076 21756
rect 27804 21698 27860 21756
rect 27804 21646 27806 21698
rect 27858 21646 27860 21698
rect 27804 21634 27860 21646
rect 27020 21534 27022 21586
rect 27074 21534 27076 21586
rect 27020 20914 27076 21534
rect 27916 21364 27972 22092
rect 27916 21298 27972 21308
rect 27020 20862 27022 20914
rect 27074 20862 27076 20914
rect 27020 20850 27076 20862
rect 28140 20188 28196 22206
rect 28252 22146 28308 22158
rect 28252 22094 28254 22146
rect 28306 22094 28308 22146
rect 28252 22036 28308 22094
rect 28252 21970 28308 21980
rect 29372 22036 29428 22318
rect 37660 22370 37716 22382
rect 37660 22318 37662 22370
rect 37714 22318 37716 22370
rect 29596 22148 29652 22158
rect 29596 22054 29652 22092
rect 29372 21970 29428 21980
rect 29932 22036 29988 22046
rect 29932 21474 29988 21980
rect 37660 22036 37716 22318
rect 37884 22148 37940 23102
rect 40012 22932 40068 22942
rect 40012 22838 40068 22876
rect 40012 22482 40068 22494
rect 40012 22430 40014 22482
rect 40066 22430 40068 22482
rect 40012 22260 40068 22430
rect 40012 22194 40068 22204
rect 37884 22082 37940 22092
rect 37660 21970 37716 21980
rect 37660 21588 37716 21598
rect 37660 21494 37716 21532
rect 40012 21588 40068 21598
rect 29932 21422 29934 21474
rect 29986 21422 29988 21474
rect 29932 21410 29988 21422
rect 40012 21474 40068 21532
rect 40012 21422 40014 21474
rect 40066 21422 40068 21474
rect 40012 21410 40068 21422
rect 35196 21196 35460 21206
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35196 21130 35460 21140
rect 26348 20018 26740 20020
rect 26348 19966 26350 20018
rect 26402 19966 26740 20018
rect 26348 19964 26740 19966
rect 28028 20132 28196 20188
rect 25116 19122 25172 19134
rect 25116 19070 25118 19122
rect 25170 19070 25172 19122
rect 23548 18834 23604 18844
rect 24892 19010 24948 19022
rect 24892 18958 24894 19010
rect 24946 18958 24948 19010
rect 24892 18900 24948 18958
rect 24892 18834 24948 18844
rect 25004 19010 25060 19022
rect 25004 18958 25006 19010
rect 25058 18958 25060 19010
rect 22988 18674 23212 18676
rect 22988 18622 22990 18674
rect 23042 18622 23212 18674
rect 22988 18620 23212 18622
rect 22988 18610 23044 18620
rect 23212 18610 23268 18620
rect 24108 18676 24164 18686
rect 24108 18582 24164 18620
rect 24556 18676 24612 18686
rect 24556 18582 24612 18620
rect 23884 18564 23940 18574
rect 23884 18470 23940 18508
rect 22540 18398 22542 18450
rect 22594 18398 22596 18450
rect 22540 18386 22596 18398
rect 22652 18452 22708 18462
rect 22428 15262 22430 15314
rect 22482 15262 22484 15314
rect 22428 14532 22484 15262
rect 22428 14466 22484 14476
rect 22652 18340 22708 18396
rect 23212 18452 23268 18462
rect 23212 18358 23268 18396
rect 23548 18450 23604 18462
rect 23548 18398 23550 18450
rect 23602 18398 23604 18450
rect 22764 18340 22820 18350
rect 22652 18338 22820 18340
rect 22652 18286 22766 18338
rect 22818 18286 22820 18338
rect 22652 18284 22820 18286
rect 22652 14530 22708 18284
rect 22764 18274 22820 18284
rect 23100 18338 23156 18350
rect 23100 18286 23102 18338
rect 23154 18286 23156 18338
rect 23100 17892 23156 18286
rect 23548 18340 23604 18398
rect 23548 18274 23604 18284
rect 23996 18452 24052 18462
rect 22764 17836 23156 17892
rect 22764 17778 22820 17836
rect 22764 17726 22766 17778
rect 22818 17726 22820 17778
rect 22764 17714 22820 17726
rect 23996 17106 24052 18396
rect 24444 18450 24500 18462
rect 24444 18398 24446 18450
rect 24498 18398 24500 18450
rect 24444 18340 24500 18398
rect 24444 18274 24500 18284
rect 24780 18450 24836 18462
rect 24780 18398 24782 18450
rect 24834 18398 24836 18450
rect 24220 18226 24276 18238
rect 24220 18174 24222 18226
rect 24274 18174 24276 18226
rect 23996 17054 23998 17106
rect 24050 17054 24052 17106
rect 23996 17042 24052 17054
rect 24108 17780 24164 17790
rect 24108 16994 24164 17724
rect 24108 16942 24110 16994
rect 24162 16942 24164 16994
rect 24108 16930 24164 16942
rect 24220 15540 24276 18174
rect 24780 17668 24836 18398
rect 25004 18340 25060 18958
rect 25004 18274 25060 18284
rect 24892 17780 24948 17790
rect 24892 17686 24948 17724
rect 24780 17602 24836 17612
rect 25116 17332 25172 19070
rect 25900 19124 25956 19134
rect 25900 19030 25956 19068
rect 26012 19124 26068 19134
rect 26236 19124 26292 19134
rect 26012 19122 26292 19124
rect 26012 19070 26014 19122
rect 26066 19070 26238 19122
rect 26290 19070 26292 19122
rect 26012 19068 26292 19070
rect 26012 19058 26068 19068
rect 26236 19058 26292 19068
rect 25228 18676 25284 18686
rect 25228 17554 25284 18620
rect 25340 18452 25396 18462
rect 25564 18452 25620 18462
rect 25340 18450 25564 18452
rect 25340 18398 25342 18450
rect 25394 18398 25564 18450
rect 25340 18396 25564 18398
rect 25340 18386 25396 18396
rect 25452 18228 25508 18238
rect 25452 17666 25508 18172
rect 25452 17614 25454 17666
rect 25506 17614 25508 17666
rect 25452 17602 25508 17614
rect 25228 17502 25230 17554
rect 25282 17502 25284 17554
rect 25228 17490 25284 17502
rect 25340 17442 25396 17454
rect 25340 17390 25342 17442
rect 25394 17390 25396 17442
rect 25340 17332 25396 17390
rect 25116 17276 25396 17332
rect 25340 17108 25396 17118
rect 25564 17108 25620 18396
rect 26236 18452 26292 18462
rect 26348 18452 26404 19964
rect 27020 19908 27076 19918
rect 26796 19906 27076 19908
rect 26796 19854 27022 19906
rect 27074 19854 27076 19906
rect 26796 19852 27076 19854
rect 26796 19458 26852 19852
rect 27020 19842 27076 19852
rect 26796 19406 26798 19458
rect 26850 19406 26852 19458
rect 26796 19394 26852 19406
rect 26292 18396 26404 18452
rect 26460 19010 26516 19022
rect 26460 18958 26462 19010
rect 26514 18958 26516 19010
rect 26236 18386 26292 18396
rect 26012 18340 26068 18350
rect 26012 18246 26068 18284
rect 25788 17668 25844 17678
rect 25788 17574 25844 17612
rect 26460 17668 26516 18958
rect 26684 19010 26740 19022
rect 26684 18958 26686 19010
rect 26738 18958 26740 19010
rect 26684 18788 26740 18958
rect 26684 18722 26740 18732
rect 26460 17602 26516 17612
rect 26572 18116 26628 18126
rect 26572 17666 26628 18060
rect 28028 17890 28084 20132
rect 37660 20020 37716 20030
rect 37660 19926 37716 19964
rect 29148 19908 29204 19918
rect 29148 19124 29204 19852
rect 29148 19058 29204 19068
rect 29596 19906 29652 19918
rect 29596 19854 29598 19906
rect 29650 19854 29652 19906
rect 28588 18452 28644 18462
rect 28588 18358 28644 18396
rect 29596 18452 29652 19854
rect 40012 19794 40068 19806
rect 40012 19742 40014 19794
rect 40066 19742 40068 19794
rect 35196 19628 35460 19638
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35196 19562 35460 19572
rect 40012 19572 40068 19742
rect 40012 19506 40068 19516
rect 40012 19346 40068 19358
rect 40012 19294 40014 19346
rect 40066 19294 40068 19346
rect 37884 19234 37940 19246
rect 37884 19182 37886 19234
rect 37938 19182 37940 19234
rect 29596 18386 29652 18396
rect 37660 18450 37716 18462
rect 37660 18398 37662 18450
rect 37714 18398 37716 18450
rect 28140 18338 28196 18350
rect 28140 18286 28142 18338
rect 28194 18286 28196 18338
rect 28140 18228 28196 18286
rect 28140 18162 28196 18172
rect 35196 18060 35460 18070
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35196 17994 35460 18004
rect 28028 17838 28030 17890
rect 28082 17838 28084 17890
rect 28028 17826 28084 17838
rect 37660 17892 37716 18398
rect 37884 18228 37940 19182
rect 40012 18900 40068 19294
rect 40012 18834 40068 18844
rect 37884 18162 37940 18172
rect 40012 18228 40068 18238
rect 40012 18134 40068 18172
rect 37660 17826 37716 17836
rect 40012 17778 40068 17790
rect 40012 17726 40014 17778
rect 40066 17726 40068 17778
rect 26572 17614 26574 17666
rect 26626 17614 26628 17666
rect 26572 17602 26628 17614
rect 27020 17668 27076 17678
rect 28364 17668 28420 17678
rect 27020 17666 28420 17668
rect 27020 17614 27022 17666
rect 27074 17614 28366 17666
rect 28418 17614 28420 17666
rect 27020 17612 28420 17614
rect 27020 17602 27076 17612
rect 28364 17602 28420 17612
rect 28476 17668 28532 17678
rect 28476 17574 28532 17612
rect 29484 17668 29540 17678
rect 26796 17442 26852 17454
rect 26796 17390 26798 17442
rect 26850 17390 26852 17442
rect 25396 17052 25620 17108
rect 26236 17108 26292 17118
rect 25340 17014 25396 17052
rect 26236 16884 26292 17052
rect 26572 16884 26628 16894
rect 26236 16882 26628 16884
rect 26236 16830 26574 16882
rect 26626 16830 26628 16882
rect 26236 16828 26628 16830
rect 24220 15474 24276 15484
rect 25676 15540 25732 15550
rect 25676 15446 25732 15484
rect 26124 15540 26180 15550
rect 26124 15446 26180 15484
rect 25900 15314 25956 15326
rect 25900 15262 25902 15314
rect 25954 15262 25956 15314
rect 25900 14980 25956 15262
rect 25900 14914 25956 14924
rect 26012 15202 26068 15214
rect 26012 15150 26014 15202
rect 26066 15150 26068 15202
rect 26012 14756 26068 15150
rect 26236 15148 26292 16828
rect 26572 16818 26628 16828
rect 26796 15540 26852 17390
rect 26908 17444 26964 17454
rect 27132 17444 27188 17454
rect 27916 17444 27972 17454
rect 26908 17442 27076 17444
rect 26908 17390 26910 17442
rect 26962 17390 27076 17442
rect 26908 17388 27076 17390
rect 26908 17378 26964 17388
rect 27020 17108 27076 17388
rect 27132 17442 27972 17444
rect 27132 17390 27134 17442
rect 27186 17390 27918 17442
rect 27970 17390 27972 17442
rect 27132 17388 27972 17390
rect 27132 17378 27188 17388
rect 27916 17378 27972 17388
rect 27020 17052 27412 17108
rect 27356 16994 27412 17052
rect 27356 16942 27358 16994
rect 27410 16942 27412 16994
rect 27356 16930 27412 16942
rect 29484 16770 29540 17612
rect 37660 17668 37716 17678
rect 37660 17574 37716 17612
rect 40012 17556 40068 17726
rect 40012 17490 40068 17500
rect 29484 16718 29486 16770
rect 29538 16718 29540 16770
rect 29484 16706 29540 16718
rect 35196 16492 35460 16502
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35196 16426 35460 16436
rect 26796 15474 26852 15484
rect 37660 15314 37716 15326
rect 37660 15262 37662 15314
rect 37714 15262 37716 15314
rect 26236 15092 26628 15148
rect 25676 14700 26068 14756
rect 23324 14644 23380 14654
rect 23100 14642 23380 14644
rect 23100 14590 23326 14642
rect 23378 14590 23380 14642
rect 23100 14588 23380 14590
rect 22652 14478 22654 14530
rect 22706 14478 22708 14530
rect 22540 14306 22596 14318
rect 22540 14254 22542 14306
rect 22594 14254 22596 14306
rect 22540 13858 22596 14254
rect 22652 14308 22708 14478
rect 22876 14532 22932 14542
rect 23100 14532 23156 14588
rect 23324 14578 23380 14588
rect 25004 14644 25060 14654
rect 22876 14530 23156 14532
rect 22876 14478 22878 14530
rect 22930 14478 23156 14530
rect 22876 14476 23156 14478
rect 23660 14532 23716 14542
rect 22876 14466 22932 14476
rect 23660 14438 23716 14476
rect 25004 14530 25060 14588
rect 25676 14642 25732 14700
rect 25676 14590 25678 14642
rect 25730 14590 25732 14642
rect 25676 14578 25732 14590
rect 26572 14644 26628 15092
rect 26572 14578 26628 14588
rect 26908 14980 26964 14990
rect 25004 14478 25006 14530
rect 25058 14478 25060 14530
rect 23212 14420 23268 14430
rect 23212 14326 23268 14364
rect 23548 14418 23604 14430
rect 23548 14366 23550 14418
rect 23602 14366 23604 14418
rect 22652 14242 22708 14252
rect 22540 13806 22542 13858
rect 22594 13806 22596 13858
rect 22540 13794 22596 13806
rect 21868 13746 22036 13748
rect 21868 13694 21870 13746
rect 21922 13694 22036 13746
rect 21868 13692 22036 13694
rect 21868 13524 21924 13692
rect 23548 13636 23604 14366
rect 23548 13570 23604 13580
rect 24220 13860 24276 13870
rect 21644 13468 21812 13524
rect 20636 12962 21252 12964
rect 20636 12910 20638 12962
rect 20690 12910 21252 12962
rect 20636 12908 21252 12910
rect 21420 13412 21476 13422
rect 21420 12962 21476 13356
rect 21756 13300 21812 13468
rect 21868 13458 21924 13468
rect 21756 13244 22148 13300
rect 22092 13074 22148 13244
rect 22092 13022 22094 13074
rect 22146 13022 22148 13074
rect 22092 13010 22148 13022
rect 24220 13074 24276 13804
rect 24220 13022 24222 13074
rect 24274 13022 24276 13074
rect 21420 12910 21422 12962
rect 21474 12910 21476 12962
rect 20636 12898 20692 12908
rect 21420 12898 21476 12910
rect 20524 12740 20580 12750
rect 20412 12738 20580 12740
rect 20412 12686 20526 12738
rect 20578 12686 20580 12738
rect 20412 12684 20580 12686
rect 19836 12572 20100 12582
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 19836 12506 20100 12516
rect 19836 11004 20100 11014
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 19836 10938 20100 10948
rect 19836 9436 20100 9446
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 19836 9370 20100 9380
rect 19836 7868 20100 7878
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 19836 7802 20100 7812
rect 19836 6300 20100 6310
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 19836 6234 20100 6244
rect 19836 4732 20100 4742
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 19836 4666 20100 4676
rect 20412 4338 20468 12684
rect 20524 12674 20580 12684
rect 24220 8428 24276 13022
rect 24668 13636 24724 13646
rect 24668 8428 24724 13580
rect 25004 13076 25060 14478
rect 26908 13970 26964 14924
rect 35196 14924 35460 14934
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35196 14858 35460 14868
rect 26908 13918 26910 13970
rect 26962 13918 26964 13970
rect 26908 13906 26964 13918
rect 27020 14756 27076 14766
rect 25564 13858 25620 13870
rect 25564 13806 25566 13858
rect 25618 13806 25620 13858
rect 25228 13746 25284 13758
rect 25228 13694 25230 13746
rect 25282 13694 25284 13746
rect 25228 13636 25284 13694
rect 25228 13570 25284 13580
rect 25452 13076 25508 13086
rect 25004 13074 25508 13076
rect 25004 13022 25006 13074
rect 25058 13022 25454 13074
rect 25506 13022 25508 13074
rect 25004 13020 25508 13022
rect 25004 13010 25060 13020
rect 25452 13010 25508 13020
rect 25564 8428 25620 13806
rect 27020 13858 27076 14700
rect 27804 14756 27860 14766
rect 27804 14642 27860 14700
rect 37660 14756 37716 15262
rect 40012 15202 40068 15214
rect 40012 15150 40014 15202
rect 40066 15150 40068 15202
rect 40012 14868 40068 15150
rect 40012 14802 40068 14812
rect 37660 14690 37716 14700
rect 27804 14590 27806 14642
rect 27858 14590 27860 14642
rect 27804 14578 27860 14590
rect 28252 14644 28308 14654
rect 28252 14550 28308 14588
rect 27020 13806 27022 13858
rect 27074 13806 27076 13858
rect 27020 13794 27076 13806
rect 35196 13356 35460 13366
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35196 13290 35460 13300
rect 35196 11788 35460 11798
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35196 11722 35460 11732
rect 35196 10220 35460 10230
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35196 10154 35460 10164
rect 35196 8652 35460 8662
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35196 8586 35460 8596
rect 20412 4286 20414 4338
rect 20466 4286 20468 4338
rect 20412 4274 20468 4286
rect 23548 8372 24276 8428
rect 24556 8372 24724 8428
rect 25340 8372 25620 8428
rect 19180 3490 19236 3500
rect 20188 4116 20244 4126
rect 19404 3444 19460 3454
rect 19404 3442 19572 3444
rect 19404 3390 19406 3442
rect 19458 3390 19572 3442
rect 19404 3388 19572 3390
rect 19404 3378 19460 3388
rect 19516 800 19572 3388
rect 19836 3164 20100 3174
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 19836 3098 20100 3108
rect 20188 800 20244 4060
rect 21420 4116 21476 4126
rect 21420 4022 21476 4060
rect 23548 3554 23604 8372
rect 23548 3502 23550 3554
rect 23602 3502 23604 3554
rect 23548 3490 23604 3502
rect 23772 3668 23828 3678
rect 22204 3442 22260 3454
rect 22204 3390 22206 3442
rect 22258 3390 22260 3442
rect 22204 800 22260 3390
rect 23772 980 23828 3612
rect 24556 3554 24612 8372
rect 25340 4338 25396 8372
rect 35196 7084 35460 7094
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35196 7018 35460 7028
rect 35196 5516 35460 5526
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35196 5450 35460 5460
rect 25340 4286 25342 4338
rect 25394 4286 25396 4338
rect 25340 4274 25396 4286
rect 24556 3502 24558 3554
rect 24610 3502 24612 3554
rect 24556 3490 24612 3502
rect 24892 4116 24948 4126
rect 23548 924 23828 980
rect 23548 800 23604 924
rect 24892 800 24948 4060
rect 26236 4116 26292 4126
rect 26236 4022 26292 4060
rect 35196 3948 35460 3958
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35196 3882 35460 3892
rect 25564 3668 25620 3678
rect 25564 3574 25620 3612
rect 16128 0 16240 800
rect 19488 0 19600 800
rect 20160 0 20272 800
rect 22176 0 22288 800
rect 23520 0 23632 800
rect 24864 0 24976 800
<< via2 >>
rect 4476 38442 4532 38444
rect 4476 38390 4478 38442
rect 4478 38390 4530 38442
rect 4530 38390 4532 38442
rect 4476 38388 4532 38390
rect 4580 38442 4636 38444
rect 4580 38390 4582 38442
rect 4582 38390 4634 38442
rect 4634 38390 4636 38442
rect 4580 38388 4636 38390
rect 4684 38442 4740 38444
rect 4684 38390 4686 38442
rect 4686 38390 4738 38442
rect 4738 38390 4740 38442
rect 4684 38388 4740 38390
rect 17500 38220 17556 38276
rect 18620 38274 18676 38276
rect 18620 38222 18622 38274
rect 18622 38222 18674 38274
rect 18674 38222 18676 38274
rect 18620 38220 18676 38222
rect 19516 38108 19572 38164
rect 21868 38162 21924 38164
rect 21868 38110 21870 38162
rect 21870 38110 21922 38162
rect 21922 38110 21924 38162
rect 21868 38108 21924 38110
rect 14140 37436 14196 37492
rect 4476 36874 4532 36876
rect 4476 36822 4478 36874
rect 4478 36822 4530 36874
rect 4530 36822 4532 36874
rect 4476 36820 4532 36822
rect 4580 36874 4636 36876
rect 4580 36822 4582 36874
rect 4582 36822 4634 36874
rect 4634 36822 4636 36874
rect 4580 36820 4636 36822
rect 4684 36874 4740 36876
rect 4684 36822 4686 36874
rect 4686 36822 4738 36874
rect 4738 36822 4740 36874
rect 4684 36820 4740 36822
rect 4476 35306 4532 35308
rect 4476 35254 4478 35306
rect 4478 35254 4530 35306
rect 4530 35254 4532 35306
rect 4476 35252 4532 35254
rect 4580 35306 4636 35308
rect 4580 35254 4582 35306
rect 4582 35254 4634 35306
rect 4634 35254 4636 35306
rect 4580 35252 4636 35254
rect 4684 35306 4740 35308
rect 4684 35254 4686 35306
rect 4686 35254 4738 35306
rect 4738 35254 4740 35306
rect 4684 35252 4740 35254
rect 4476 33738 4532 33740
rect 4476 33686 4478 33738
rect 4478 33686 4530 33738
rect 4530 33686 4532 33738
rect 4476 33684 4532 33686
rect 4580 33738 4636 33740
rect 4580 33686 4582 33738
rect 4582 33686 4634 33738
rect 4634 33686 4636 33738
rect 4580 33684 4636 33686
rect 4684 33738 4740 33740
rect 4684 33686 4686 33738
rect 4686 33686 4738 33738
rect 4738 33686 4740 33738
rect 4684 33684 4740 33686
rect 4476 32170 4532 32172
rect 4476 32118 4478 32170
rect 4478 32118 4530 32170
rect 4530 32118 4532 32170
rect 4476 32116 4532 32118
rect 4580 32170 4636 32172
rect 4580 32118 4582 32170
rect 4582 32118 4634 32170
rect 4634 32118 4636 32170
rect 4580 32116 4636 32118
rect 4684 32170 4740 32172
rect 4684 32118 4686 32170
rect 4686 32118 4738 32170
rect 4738 32118 4740 32170
rect 4684 32116 4740 32118
rect 4476 30602 4532 30604
rect 4476 30550 4478 30602
rect 4478 30550 4530 30602
rect 4530 30550 4532 30602
rect 4476 30548 4532 30550
rect 4580 30602 4636 30604
rect 4580 30550 4582 30602
rect 4582 30550 4634 30602
rect 4634 30550 4636 30602
rect 4580 30548 4636 30550
rect 4684 30602 4740 30604
rect 4684 30550 4686 30602
rect 4686 30550 4738 30602
rect 4738 30550 4740 30602
rect 4684 30548 4740 30550
rect 4476 29034 4532 29036
rect 4476 28982 4478 29034
rect 4478 28982 4530 29034
rect 4530 28982 4532 29034
rect 4476 28980 4532 28982
rect 4580 29034 4636 29036
rect 4580 28982 4582 29034
rect 4582 28982 4634 29034
rect 4634 28982 4636 29034
rect 4580 28980 4636 28982
rect 4684 29034 4740 29036
rect 4684 28982 4686 29034
rect 4686 28982 4738 29034
rect 4738 28982 4740 29034
rect 4684 28980 4740 28982
rect 10780 27858 10836 27860
rect 10780 27806 10782 27858
rect 10782 27806 10834 27858
rect 10834 27806 10836 27858
rect 10780 27804 10836 27806
rect 4172 27580 4228 27636
rect 1932 26236 1988 26292
rect 1932 23548 1988 23604
rect 4476 27466 4532 27468
rect 4476 27414 4478 27466
rect 4478 27414 4530 27466
rect 4530 27414 4532 27466
rect 4476 27412 4532 27414
rect 4580 27466 4636 27468
rect 4580 27414 4582 27466
rect 4582 27414 4634 27466
rect 4634 27414 4636 27466
rect 4580 27412 4636 27414
rect 4684 27466 4740 27468
rect 4684 27414 4686 27466
rect 4686 27414 4738 27466
rect 4738 27414 4740 27466
rect 4684 27412 4740 27414
rect 14028 28588 14084 28644
rect 14028 27858 14084 27860
rect 14028 27806 14030 27858
rect 14030 27806 14082 27858
rect 14082 27806 14084 27858
rect 14028 27804 14084 27806
rect 11452 27244 11508 27300
rect 13804 27132 13860 27188
rect 13916 27020 13972 27076
rect 4284 26124 4340 26180
rect 11452 26178 11508 26180
rect 11452 26126 11454 26178
rect 11454 26126 11506 26178
rect 11506 26126 11508 26178
rect 11452 26124 11508 26126
rect 4476 25898 4532 25900
rect 4476 25846 4478 25898
rect 4478 25846 4530 25898
rect 4530 25846 4532 25898
rect 4476 25844 4532 25846
rect 4580 25898 4636 25900
rect 4580 25846 4582 25898
rect 4582 25846 4634 25898
rect 4634 25846 4636 25898
rect 4580 25844 4636 25846
rect 4684 25898 4740 25900
rect 4684 25846 4686 25898
rect 4686 25846 4738 25898
rect 4738 25846 4740 25898
rect 4684 25844 4740 25846
rect 14140 26962 14196 26964
rect 14140 26910 14142 26962
rect 14142 26910 14194 26962
rect 14194 26910 14196 26962
rect 14140 26908 14196 26910
rect 15260 37490 15316 37492
rect 15260 37438 15262 37490
rect 15262 37438 15314 37490
rect 15314 37438 15316 37490
rect 15260 37436 15316 37438
rect 19628 37996 19684 38052
rect 20748 38050 20804 38052
rect 20748 37998 20750 38050
rect 20750 37998 20802 38050
rect 20802 37998 20804 38050
rect 20748 37996 20804 37998
rect 19836 37658 19892 37660
rect 19836 37606 19838 37658
rect 19838 37606 19890 37658
rect 19890 37606 19892 37658
rect 19836 37604 19892 37606
rect 19940 37658 19996 37660
rect 19940 37606 19942 37658
rect 19942 37606 19994 37658
rect 19994 37606 19996 37658
rect 19940 37604 19996 37606
rect 20044 37658 20100 37660
rect 20044 37606 20046 37658
rect 20046 37606 20098 37658
rect 20098 37606 20100 37658
rect 20044 37604 20100 37606
rect 22876 38220 22932 38276
rect 19836 36090 19892 36092
rect 19836 36038 19838 36090
rect 19838 36038 19890 36090
rect 19890 36038 19892 36090
rect 19836 36036 19892 36038
rect 19940 36090 19996 36092
rect 19940 36038 19942 36090
rect 19942 36038 19994 36090
rect 19994 36038 19996 36090
rect 19940 36036 19996 36038
rect 20044 36090 20100 36092
rect 20044 36038 20046 36090
rect 20046 36038 20098 36090
rect 20098 36038 20100 36090
rect 20044 36036 20100 36038
rect 16716 28642 16772 28644
rect 16716 28590 16718 28642
rect 16718 28590 16770 28642
rect 16770 28590 16772 28642
rect 16716 28588 16772 28590
rect 14700 27746 14756 27748
rect 14700 27694 14702 27746
rect 14702 27694 14754 27746
rect 14754 27694 14756 27746
rect 14700 27692 14756 27694
rect 15932 27692 15988 27748
rect 15148 27298 15204 27300
rect 15148 27246 15150 27298
rect 15150 27246 15202 27298
rect 15202 27246 15204 27298
rect 15148 27244 15204 27246
rect 19836 34522 19892 34524
rect 19836 34470 19838 34522
rect 19838 34470 19890 34522
rect 19890 34470 19892 34522
rect 19836 34468 19892 34470
rect 19940 34522 19996 34524
rect 19940 34470 19942 34522
rect 19942 34470 19994 34522
rect 19994 34470 19996 34522
rect 19940 34468 19996 34470
rect 20044 34522 20100 34524
rect 20044 34470 20046 34522
rect 20046 34470 20098 34522
rect 20098 34470 20100 34522
rect 20044 34468 20100 34470
rect 19836 32954 19892 32956
rect 19836 32902 19838 32954
rect 19838 32902 19890 32954
rect 19890 32902 19892 32954
rect 19836 32900 19892 32902
rect 19940 32954 19996 32956
rect 19940 32902 19942 32954
rect 19942 32902 19994 32954
rect 19994 32902 19996 32954
rect 19940 32900 19996 32902
rect 20044 32954 20100 32956
rect 20044 32902 20046 32954
rect 20046 32902 20098 32954
rect 20098 32902 20100 32954
rect 20044 32900 20100 32902
rect 19836 31386 19892 31388
rect 19836 31334 19838 31386
rect 19838 31334 19890 31386
rect 19890 31334 19892 31386
rect 19836 31332 19892 31334
rect 19940 31386 19996 31388
rect 19940 31334 19942 31386
rect 19942 31334 19994 31386
rect 19994 31334 19996 31386
rect 19940 31332 19996 31334
rect 20044 31386 20100 31388
rect 20044 31334 20046 31386
rect 20046 31334 20098 31386
rect 20098 31334 20100 31386
rect 20044 31332 20100 31334
rect 19836 29818 19892 29820
rect 19836 29766 19838 29818
rect 19838 29766 19890 29818
rect 19890 29766 19892 29818
rect 19836 29764 19892 29766
rect 19940 29818 19996 29820
rect 19940 29766 19942 29818
rect 19942 29766 19994 29818
rect 19994 29766 19996 29818
rect 19940 29764 19996 29766
rect 20044 29818 20100 29820
rect 20044 29766 20046 29818
rect 20046 29766 20098 29818
rect 20098 29766 20100 29818
rect 20044 29764 20100 29766
rect 17500 28588 17556 28644
rect 14812 27132 14868 27188
rect 14476 27020 14532 27076
rect 16044 27186 16100 27188
rect 16044 27134 16046 27186
rect 16046 27134 16098 27186
rect 16098 27134 16100 27186
rect 16044 27132 16100 27134
rect 16716 27074 16772 27076
rect 16716 27022 16718 27074
rect 16718 27022 16770 27074
rect 16770 27022 16772 27074
rect 16716 27020 16772 27022
rect 14924 26908 14980 26964
rect 16940 27186 16996 27188
rect 16940 27134 16942 27186
rect 16942 27134 16994 27186
rect 16994 27134 16996 27186
rect 16940 27132 16996 27134
rect 17164 26962 17220 26964
rect 17164 26910 17166 26962
rect 17166 26910 17218 26962
rect 17218 26910 17220 26962
rect 17164 26908 17220 26910
rect 15148 26850 15204 26852
rect 15148 26798 15150 26850
rect 15150 26798 15202 26850
rect 15202 26798 15204 26850
rect 15148 26796 15204 26798
rect 14252 26290 14308 26292
rect 14252 26238 14254 26290
rect 14254 26238 14306 26290
rect 14306 26238 14308 26290
rect 14252 26236 14308 26238
rect 13804 25506 13860 25508
rect 13804 25454 13806 25506
rect 13806 25454 13858 25506
rect 13858 25454 13860 25506
rect 13804 25452 13860 25454
rect 14812 26124 14868 26180
rect 15372 26178 15428 26180
rect 15372 26126 15374 26178
rect 15374 26126 15426 26178
rect 15426 26126 15428 26178
rect 15372 26124 15428 26126
rect 13580 25394 13636 25396
rect 13580 25342 13582 25394
rect 13582 25342 13634 25394
rect 13634 25342 13636 25394
rect 13580 25340 13636 25342
rect 13468 24892 13524 24948
rect 4476 24330 4532 24332
rect 4476 24278 4478 24330
rect 4478 24278 4530 24330
rect 4530 24278 4532 24330
rect 4476 24276 4532 24278
rect 4580 24330 4636 24332
rect 4580 24278 4582 24330
rect 4582 24278 4634 24330
rect 4634 24278 4636 24330
rect 4580 24276 4636 24278
rect 4684 24330 4740 24332
rect 4684 24278 4686 24330
rect 4686 24278 4738 24330
rect 4738 24278 4740 24330
rect 4684 24276 4740 24278
rect 4284 23938 4340 23940
rect 4284 23886 4286 23938
rect 4286 23886 4338 23938
rect 4338 23886 4340 23938
rect 4284 23884 4340 23886
rect 11004 23884 11060 23940
rect 13132 23660 13188 23716
rect 13692 23884 13748 23940
rect 14364 23826 14420 23828
rect 14364 23774 14366 23826
rect 14366 23774 14418 23826
rect 14418 23774 14420 23826
rect 14364 23772 14420 23774
rect 14700 23772 14756 23828
rect 14028 23714 14084 23716
rect 14028 23662 14030 23714
rect 14030 23662 14082 23714
rect 14082 23662 14084 23714
rect 14028 23660 14084 23662
rect 14364 23548 14420 23604
rect 4172 22876 4228 22932
rect 4476 22762 4532 22764
rect 4476 22710 4478 22762
rect 4478 22710 4530 22762
rect 4530 22710 4532 22762
rect 4476 22708 4532 22710
rect 4580 22762 4636 22764
rect 4580 22710 4582 22762
rect 4582 22710 4634 22762
rect 4634 22710 4636 22762
rect 4580 22708 4636 22710
rect 4684 22762 4740 22764
rect 4684 22710 4686 22762
rect 4686 22710 4738 22762
rect 4738 22710 4740 22762
rect 4684 22708 4740 22710
rect 14140 23100 14196 23156
rect 11340 21756 11396 21812
rect 12012 21586 12068 21588
rect 12012 21534 12014 21586
rect 12014 21534 12066 21586
rect 12066 21534 12068 21586
rect 12012 21532 12068 21534
rect 4476 21194 4532 21196
rect 4476 21142 4478 21194
rect 4478 21142 4530 21194
rect 4530 21142 4532 21194
rect 4476 21140 4532 21142
rect 4580 21194 4636 21196
rect 4580 21142 4582 21194
rect 4582 21142 4634 21194
rect 4634 21142 4636 21194
rect 4580 21140 4636 21142
rect 4684 21194 4740 21196
rect 4684 21142 4686 21194
rect 4686 21142 4738 21194
rect 4738 21142 4740 21194
rect 4684 21140 4740 21142
rect 14588 21810 14644 21812
rect 14588 21758 14590 21810
rect 14590 21758 14642 21810
rect 14642 21758 14644 21810
rect 14588 21756 14644 21758
rect 18956 26962 19012 26964
rect 18956 26910 18958 26962
rect 18958 26910 19010 26962
rect 19010 26910 19012 26962
rect 18956 26908 19012 26910
rect 18956 26290 19012 26292
rect 18956 26238 18958 26290
rect 18958 26238 19010 26290
rect 19010 26238 19012 26290
rect 18956 26236 19012 26238
rect 19964 28642 20020 28644
rect 19964 28590 19966 28642
rect 19966 28590 20018 28642
rect 20018 28590 20020 28642
rect 19964 28588 20020 28590
rect 19836 28250 19892 28252
rect 19836 28198 19838 28250
rect 19838 28198 19890 28250
rect 19890 28198 19892 28250
rect 19836 28196 19892 28198
rect 19940 28250 19996 28252
rect 19940 28198 19942 28250
rect 19942 28198 19994 28250
rect 19994 28198 19996 28250
rect 19940 28196 19996 28198
rect 20044 28250 20100 28252
rect 20044 28198 20046 28250
rect 20046 28198 20098 28250
rect 20098 28198 20100 28250
rect 20044 28196 20100 28198
rect 20188 27858 20244 27860
rect 20188 27806 20190 27858
rect 20190 27806 20242 27858
rect 20242 27806 20244 27858
rect 20188 27804 20244 27806
rect 22652 27804 22708 27860
rect 19836 26682 19892 26684
rect 19836 26630 19838 26682
rect 19838 26630 19890 26682
rect 19890 26630 19892 26682
rect 19836 26628 19892 26630
rect 19940 26682 19996 26684
rect 19940 26630 19942 26682
rect 19942 26630 19994 26682
rect 19994 26630 19996 26682
rect 19940 26628 19996 26630
rect 20044 26682 20100 26684
rect 20044 26630 20046 26682
rect 20046 26630 20098 26682
rect 20098 26630 20100 26682
rect 20044 26628 20100 26630
rect 19516 26460 19572 26516
rect 19964 26460 20020 26516
rect 19068 26348 19124 26404
rect 17388 24946 17444 24948
rect 17388 24894 17390 24946
rect 17390 24894 17442 24946
rect 17442 24894 17444 24946
rect 17388 24892 17444 24894
rect 15372 23660 15428 23716
rect 16604 23714 16660 23716
rect 16604 23662 16606 23714
rect 16606 23662 16658 23714
rect 16658 23662 16660 23714
rect 16604 23660 16660 23662
rect 15596 23266 15652 23268
rect 15596 23214 15598 23266
rect 15598 23214 15650 23266
rect 15650 23214 15652 23266
rect 15596 23212 15652 23214
rect 15372 23154 15428 23156
rect 15372 23102 15374 23154
rect 15374 23102 15426 23154
rect 15426 23102 15428 23154
rect 15372 23100 15428 23102
rect 16044 23154 16100 23156
rect 16044 23102 16046 23154
rect 16046 23102 16098 23154
rect 16098 23102 16100 23154
rect 16044 23100 16100 23102
rect 15260 22652 15316 22708
rect 14924 21698 14980 21700
rect 14924 21646 14926 21698
rect 14926 21646 14978 21698
rect 14978 21646 14980 21698
rect 14924 21644 14980 21646
rect 4476 19626 4532 19628
rect 4476 19574 4478 19626
rect 4478 19574 4530 19626
rect 4530 19574 4532 19626
rect 4476 19572 4532 19574
rect 4580 19626 4636 19628
rect 4580 19574 4582 19626
rect 4582 19574 4634 19626
rect 4634 19574 4636 19626
rect 4580 19572 4636 19574
rect 4684 19626 4740 19628
rect 4684 19574 4686 19626
rect 4686 19574 4738 19626
rect 4738 19574 4740 19626
rect 4684 19572 4740 19574
rect 14700 19404 14756 19460
rect 4476 18058 4532 18060
rect 4476 18006 4478 18058
rect 4478 18006 4530 18058
rect 4530 18006 4532 18058
rect 4476 18004 4532 18006
rect 4580 18058 4636 18060
rect 4580 18006 4582 18058
rect 4582 18006 4634 18058
rect 4634 18006 4636 18058
rect 4580 18004 4636 18006
rect 4684 18058 4740 18060
rect 4684 18006 4686 18058
rect 4686 18006 4738 18058
rect 4738 18006 4740 18058
rect 4684 18004 4740 18006
rect 12908 17724 12964 17780
rect 15372 21756 15428 21812
rect 16828 23042 16884 23044
rect 16828 22990 16830 23042
rect 16830 22990 16882 23042
rect 16882 22990 16884 23042
rect 16828 22988 16884 22990
rect 17276 22594 17332 22596
rect 17276 22542 17278 22594
rect 17278 22542 17330 22594
rect 17330 22542 17332 22594
rect 17276 22540 17332 22542
rect 15932 21810 15988 21812
rect 15932 21758 15934 21810
rect 15934 21758 15986 21810
rect 15986 21758 15988 21810
rect 15932 21756 15988 21758
rect 15708 21644 15764 21700
rect 16940 22204 16996 22260
rect 17164 21756 17220 21812
rect 16828 21644 16884 21700
rect 17612 23660 17668 23716
rect 17948 24668 18004 24724
rect 18732 26178 18788 26180
rect 18732 26126 18734 26178
rect 18734 26126 18786 26178
rect 18786 26126 18788 26178
rect 18732 26124 18788 26126
rect 18284 26066 18340 26068
rect 18284 26014 18286 26066
rect 18286 26014 18338 26066
rect 18338 26014 18340 26066
rect 18284 26012 18340 26014
rect 18732 25900 18788 25956
rect 18620 25788 18676 25844
rect 18284 25394 18340 25396
rect 18284 25342 18286 25394
rect 18286 25342 18338 25394
rect 18338 25342 18340 25394
rect 18284 25340 18340 25342
rect 18172 25228 18228 25284
rect 17500 23042 17556 23044
rect 17500 22990 17502 23042
rect 17502 22990 17554 23042
rect 17554 22990 17556 23042
rect 17500 22988 17556 22990
rect 17612 22258 17668 22260
rect 17612 22206 17614 22258
rect 17614 22206 17666 22258
rect 17666 22206 17668 22258
rect 17612 22204 17668 22206
rect 17836 23212 17892 23268
rect 18284 24834 18340 24836
rect 18284 24782 18286 24834
rect 18286 24782 18338 24834
rect 18338 24782 18340 24834
rect 18284 24780 18340 24782
rect 18396 24722 18452 24724
rect 18396 24670 18398 24722
rect 18398 24670 18450 24722
rect 18450 24670 18452 24722
rect 18396 24668 18452 24670
rect 19852 26402 19908 26404
rect 19852 26350 19854 26402
rect 19854 26350 19906 26402
rect 19906 26350 19908 26402
rect 19852 26348 19908 26350
rect 19180 26066 19236 26068
rect 19180 26014 19182 26066
rect 19182 26014 19234 26066
rect 19234 26014 19236 26066
rect 19180 26012 19236 26014
rect 19068 25788 19124 25844
rect 18732 25452 18788 25508
rect 18732 25282 18788 25284
rect 18732 25230 18734 25282
rect 18734 25230 18786 25282
rect 18786 25230 18788 25282
rect 18732 25228 18788 25230
rect 19628 26012 19684 26068
rect 19180 25506 19236 25508
rect 19180 25454 19182 25506
rect 19182 25454 19234 25506
rect 19234 25454 19236 25506
rect 19180 25452 19236 25454
rect 21756 27692 21812 27748
rect 23548 27858 23604 27860
rect 23548 27806 23550 27858
rect 23550 27806 23602 27858
rect 23602 27806 23604 27858
rect 23548 27804 23604 27806
rect 22988 27746 23044 27748
rect 22988 27694 22990 27746
rect 22990 27694 23042 27746
rect 23042 27694 23044 27746
rect 22988 27692 23044 27694
rect 35196 38442 35252 38444
rect 35196 38390 35198 38442
rect 35198 38390 35250 38442
rect 35250 38390 35252 38442
rect 35196 38388 35252 38390
rect 35300 38442 35356 38444
rect 35300 38390 35302 38442
rect 35302 38390 35354 38442
rect 35354 38390 35356 38442
rect 35300 38388 35356 38390
rect 35404 38442 35460 38444
rect 35404 38390 35406 38442
rect 35406 38390 35458 38442
rect 35458 38390 35460 38442
rect 35404 38388 35460 38390
rect 25564 38274 25620 38276
rect 25564 38222 25566 38274
rect 25566 38222 25618 38274
rect 25618 38222 25620 38274
rect 25564 38220 25620 38222
rect 24892 37436 24948 37492
rect 26236 37490 26292 37492
rect 26236 37438 26238 37490
rect 26238 37438 26290 37490
rect 26290 37438 26292 37490
rect 26236 37436 26292 37438
rect 24556 27692 24612 27748
rect 25452 27804 25508 27860
rect 20972 26796 21028 26852
rect 22540 26796 22596 26852
rect 20972 26290 21028 26292
rect 20972 26238 20974 26290
rect 20974 26238 21026 26290
rect 21026 26238 21028 26290
rect 20972 26236 21028 26238
rect 20524 26124 20580 26180
rect 21420 26348 21476 26404
rect 20524 25676 20580 25732
rect 19628 25340 19684 25396
rect 19068 25228 19124 25284
rect 19404 25282 19460 25284
rect 19404 25230 19406 25282
rect 19406 25230 19458 25282
rect 19458 25230 19460 25282
rect 19404 25228 19460 25230
rect 21084 25564 21140 25620
rect 20748 25282 20804 25284
rect 20748 25230 20750 25282
rect 20750 25230 20802 25282
rect 20802 25230 20804 25282
rect 20748 25228 20804 25230
rect 19836 25114 19892 25116
rect 19836 25062 19838 25114
rect 19838 25062 19890 25114
rect 19890 25062 19892 25114
rect 19836 25060 19892 25062
rect 19940 25114 19996 25116
rect 19940 25062 19942 25114
rect 19942 25062 19994 25114
rect 19994 25062 19996 25114
rect 19940 25060 19996 25062
rect 20044 25114 20100 25116
rect 20044 25062 20046 25114
rect 20046 25062 20098 25114
rect 20098 25062 20100 25114
rect 20044 25060 20100 25062
rect 19404 24946 19460 24948
rect 19404 24894 19406 24946
rect 19406 24894 19458 24946
rect 19458 24894 19460 24946
rect 19404 24892 19460 24894
rect 19068 24722 19124 24724
rect 19068 24670 19070 24722
rect 19070 24670 19122 24722
rect 19122 24670 19124 24722
rect 19068 24668 19124 24670
rect 17836 22258 17892 22260
rect 17836 22206 17838 22258
rect 17838 22206 17890 22258
rect 17890 22206 17892 22258
rect 17836 22204 17892 22206
rect 17724 21756 17780 21812
rect 17948 21698 18004 21700
rect 17948 21646 17950 21698
rect 17950 21646 18002 21698
rect 18002 21646 18004 21698
rect 17948 21644 18004 21646
rect 17388 21420 17444 21476
rect 18172 23826 18228 23828
rect 18172 23774 18174 23826
rect 18174 23774 18226 23826
rect 18226 23774 18228 23826
rect 18172 23772 18228 23774
rect 19836 23546 19892 23548
rect 19836 23494 19838 23546
rect 19838 23494 19890 23546
rect 19890 23494 19892 23546
rect 19836 23492 19892 23494
rect 19940 23546 19996 23548
rect 19940 23494 19942 23546
rect 19942 23494 19994 23546
rect 19994 23494 19996 23546
rect 19940 23492 19996 23494
rect 20044 23546 20100 23548
rect 20044 23494 20046 23546
rect 20046 23494 20098 23546
rect 20098 23494 20100 23546
rect 20044 23492 20100 23494
rect 20412 24722 20468 24724
rect 20412 24670 20414 24722
rect 20414 24670 20466 24722
rect 20466 24670 20468 24722
rect 20412 24668 20468 24670
rect 18732 23100 18788 23156
rect 19068 22988 19124 23044
rect 18844 22876 18900 22932
rect 19180 22876 19236 22932
rect 18284 22540 18340 22596
rect 18844 22594 18900 22596
rect 18844 22542 18846 22594
rect 18846 22542 18898 22594
rect 18898 22542 18900 22594
rect 18844 22540 18900 22542
rect 19068 22316 19124 22372
rect 18844 22204 18900 22260
rect 18172 21756 18228 21812
rect 18172 21420 18228 21476
rect 17164 19740 17220 19796
rect 14476 18172 14532 18228
rect 12908 16994 12964 16996
rect 12908 16942 12910 16994
rect 12910 16942 12962 16994
rect 12962 16942 12964 16994
rect 12908 16940 12964 16942
rect 15036 18338 15092 18340
rect 15036 18286 15038 18338
rect 15038 18286 15090 18338
rect 15090 18286 15092 18338
rect 15036 18284 15092 18286
rect 15148 17666 15204 17668
rect 15148 17614 15150 17666
rect 15150 17614 15202 17666
rect 15202 17614 15204 17666
rect 15148 17612 15204 17614
rect 14476 16940 14532 16996
rect 12236 16882 12292 16884
rect 12236 16830 12238 16882
rect 12238 16830 12290 16882
rect 12290 16830 12292 16882
rect 12236 16828 12292 16830
rect 15372 17388 15428 17444
rect 4476 16490 4532 16492
rect 4476 16438 4478 16490
rect 4478 16438 4530 16490
rect 4530 16438 4532 16490
rect 4476 16436 4532 16438
rect 4580 16490 4636 16492
rect 4580 16438 4582 16490
rect 4582 16438 4634 16490
rect 4634 16438 4636 16490
rect 4580 16436 4636 16438
rect 4684 16490 4740 16492
rect 4684 16438 4686 16490
rect 4686 16438 4738 16490
rect 4738 16438 4740 16490
rect 4684 16436 4740 16438
rect 16940 19234 16996 19236
rect 16940 19182 16942 19234
rect 16942 19182 16994 19234
rect 16994 19182 16996 19234
rect 16940 19180 16996 19182
rect 15932 19068 15988 19124
rect 18620 21420 18676 21476
rect 18396 20188 18452 20244
rect 18060 20018 18116 20020
rect 18060 19966 18062 20018
rect 18062 19966 18114 20018
rect 18114 19966 18116 20018
rect 18060 19964 18116 19966
rect 17612 19404 17668 19460
rect 16492 18396 16548 18452
rect 16268 18338 16324 18340
rect 16268 18286 16270 18338
rect 16270 18286 16322 18338
rect 16322 18286 16324 18338
rect 16268 18284 16324 18286
rect 15596 18226 15652 18228
rect 15596 18174 15598 18226
rect 15598 18174 15650 18226
rect 15650 18174 15652 18226
rect 15596 18172 15652 18174
rect 17500 18450 17556 18452
rect 17500 18398 17502 18450
rect 17502 18398 17554 18450
rect 17554 18398 17556 18450
rect 17500 18396 17556 18398
rect 15596 17666 15652 17668
rect 15596 17614 15598 17666
rect 15598 17614 15650 17666
rect 15650 17614 15652 17666
rect 15596 17612 15652 17614
rect 16716 18284 16772 18340
rect 17724 18956 17780 19012
rect 17836 18674 17892 18676
rect 17836 18622 17838 18674
rect 17838 18622 17890 18674
rect 17890 18622 17892 18674
rect 17836 18620 17892 18622
rect 17724 18396 17780 18452
rect 17052 17554 17108 17556
rect 17052 17502 17054 17554
rect 17054 17502 17106 17554
rect 17106 17502 17108 17554
rect 17052 17500 17108 17502
rect 18172 19292 18228 19348
rect 18956 20412 19012 20468
rect 19068 20076 19124 20132
rect 19628 22652 19684 22708
rect 20188 22652 20244 22708
rect 19628 21868 19684 21924
rect 19836 21978 19892 21980
rect 19836 21926 19838 21978
rect 19838 21926 19890 21978
rect 19890 21926 19892 21978
rect 19836 21924 19892 21926
rect 19940 21978 19996 21980
rect 19940 21926 19942 21978
rect 19942 21926 19994 21978
rect 19994 21926 19996 21978
rect 19940 21924 19996 21926
rect 20044 21978 20100 21980
rect 20044 21926 20046 21978
rect 20046 21926 20098 21978
rect 20098 21926 20100 21978
rect 20188 21980 20244 22036
rect 20044 21924 20100 21926
rect 19292 21644 19348 21700
rect 20188 21756 20244 21812
rect 20076 20802 20132 20804
rect 20076 20750 20078 20802
rect 20078 20750 20130 20802
rect 20130 20750 20132 20802
rect 20076 20748 20132 20750
rect 19292 19852 19348 19908
rect 19404 20412 19460 20468
rect 18620 19404 18676 19460
rect 18508 19180 18564 19236
rect 18172 18508 18228 18564
rect 18732 19068 18788 19124
rect 18620 18396 18676 18452
rect 19836 20410 19892 20412
rect 19836 20358 19838 20410
rect 19838 20358 19890 20410
rect 19890 20358 19892 20410
rect 19836 20356 19892 20358
rect 19940 20410 19996 20412
rect 19940 20358 19942 20410
rect 19942 20358 19994 20410
rect 19994 20358 19996 20410
rect 19940 20356 19996 20358
rect 20044 20410 20100 20412
rect 20044 20358 20046 20410
rect 20046 20358 20098 20410
rect 20098 20358 20100 20410
rect 20044 20356 20100 20358
rect 20300 21532 20356 21588
rect 19964 19964 20020 20020
rect 19292 18956 19348 19012
rect 19404 19068 19460 19124
rect 20076 19122 20132 19124
rect 20076 19070 20078 19122
rect 20078 19070 20130 19122
rect 20130 19070 20132 19122
rect 20076 19068 20132 19070
rect 19836 18842 19892 18844
rect 19836 18790 19838 18842
rect 19838 18790 19890 18842
rect 19890 18790 19892 18842
rect 19836 18788 19892 18790
rect 19940 18842 19996 18844
rect 19940 18790 19942 18842
rect 19942 18790 19994 18842
rect 19994 18790 19996 18842
rect 19940 18788 19996 18790
rect 20044 18842 20100 18844
rect 20044 18790 20046 18842
rect 20046 18790 20098 18842
rect 20098 18790 20100 18842
rect 20044 18788 20100 18790
rect 19180 18396 19236 18452
rect 18844 17612 18900 17668
rect 18060 17500 18116 17556
rect 18508 17554 18564 17556
rect 18508 17502 18510 17554
rect 18510 17502 18562 17554
rect 18562 17502 18564 17554
rect 18508 17500 18564 17502
rect 15484 16828 15540 16884
rect 13916 15148 13972 15204
rect 4476 14922 4532 14924
rect 4476 14870 4478 14922
rect 4478 14870 4530 14922
rect 4530 14870 4532 14922
rect 4476 14868 4532 14870
rect 4580 14922 4636 14924
rect 4580 14870 4582 14922
rect 4582 14870 4634 14922
rect 4634 14870 4636 14922
rect 4580 14868 4636 14870
rect 4684 14922 4740 14924
rect 4684 14870 4686 14922
rect 4686 14870 4738 14922
rect 4738 14870 4740 14922
rect 4684 14868 4740 14870
rect 13356 14252 13412 14308
rect 15484 14252 15540 14308
rect 16492 15372 16548 15428
rect 18956 17388 19012 17444
rect 17388 15372 17444 15428
rect 18172 15260 18228 15316
rect 18844 15314 18900 15316
rect 18844 15262 18846 15314
rect 18846 15262 18898 15314
rect 18898 15262 18900 15314
rect 18844 15260 18900 15262
rect 16268 15202 16324 15204
rect 16268 15150 16270 15202
rect 16270 15150 16322 15202
rect 16322 15150 16324 15202
rect 16268 15148 16324 15150
rect 18396 15202 18452 15204
rect 18396 15150 18398 15202
rect 18398 15150 18450 15202
rect 18450 15150 18452 15202
rect 18396 15148 18452 15150
rect 19852 18620 19908 18676
rect 20636 23436 20692 23492
rect 20524 23154 20580 23156
rect 20524 23102 20526 23154
rect 20526 23102 20578 23154
rect 20578 23102 20580 23154
rect 20524 23100 20580 23102
rect 22540 26236 22596 26292
rect 21980 25900 22036 25956
rect 21532 25788 21588 25844
rect 21756 25730 21812 25732
rect 21756 25678 21758 25730
rect 21758 25678 21810 25730
rect 21810 25678 21812 25730
rect 21756 25676 21812 25678
rect 21644 25564 21700 25620
rect 21644 25228 21700 25284
rect 21868 25282 21924 25284
rect 21868 25230 21870 25282
rect 21870 25230 21922 25282
rect 21922 25230 21924 25282
rect 21868 25228 21924 25230
rect 22316 25506 22372 25508
rect 22316 25454 22318 25506
rect 22318 25454 22370 25506
rect 22370 25454 22372 25506
rect 22316 25452 22372 25454
rect 22092 24892 22148 24948
rect 21308 23436 21364 23492
rect 21420 22930 21476 22932
rect 21420 22878 21422 22930
rect 21422 22878 21474 22930
rect 21474 22878 21476 22930
rect 21420 22876 21476 22878
rect 20748 22652 20804 22708
rect 21308 22652 21364 22708
rect 20748 22370 20804 22372
rect 20748 22318 20750 22370
rect 20750 22318 20802 22370
rect 20802 22318 20804 22370
rect 20748 22316 20804 22318
rect 20524 19964 20580 20020
rect 21420 22316 21476 22372
rect 21980 23324 22036 23380
rect 21644 22652 21700 22708
rect 21308 21756 21364 21812
rect 21868 21868 21924 21924
rect 23772 26514 23828 26516
rect 23772 26462 23774 26514
rect 23774 26462 23826 26514
rect 23826 26462 23828 26514
rect 23772 26460 23828 26462
rect 23212 26290 23268 26292
rect 23212 26238 23214 26290
rect 23214 26238 23266 26290
rect 23266 26238 23268 26290
rect 23212 26236 23268 26238
rect 35196 36874 35252 36876
rect 35196 36822 35198 36874
rect 35198 36822 35250 36874
rect 35250 36822 35252 36874
rect 35196 36820 35252 36822
rect 35300 36874 35356 36876
rect 35300 36822 35302 36874
rect 35302 36822 35354 36874
rect 35354 36822 35356 36874
rect 35300 36820 35356 36822
rect 35404 36874 35460 36876
rect 35404 36822 35406 36874
rect 35406 36822 35458 36874
rect 35458 36822 35460 36874
rect 35404 36820 35460 36822
rect 35196 35306 35252 35308
rect 35196 35254 35198 35306
rect 35198 35254 35250 35306
rect 35250 35254 35252 35306
rect 35196 35252 35252 35254
rect 35300 35306 35356 35308
rect 35300 35254 35302 35306
rect 35302 35254 35354 35306
rect 35354 35254 35356 35306
rect 35300 35252 35356 35254
rect 35404 35306 35460 35308
rect 35404 35254 35406 35306
rect 35406 35254 35458 35306
rect 35458 35254 35460 35306
rect 35404 35252 35460 35254
rect 35196 33738 35252 33740
rect 35196 33686 35198 33738
rect 35198 33686 35250 33738
rect 35250 33686 35252 33738
rect 35196 33684 35252 33686
rect 35300 33738 35356 33740
rect 35300 33686 35302 33738
rect 35302 33686 35354 33738
rect 35354 33686 35356 33738
rect 35300 33684 35356 33686
rect 35404 33738 35460 33740
rect 35404 33686 35406 33738
rect 35406 33686 35458 33738
rect 35458 33686 35460 33738
rect 35404 33684 35460 33686
rect 35196 32170 35252 32172
rect 35196 32118 35198 32170
rect 35198 32118 35250 32170
rect 35250 32118 35252 32170
rect 35196 32116 35252 32118
rect 35300 32170 35356 32172
rect 35300 32118 35302 32170
rect 35302 32118 35354 32170
rect 35354 32118 35356 32170
rect 35300 32116 35356 32118
rect 35404 32170 35460 32172
rect 35404 32118 35406 32170
rect 35406 32118 35458 32170
rect 35458 32118 35460 32170
rect 35404 32116 35460 32118
rect 35196 30602 35252 30604
rect 35196 30550 35198 30602
rect 35198 30550 35250 30602
rect 35250 30550 35252 30602
rect 35196 30548 35252 30550
rect 35300 30602 35356 30604
rect 35300 30550 35302 30602
rect 35302 30550 35354 30602
rect 35354 30550 35356 30602
rect 35300 30548 35356 30550
rect 35404 30602 35460 30604
rect 35404 30550 35406 30602
rect 35406 30550 35458 30602
rect 35458 30550 35460 30602
rect 35404 30548 35460 30550
rect 35196 29034 35252 29036
rect 35196 28982 35198 29034
rect 35198 28982 35250 29034
rect 35250 28982 35252 29034
rect 35196 28980 35252 28982
rect 35300 29034 35356 29036
rect 35300 28982 35302 29034
rect 35302 28982 35354 29034
rect 35354 28982 35356 29034
rect 35300 28980 35356 28982
rect 35404 29034 35460 29036
rect 35404 28982 35406 29034
rect 35406 28982 35458 29034
rect 35458 28982 35460 29034
rect 35404 28980 35460 28982
rect 26012 27804 26068 27860
rect 35196 27466 35252 27468
rect 35196 27414 35198 27466
rect 35198 27414 35250 27466
rect 35250 27414 35252 27466
rect 35196 27412 35252 27414
rect 35300 27466 35356 27468
rect 35300 27414 35302 27466
rect 35302 27414 35354 27466
rect 35354 27414 35356 27466
rect 35300 27412 35356 27414
rect 35404 27466 35460 27468
rect 35404 27414 35406 27466
rect 35406 27414 35458 27466
rect 35458 27414 35460 27466
rect 35404 27412 35460 27414
rect 27580 27020 27636 27076
rect 25564 26460 25620 26516
rect 26348 26796 26404 26852
rect 23548 25564 23604 25620
rect 25676 26124 25732 26180
rect 22764 25228 22820 25284
rect 23436 25452 23492 25508
rect 22316 22540 22372 22596
rect 22316 21980 22372 22036
rect 21532 20578 21588 20580
rect 21532 20526 21534 20578
rect 21534 20526 21586 20578
rect 21586 20526 21588 20578
rect 21532 20524 21588 20526
rect 20972 20018 21028 20020
rect 20972 19966 20974 20018
rect 20974 19966 21026 20018
rect 21026 19966 21028 20018
rect 20972 19964 21028 19966
rect 21756 20130 21812 20132
rect 21756 20078 21758 20130
rect 21758 20078 21810 20130
rect 21810 20078 21812 20130
rect 21756 20076 21812 20078
rect 21420 19964 21476 20020
rect 22092 19964 22148 20020
rect 21308 19852 21364 19908
rect 20636 19794 20692 19796
rect 20636 19742 20638 19794
rect 20638 19742 20690 19794
rect 20690 19742 20692 19794
rect 20636 19740 20692 19742
rect 21196 19740 21252 19796
rect 20300 18620 20356 18676
rect 20748 18732 20804 18788
rect 20076 18396 20132 18452
rect 19404 18284 19460 18340
rect 19628 18172 19684 18228
rect 19404 17666 19460 17668
rect 19404 17614 19406 17666
rect 19406 17614 19458 17666
rect 19458 17614 19460 17666
rect 19404 17612 19460 17614
rect 20860 18396 20916 18452
rect 22316 21756 22372 21812
rect 22316 20524 22372 20580
rect 22540 22370 22596 22372
rect 22540 22318 22542 22370
rect 22542 22318 22594 22370
rect 22594 22318 22596 22370
rect 22540 22316 22596 22318
rect 22988 21532 23044 21588
rect 21756 18844 21812 18900
rect 20188 18226 20244 18228
rect 20188 18174 20190 18226
rect 20190 18174 20242 18226
rect 20242 18174 20244 18226
rect 20188 18172 20244 18174
rect 21420 18226 21476 18228
rect 21420 18174 21422 18226
rect 21422 18174 21474 18226
rect 21474 18174 21476 18226
rect 21420 18172 21476 18174
rect 22876 20802 22932 20804
rect 22876 20750 22878 20802
rect 22878 20750 22930 20802
rect 22930 20750 22932 20802
rect 22876 20748 22932 20750
rect 22428 19122 22484 19124
rect 22428 19070 22430 19122
rect 22430 19070 22482 19122
rect 22482 19070 22484 19122
rect 22428 19068 22484 19070
rect 22204 18732 22260 18788
rect 22092 18620 22148 18676
rect 21980 18284 22036 18340
rect 21756 18060 21812 18116
rect 20300 17724 20356 17780
rect 19836 17274 19892 17276
rect 19836 17222 19838 17274
rect 19838 17222 19890 17274
rect 19890 17222 19892 17274
rect 19836 17220 19892 17222
rect 19940 17274 19996 17276
rect 19940 17222 19942 17274
rect 19942 17222 19994 17274
rect 19994 17222 19996 17274
rect 19940 17220 19996 17222
rect 20044 17274 20100 17276
rect 20044 17222 20046 17274
rect 20046 17222 20098 17274
rect 20098 17222 20100 17274
rect 20044 17220 20100 17222
rect 21980 17052 22036 17108
rect 19836 15706 19892 15708
rect 19836 15654 19838 15706
rect 19838 15654 19890 15706
rect 19890 15654 19892 15706
rect 19836 15652 19892 15654
rect 19940 15706 19996 15708
rect 19940 15654 19942 15706
rect 19942 15654 19994 15706
rect 19994 15654 19996 15706
rect 19940 15652 19996 15654
rect 20044 15706 20100 15708
rect 20044 15654 20046 15706
rect 20046 15654 20098 15706
rect 20098 15654 20100 15706
rect 20044 15652 20100 15654
rect 21868 15426 21924 15428
rect 21868 15374 21870 15426
rect 21870 15374 21922 15426
rect 21922 15374 21924 15426
rect 21868 15372 21924 15374
rect 19964 15148 20020 15204
rect 18284 14476 18340 14532
rect 16268 14252 16324 14308
rect 4476 13354 4532 13356
rect 4476 13302 4478 13354
rect 4478 13302 4530 13354
rect 4530 13302 4532 13354
rect 4476 13300 4532 13302
rect 4580 13354 4636 13356
rect 4580 13302 4582 13354
rect 4582 13302 4634 13354
rect 4634 13302 4636 13354
rect 4580 13300 4636 13302
rect 4684 13354 4740 13356
rect 4684 13302 4686 13354
rect 4686 13302 4738 13354
rect 4738 13302 4740 13354
rect 4684 13300 4740 13302
rect 16828 14252 16884 14308
rect 17612 14252 17668 14308
rect 16044 12460 16100 12516
rect 17388 12460 17444 12516
rect 4476 11786 4532 11788
rect 4476 11734 4478 11786
rect 4478 11734 4530 11786
rect 4530 11734 4532 11786
rect 4476 11732 4532 11734
rect 4580 11786 4636 11788
rect 4580 11734 4582 11786
rect 4582 11734 4634 11786
rect 4634 11734 4636 11786
rect 4580 11732 4636 11734
rect 4684 11786 4740 11788
rect 4684 11734 4686 11786
rect 4686 11734 4738 11786
rect 4738 11734 4740 11786
rect 4684 11732 4740 11734
rect 4476 10218 4532 10220
rect 4476 10166 4478 10218
rect 4478 10166 4530 10218
rect 4530 10166 4532 10218
rect 4476 10164 4532 10166
rect 4580 10218 4636 10220
rect 4580 10166 4582 10218
rect 4582 10166 4634 10218
rect 4634 10166 4636 10218
rect 4580 10164 4636 10166
rect 4684 10218 4740 10220
rect 4684 10166 4686 10218
rect 4686 10166 4738 10218
rect 4738 10166 4740 10218
rect 4684 10164 4740 10166
rect 4476 8650 4532 8652
rect 4476 8598 4478 8650
rect 4478 8598 4530 8650
rect 4530 8598 4532 8650
rect 4476 8596 4532 8598
rect 4580 8650 4636 8652
rect 4580 8598 4582 8650
rect 4582 8598 4634 8650
rect 4634 8598 4636 8650
rect 4580 8596 4636 8598
rect 4684 8650 4740 8652
rect 4684 8598 4686 8650
rect 4686 8598 4738 8650
rect 4738 8598 4740 8650
rect 4684 8596 4740 8598
rect 4476 7082 4532 7084
rect 4476 7030 4478 7082
rect 4478 7030 4530 7082
rect 4530 7030 4532 7082
rect 4476 7028 4532 7030
rect 4580 7082 4636 7084
rect 4580 7030 4582 7082
rect 4582 7030 4634 7082
rect 4634 7030 4636 7082
rect 4580 7028 4636 7030
rect 4684 7082 4740 7084
rect 4684 7030 4686 7082
rect 4686 7030 4738 7082
rect 4738 7030 4740 7082
rect 4684 7028 4740 7030
rect 4476 5514 4532 5516
rect 4476 5462 4478 5514
rect 4478 5462 4530 5514
rect 4530 5462 4532 5514
rect 4476 5460 4532 5462
rect 4580 5514 4636 5516
rect 4580 5462 4582 5514
rect 4582 5462 4634 5514
rect 4634 5462 4636 5514
rect 4580 5460 4636 5462
rect 4684 5514 4740 5516
rect 4684 5462 4686 5514
rect 4686 5462 4738 5514
rect 4738 5462 4740 5514
rect 4684 5460 4740 5462
rect 16156 4172 16212 4228
rect 4476 3946 4532 3948
rect 4476 3894 4478 3946
rect 4478 3894 4530 3946
rect 4530 3894 4532 3946
rect 4476 3892 4532 3894
rect 4580 3946 4636 3948
rect 4580 3894 4582 3946
rect 4582 3894 4634 3946
rect 4634 3894 4636 3946
rect 4580 3892 4636 3894
rect 4684 3946 4740 3948
rect 4684 3894 4686 3946
rect 4686 3894 4738 3946
rect 4738 3894 4740 3946
rect 4684 3892 4740 3894
rect 18508 4226 18564 4228
rect 18508 4174 18510 4226
rect 18510 4174 18562 4226
rect 18562 4174 18564 4226
rect 18508 4172 18564 4174
rect 18060 3554 18116 3556
rect 18060 3502 18062 3554
rect 18062 3502 18114 3554
rect 18114 3502 18116 3554
rect 18060 3500 18116 3502
rect 19852 14530 19908 14532
rect 19852 14478 19854 14530
rect 19854 14478 19906 14530
rect 19906 14478 19908 14530
rect 19852 14476 19908 14478
rect 20188 14530 20244 14532
rect 20188 14478 20190 14530
rect 20190 14478 20242 14530
rect 20242 14478 20244 14530
rect 20188 14476 20244 14478
rect 21868 14530 21924 14532
rect 21868 14478 21870 14530
rect 21870 14478 21922 14530
rect 21922 14478 21924 14530
rect 21868 14476 21924 14478
rect 19964 14418 20020 14420
rect 19964 14366 19966 14418
rect 19966 14366 20018 14418
rect 20018 14366 20020 14418
rect 19964 14364 20020 14366
rect 21420 14364 21476 14420
rect 20636 14306 20692 14308
rect 20636 14254 20638 14306
rect 20638 14254 20690 14306
rect 20690 14254 20692 14306
rect 20636 14252 20692 14254
rect 19836 14138 19892 14140
rect 19836 14086 19838 14138
rect 19838 14086 19890 14138
rect 19890 14086 19892 14138
rect 19836 14084 19892 14086
rect 19940 14138 19996 14140
rect 19940 14086 19942 14138
rect 19942 14086 19994 14138
rect 19994 14086 19996 14138
rect 19940 14084 19996 14086
rect 20044 14138 20100 14140
rect 20044 14086 20046 14138
rect 20046 14086 20098 14138
rect 20098 14086 20100 14138
rect 20044 14084 20100 14086
rect 21308 13858 21364 13860
rect 21308 13806 21310 13858
rect 21310 13806 21362 13858
rect 21362 13806 21364 13858
rect 21308 13804 21364 13806
rect 19628 13132 19684 13188
rect 20524 13186 20580 13188
rect 20524 13134 20526 13186
rect 20526 13134 20578 13186
rect 20578 13134 20580 13186
rect 20524 13132 20580 13134
rect 21756 14306 21812 14308
rect 21756 14254 21758 14306
rect 21758 14254 21810 14306
rect 21810 14254 21812 14306
rect 21756 14252 21812 14254
rect 22204 14530 22260 14532
rect 22204 14478 22206 14530
rect 22206 14478 22258 14530
rect 22258 14478 22260 14530
rect 22204 14476 22260 14478
rect 24668 23042 24724 23044
rect 24668 22990 24670 23042
rect 24670 22990 24722 23042
rect 24722 22990 24724 23042
rect 24668 22988 24724 22990
rect 23996 21868 24052 21924
rect 26236 24946 26292 24948
rect 26236 24894 26238 24946
rect 26238 24894 26290 24946
rect 26290 24894 26292 24946
rect 26236 24892 26292 24894
rect 28364 27020 28420 27076
rect 27356 26850 27412 26852
rect 27356 26798 27358 26850
rect 27358 26798 27410 26850
rect 27410 26798 27412 26850
rect 27356 26796 27412 26798
rect 27020 25452 27076 25508
rect 37660 27074 37716 27076
rect 37660 27022 37662 27074
rect 37662 27022 37714 27074
rect 37714 27022 37716 27074
rect 37660 27020 37716 27022
rect 28812 26178 28868 26180
rect 28812 26126 28814 26178
rect 28814 26126 28866 26178
rect 28866 26126 28868 26178
rect 28812 26124 28868 26126
rect 27804 25564 27860 25620
rect 28588 25618 28644 25620
rect 28588 25566 28590 25618
rect 28590 25566 28642 25618
rect 28642 25566 28644 25618
rect 28588 25564 28644 25566
rect 35196 25898 35252 25900
rect 35196 25846 35198 25898
rect 35198 25846 35250 25898
rect 35250 25846 35252 25898
rect 35196 25844 35252 25846
rect 35300 25898 35356 25900
rect 35300 25846 35302 25898
rect 35302 25846 35354 25898
rect 35354 25846 35356 25898
rect 35300 25844 35356 25846
rect 35404 25898 35460 25900
rect 35404 25846 35406 25898
rect 35406 25846 35458 25898
rect 35458 25846 35460 25898
rect 35404 25844 35460 25846
rect 40012 26236 40068 26292
rect 37660 25564 37716 25620
rect 40012 25564 40068 25620
rect 26124 23714 26180 23716
rect 26124 23662 26126 23714
rect 26126 23662 26178 23714
rect 26178 23662 26180 23714
rect 26124 23660 26180 23662
rect 26460 23714 26516 23716
rect 26460 23662 26462 23714
rect 26462 23662 26514 23714
rect 26514 23662 26516 23714
rect 26460 23660 26516 23662
rect 35196 24330 35252 24332
rect 35196 24278 35198 24330
rect 35198 24278 35250 24330
rect 35250 24278 35252 24330
rect 35196 24276 35252 24278
rect 35300 24330 35356 24332
rect 35300 24278 35302 24330
rect 35302 24278 35354 24330
rect 35354 24278 35356 24330
rect 35300 24276 35356 24278
rect 35404 24330 35460 24332
rect 35404 24278 35406 24330
rect 35406 24278 35458 24330
rect 35458 24278 35460 24330
rect 35404 24276 35460 24278
rect 27916 23660 27972 23716
rect 28364 23660 28420 23716
rect 24556 21756 24612 21812
rect 25340 21868 25396 21924
rect 25452 21980 25508 22036
rect 25900 21756 25956 21812
rect 24668 21644 24724 21700
rect 25340 21698 25396 21700
rect 25340 21646 25342 21698
rect 25342 21646 25394 21698
rect 25394 21646 25396 21698
rect 25340 21644 25396 21646
rect 25564 21532 25620 21588
rect 25228 21420 25284 21476
rect 25340 21308 25396 21364
rect 25340 20188 25396 20244
rect 23660 20130 23716 20132
rect 23660 20078 23662 20130
rect 23662 20078 23714 20130
rect 23714 20078 23716 20130
rect 23660 20076 23716 20078
rect 23772 20018 23828 20020
rect 23772 19966 23774 20018
rect 23774 19966 23826 20018
rect 23826 19966 23828 20018
rect 23772 19964 23828 19966
rect 40012 23548 40068 23604
rect 37324 22988 37380 23044
rect 35196 22762 35252 22764
rect 35196 22710 35198 22762
rect 35198 22710 35250 22762
rect 35250 22710 35252 22762
rect 35196 22708 35252 22710
rect 35300 22762 35356 22764
rect 35300 22710 35302 22762
rect 35302 22710 35354 22762
rect 35354 22710 35356 22762
rect 35300 22708 35356 22710
rect 35404 22762 35460 22764
rect 35404 22710 35406 22762
rect 35406 22710 35458 22762
rect 35458 22710 35460 22762
rect 35404 22708 35460 22710
rect 26572 21756 26628 21812
rect 26684 21868 26740 21924
rect 25676 20018 25732 20020
rect 25676 19966 25678 20018
rect 25678 19966 25730 20018
rect 25730 19966 25732 20018
rect 25676 19964 25732 19966
rect 27916 21308 27972 21364
rect 28252 21980 28308 22036
rect 29596 22146 29652 22148
rect 29596 22094 29598 22146
rect 29598 22094 29650 22146
rect 29650 22094 29652 22146
rect 29596 22092 29652 22094
rect 29372 21980 29428 22036
rect 29932 21980 29988 22036
rect 40012 22930 40068 22932
rect 40012 22878 40014 22930
rect 40014 22878 40066 22930
rect 40066 22878 40068 22930
rect 40012 22876 40068 22878
rect 40012 22204 40068 22260
rect 37884 22092 37940 22148
rect 37660 21980 37716 22036
rect 37660 21586 37716 21588
rect 37660 21534 37662 21586
rect 37662 21534 37714 21586
rect 37714 21534 37716 21586
rect 37660 21532 37716 21534
rect 40012 21532 40068 21588
rect 35196 21194 35252 21196
rect 35196 21142 35198 21194
rect 35198 21142 35250 21194
rect 35250 21142 35252 21194
rect 35196 21140 35252 21142
rect 35300 21194 35356 21196
rect 35300 21142 35302 21194
rect 35302 21142 35354 21194
rect 35354 21142 35356 21194
rect 35300 21140 35356 21142
rect 35404 21194 35460 21196
rect 35404 21142 35406 21194
rect 35406 21142 35458 21194
rect 35458 21142 35460 21194
rect 35404 21140 35460 21142
rect 23548 18844 23604 18900
rect 24892 18844 24948 18900
rect 23212 18620 23268 18676
rect 24108 18674 24164 18676
rect 24108 18622 24110 18674
rect 24110 18622 24162 18674
rect 24162 18622 24164 18674
rect 24108 18620 24164 18622
rect 24556 18674 24612 18676
rect 24556 18622 24558 18674
rect 24558 18622 24610 18674
rect 24610 18622 24612 18674
rect 24556 18620 24612 18622
rect 23884 18562 23940 18564
rect 23884 18510 23886 18562
rect 23886 18510 23938 18562
rect 23938 18510 23940 18562
rect 23884 18508 23940 18510
rect 22652 18396 22708 18452
rect 22428 14476 22484 14532
rect 23212 18450 23268 18452
rect 23212 18398 23214 18450
rect 23214 18398 23266 18450
rect 23266 18398 23268 18450
rect 23212 18396 23268 18398
rect 23548 18284 23604 18340
rect 23996 18396 24052 18452
rect 24444 18284 24500 18340
rect 24108 17724 24164 17780
rect 25004 18284 25060 18340
rect 24892 17778 24948 17780
rect 24892 17726 24894 17778
rect 24894 17726 24946 17778
rect 24946 17726 24948 17778
rect 24892 17724 24948 17726
rect 24780 17612 24836 17668
rect 25900 19122 25956 19124
rect 25900 19070 25902 19122
rect 25902 19070 25954 19122
rect 25954 19070 25956 19122
rect 25900 19068 25956 19070
rect 25228 18620 25284 18676
rect 25564 18396 25620 18452
rect 25452 18172 25508 18228
rect 26236 18396 26292 18452
rect 26012 18338 26068 18340
rect 26012 18286 26014 18338
rect 26014 18286 26066 18338
rect 26066 18286 26068 18338
rect 26012 18284 26068 18286
rect 25788 17666 25844 17668
rect 25788 17614 25790 17666
rect 25790 17614 25842 17666
rect 25842 17614 25844 17666
rect 25788 17612 25844 17614
rect 26684 18732 26740 18788
rect 26460 17612 26516 17668
rect 26572 18060 26628 18116
rect 37660 20018 37716 20020
rect 37660 19966 37662 20018
rect 37662 19966 37714 20018
rect 37714 19966 37716 20018
rect 37660 19964 37716 19966
rect 29148 19906 29204 19908
rect 29148 19854 29150 19906
rect 29150 19854 29202 19906
rect 29202 19854 29204 19906
rect 29148 19852 29204 19854
rect 29148 19068 29204 19124
rect 28588 18450 28644 18452
rect 28588 18398 28590 18450
rect 28590 18398 28642 18450
rect 28642 18398 28644 18450
rect 28588 18396 28644 18398
rect 35196 19626 35252 19628
rect 35196 19574 35198 19626
rect 35198 19574 35250 19626
rect 35250 19574 35252 19626
rect 35196 19572 35252 19574
rect 35300 19626 35356 19628
rect 35300 19574 35302 19626
rect 35302 19574 35354 19626
rect 35354 19574 35356 19626
rect 35300 19572 35356 19574
rect 35404 19626 35460 19628
rect 35404 19574 35406 19626
rect 35406 19574 35458 19626
rect 35458 19574 35460 19626
rect 35404 19572 35460 19574
rect 40012 19516 40068 19572
rect 29596 18396 29652 18452
rect 28140 18172 28196 18228
rect 35196 18058 35252 18060
rect 35196 18006 35198 18058
rect 35198 18006 35250 18058
rect 35250 18006 35252 18058
rect 35196 18004 35252 18006
rect 35300 18058 35356 18060
rect 35300 18006 35302 18058
rect 35302 18006 35354 18058
rect 35354 18006 35356 18058
rect 35300 18004 35356 18006
rect 35404 18058 35460 18060
rect 35404 18006 35406 18058
rect 35406 18006 35458 18058
rect 35458 18006 35460 18058
rect 35404 18004 35460 18006
rect 40012 18844 40068 18900
rect 37884 18172 37940 18228
rect 40012 18226 40068 18228
rect 40012 18174 40014 18226
rect 40014 18174 40066 18226
rect 40066 18174 40068 18226
rect 40012 18172 40068 18174
rect 37660 17836 37716 17892
rect 28476 17666 28532 17668
rect 28476 17614 28478 17666
rect 28478 17614 28530 17666
rect 28530 17614 28532 17666
rect 28476 17612 28532 17614
rect 29484 17612 29540 17668
rect 25340 17106 25396 17108
rect 25340 17054 25342 17106
rect 25342 17054 25394 17106
rect 25394 17054 25396 17106
rect 25340 17052 25396 17054
rect 26236 17106 26292 17108
rect 26236 17054 26238 17106
rect 26238 17054 26290 17106
rect 26290 17054 26292 17106
rect 26236 17052 26292 17054
rect 24220 15484 24276 15540
rect 25676 15538 25732 15540
rect 25676 15486 25678 15538
rect 25678 15486 25730 15538
rect 25730 15486 25732 15538
rect 25676 15484 25732 15486
rect 26124 15538 26180 15540
rect 26124 15486 26126 15538
rect 26126 15486 26178 15538
rect 26178 15486 26180 15538
rect 26124 15484 26180 15486
rect 25900 14924 25956 14980
rect 37660 17666 37716 17668
rect 37660 17614 37662 17666
rect 37662 17614 37714 17666
rect 37714 17614 37716 17666
rect 37660 17612 37716 17614
rect 40012 17500 40068 17556
rect 35196 16490 35252 16492
rect 35196 16438 35198 16490
rect 35198 16438 35250 16490
rect 35250 16438 35252 16490
rect 35196 16436 35252 16438
rect 35300 16490 35356 16492
rect 35300 16438 35302 16490
rect 35302 16438 35354 16490
rect 35354 16438 35356 16490
rect 35300 16436 35356 16438
rect 35404 16490 35460 16492
rect 35404 16438 35406 16490
rect 35406 16438 35458 16490
rect 35458 16438 35460 16490
rect 35404 16436 35460 16438
rect 26796 15484 26852 15540
rect 25004 14588 25060 14644
rect 23660 14530 23716 14532
rect 23660 14478 23662 14530
rect 23662 14478 23714 14530
rect 23714 14478 23716 14530
rect 23660 14476 23716 14478
rect 26572 14588 26628 14644
rect 26908 14924 26964 14980
rect 23212 14418 23268 14420
rect 23212 14366 23214 14418
rect 23214 14366 23266 14418
rect 23266 14366 23268 14418
rect 23212 14364 23268 14366
rect 22652 14252 22708 14308
rect 23548 13580 23604 13636
rect 24220 13804 24276 13860
rect 21420 13356 21476 13412
rect 21868 13468 21924 13524
rect 19836 12570 19892 12572
rect 19836 12518 19838 12570
rect 19838 12518 19890 12570
rect 19890 12518 19892 12570
rect 19836 12516 19892 12518
rect 19940 12570 19996 12572
rect 19940 12518 19942 12570
rect 19942 12518 19994 12570
rect 19994 12518 19996 12570
rect 19940 12516 19996 12518
rect 20044 12570 20100 12572
rect 20044 12518 20046 12570
rect 20046 12518 20098 12570
rect 20098 12518 20100 12570
rect 20044 12516 20100 12518
rect 19836 11002 19892 11004
rect 19836 10950 19838 11002
rect 19838 10950 19890 11002
rect 19890 10950 19892 11002
rect 19836 10948 19892 10950
rect 19940 11002 19996 11004
rect 19940 10950 19942 11002
rect 19942 10950 19994 11002
rect 19994 10950 19996 11002
rect 19940 10948 19996 10950
rect 20044 11002 20100 11004
rect 20044 10950 20046 11002
rect 20046 10950 20098 11002
rect 20098 10950 20100 11002
rect 20044 10948 20100 10950
rect 19836 9434 19892 9436
rect 19836 9382 19838 9434
rect 19838 9382 19890 9434
rect 19890 9382 19892 9434
rect 19836 9380 19892 9382
rect 19940 9434 19996 9436
rect 19940 9382 19942 9434
rect 19942 9382 19994 9434
rect 19994 9382 19996 9434
rect 19940 9380 19996 9382
rect 20044 9434 20100 9436
rect 20044 9382 20046 9434
rect 20046 9382 20098 9434
rect 20098 9382 20100 9434
rect 20044 9380 20100 9382
rect 19836 7866 19892 7868
rect 19836 7814 19838 7866
rect 19838 7814 19890 7866
rect 19890 7814 19892 7866
rect 19836 7812 19892 7814
rect 19940 7866 19996 7868
rect 19940 7814 19942 7866
rect 19942 7814 19994 7866
rect 19994 7814 19996 7866
rect 19940 7812 19996 7814
rect 20044 7866 20100 7868
rect 20044 7814 20046 7866
rect 20046 7814 20098 7866
rect 20098 7814 20100 7866
rect 20044 7812 20100 7814
rect 19836 6298 19892 6300
rect 19836 6246 19838 6298
rect 19838 6246 19890 6298
rect 19890 6246 19892 6298
rect 19836 6244 19892 6246
rect 19940 6298 19996 6300
rect 19940 6246 19942 6298
rect 19942 6246 19994 6298
rect 19994 6246 19996 6298
rect 19940 6244 19996 6246
rect 20044 6298 20100 6300
rect 20044 6246 20046 6298
rect 20046 6246 20098 6298
rect 20098 6246 20100 6298
rect 20044 6244 20100 6246
rect 19836 4730 19892 4732
rect 19836 4678 19838 4730
rect 19838 4678 19890 4730
rect 19890 4678 19892 4730
rect 19836 4676 19892 4678
rect 19940 4730 19996 4732
rect 19940 4678 19942 4730
rect 19942 4678 19994 4730
rect 19994 4678 19996 4730
rect 19940 4676 19996 4678
rect 20044 4730 20100 4732
rect 20044 4678 20046 4730
rect 20046 4678 20098 4730
rect 20098 4678 20100 4730
rect 20044 4676 20100 4678
rect 24668 13634 24724 13636
rect 24668 13582 24670 13634
rect 24670 13582 24722 13634
rect 24722 13582 24724 13634
rect 24668 13580 24724 13582
rect 35196 14922 35252 14924
rect 35196 14870 35198 14922
rect 35198 14870 35250 14922
rect 35250 14870 35252 14922
rect 35196 14868 35252 14870
rect 35300 14922 35356 14924
rect 35300 14870 35302 14922
rect 35302 14870 35354 14922
rect 35354 14870 35356 14922
rect 35300 14868 35356 14870
rect 35404 14922 35460 14924
rect 35404 14870 35406 14922
rect 35406 14870 35458 14922
rect 35458 14870 35460 14922
rect 35404 14868 35460 14870
rect 27020 14700 27076 14756
rect 25228 13580 25284 13636
rect 27804 14700 27860 14756
rect 40012 14812 40068 14868
rect 37660 14700 37716 14756
rect 28252 14642 28308 14644
rect 28252 14590 28254 14642
rect 28254 14590 28306 14642
rect 28306 14590 28308 14642
rect 28252 14588 28308 14590
rect 35196 13354 35252 13356
rect 35196 13302 35198 13354
rect 35198 13302 35250 13354
rect 35250 13302 35252 13354
rect 35196 13300 35252 13302
rect 35300 13354 35356 13356
rect 35300 13302 35302 13354
rect 35302 13302 35354 13354
rect 35354 13302 35356 13354
rect 35300 13300 35356 13302
rect 35404 13354 35460 13356
rect 35404 13302 35406 13354
rect 35406 13302 35458 13354
rect 35458 13302 35460 13354
rect 35404 13300 35460 13302
rect 35196 11786 35252 11788
rect 35196 11734 35198 11786
rect 35198 11734 35250 11786
rect 35250 11734 35252 11786
rect 35196 11732 35252 11734
rect 35300 11786 35356 11788
rect 35300 11734 35302 11786
rect 35302 11734 35354 11786
rect 35354 11734 35356 11786
rect 35300 11732 35356 11734
rect 35404 11786 35460 11788
rect 35404 11734 35406 11786
rect 35406 11734 35458 11786
rect 35458 11734 35460 11786
rect 35404 11732 35460 11734
rect 35196 10218 35252 10220
rect 35196 10166 35198 10218
rect 35198 10166 35250 10218
rect 35250 10166 35252 10218
rect 35196 10164 35252 10166
rect 35300 10218 35356 10220
rect 35300 10166 35302 10218
rect 35302 10166 35354 10218
rect 35354 10166 35356 10218
rect 35300 10164 35356 10166
rect 35404 10218 35460 10220
rect 35404 10166 35406 10218
rect 35406 10166 35458 10218
rect 35458 10166 35460 10218
rect 35404 10164 35460 10166
rect 35196 8650 35252 8652
rect 35196 8598 35198 8650
rect 35198 8598 35250 8650
rect 35250 8598 35252 8650
rect 35196 8596 35252 8598
rect 35300 8650 35356 8652
rect 35300 8598 35302 8650
rect 35302 8598 35354 8650
rect 35354 8598 35356 8650
rect 35300 8596 35356 8598
rect 35404 8650 35460 8652
rect 35404 8598 35406 8650
rect 35406 8598 35458 8650
rect 35458 8598 35460 8650
rect 35404 8596 35460 8598
rect 19180 3500 19236 3556
rect 20188 4060 20244 4116
rect 19836 3162 19892 3164
rect 19836 3110 19838 3162
rect 19838 3110 19890 3162
rect 19890 3110 19892 3162
rect 19836 3108 19892 3110
rect 19940 3162 19996 3164
rect 19940 3110 19942 3162
rect 19942 3110 19994 3162
rect 19994 3110 19996 3162
rect 19940 3108 19996 3110
rect 20044 3162 20100 3164
rect 20044 3110 20046 3162
rect 20046 3110 20098 3162
rect 20098 3110 20100 3162
rect 20044 3108 20100 3110
rect 21420 4114 21476 4116
rect 21420 4062 21422 4114
rect 21422 4062 21474 4114
rect 21474 4062 21476 4114
rect 21420 4060 21476 4062
rect 23772 3612 23828 3668
rect 35196 7082 35252 7084
rect 35196 7030 35198 7082
rect 35198 7030 35250 7082
rect 35250 7030 35252 7082
rect 35196 7028 35252 7030
rect 35300 7082 35356 7084
rect 35300 7030 35302 7082
rect 35302 7030 35354 7082
rect 35354 7030 35356 7082
rect 35300 7028 35356 7030
rect 35404 7082 35460 7084
rect 35404 7030 35406 7082
rect 35406 7030 35458 7082
rect 35458 7030 35460 7082
rect 35404 7028 35460 7030
rect 35196 5514 35252 5516
rect 35196 5462 35198 5514
rect 35198 5462 35250 5514
rect 35250 5462 35252 5514
rect 35196 5460 35252 5462
rect 35300 5514 35356 5516
rect 35300 5462 35302 5514
rect 35302 5462 35354 5514
rect 35354 5462 35356 5514
rect 35300 5460 35356 5462
rect 35404 5514 35460 5516
rect 35404 5462 35406 5514
rect 35406 5462 35458 5514
rect 35458 5462 35460 5514
rect 35404 5460 35460 5462
rect 24892 4060 24948 4116
rect 26236 4114 26292 4116
rect 26236 4062 26238 4114
rect 26238 4062 26290 4114
rect 26290 4062 26292 4114
rect 26236 4060 26292 4062
rect 35196 3946 35252 3948
rect 35196 3894 35198 3946
rect 35198 3894 35250 3946
rect 35250 3894 35252 3946
rect 35196 3892 35252 3894
rect 35300 3946 35356 3948
rect 35300 3894 35302 3946
rect 35302 3894 35354 3946
rect 35354 3894 35356 3946
rect 35300 3892 35356 3894
rect 35404 3946 35460 3948
rect 35404 3894 35406 3946
rect 35406 3894 35458 3946
rect 35458 3894 35460 3946
rect 35404 3892 35460 3894
rect 25564 3666 25620 3668
rect 25564 3614 25566 3666
rect 25566 3614 25618 3666
rect 25618 3614 25620 3666
rect 25564 3612 25620 3614
<< metal3 >>
rect 4466 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4750 38444
rect 35186 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35470 38444
rect 17490 38220 17500 38276
rect 17556 38220 18620 38276
rect 18676 38220 18686 38276
rect 22866 38220 22876 38276
rect 22932 38220 25564 38276
rect 25620 38220 25630 38276
rect 19506 38108 19516 38164
rect 19572 38108 21868 38164
rect 21924 38108 21934 38164
rect 19618 37996 19628 38052
rect 19684 37996 20748 38052
rect 20804 37996 20814 38052
rect 19826 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20110 37660
rect 14130 37436 14140 37492
rect 14196 37436 15260 37492
rect 15316 37436 15326 37492
rect 24882 37436 24892 37492
rect 24948 37436 26236 37492
rect 26292 37436 26302 37492
rect 4466 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4750 36876
rect 35186 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35470 36876
rect 19826 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20110 36092
rect 4466 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4750 35308
rect 35186 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35470 35308
rect 19826 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20110 34524
rect 4466 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4750 33740
rect 35186 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35470 33740
rect 19826 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20110 32956
rect 4466 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4750 32172
rect 35186 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35470 32172
rect 19826 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20110 31388
rect 4466 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4750 30604
rect 35186 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35470 30604
rect 19826 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20110 29820
rect 4466 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4750 29036
rect 35186 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35470 29036
rect 14018 28588 14028 28644
rect 14084 28588 16716 28644
rect 16772 28588 17500 28644
rect 17556 28588 19964 28644
rect 20020 28588 20030 28644
rect 19826 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20110 28252
rect 10770 27804 10780 27860
rect 10836 27804 14028 27860
rect 14084 27804 14094 27860
rect 20178 27804 20188 27860
rect 20244 27804 22652 27860
rect 22708 27804 23548 27860
rect 23604 27804 25452 27860
rect 25508 27804 26012 27860
rect 26068 27804 26078 27860
rect 14690 27692 14700 27748
rect 14756 27692 15932 27748
rect 15988 27692 15998 27748
rect 21746 27692 21756 27748
rect 21812 27692 22988 27748
rect 23044 27692 24556 27748
rect 24612 27692 24622 27748
rect 0 27636 800 27664
rect 0 27580 4172 27636
rect 4228 27580 4238 27636
rect 0 27552 800 27580
rect 4466 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4750 27468
rect 35186 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35470 27468
rect 11442 27244 11452 27300
rect 11508 27244 15148 27300
rect 15204 27244 15214 27300
rect 13794 27132 13804 27188
rect 13860 27132 14812 27188
rect 14868 27132 14878 27188
rect 16034 27132 16044 27188
rect 16100 27132 16940 27188
rect 16996 27132 17006 27188
rect 14812 27076 14868 27132
rect 13906 27020 13916 27076
rect 13972 27020 14476 27076
rect 14532 27020 14542 27076
rect 14812 27020 16716 27076
rect 16772 27020 16782 27076
rect 27570 27020 27580 27076
rect 27636 27020 28364 27076
rect 28420 27020 37660 27076
rect 37716 27020 37726 27076
rect 14130 26908 14140 26964
rect 14196 26908 14924 26964
rect 14980 26908 14990 26964
rect 17154 26908 17164 26964
rect 17220 26908 18956 26964
rect 19012 26908 19022 26964
rect 15138 26796 15148 26852
rect 15204 26796 20972 26852
rect 21028 26796 22540 26852
rect 22596 26796 22606 26852
rect 26338 26796 26348 26852
rect 26404 26796 27356 26852
rect 27412 26796 27422 26852
rect 19826 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20110 26684
rect 19506 26460 19516 26516
rect 19572 26460 19964 26516
rect 20020 26460 20030 26516
rect 23762 26460 23772 26516
rect 23828 26460 25564 26516
rect 25620 26460 25630 26516
rect 19058 26348 19068 26404
rect 19124 26348 19852 26404
rect 19908 26348 19918 26404
rect 20972 26348 21420 26404
rect 21476 26348 21486 26404
rect 0 26292 800 26320
rect 20972 26292 21028 26348
rect 41200 26292 42000 26320
rect 0 26236 1932 26292
rect 1988 26236 1998 26292
rect 14242 26236 14252 26292
rect 14308 26236 15148 26292
rect 18946 26236 18956 26292
rect 19012 26236 20972 26292
rect 21028 26236 21038 26292
rect 22530 26236 22540 26292
rect 22596 26236 23212 26292
rect 23268 26236 23278 26292
rect 40002 26236 40012 26292
rect 40068 26236 42000 26292
rect 0 26208 800 26236
rect 15092 26180 15148 26236
rect 41200 26208 42000 26236
rect 4274 26124 4284 26180
rect 4340 26124 11452 26180
rect 11508 26124 14812 26180
rect 14868 26124 14878 26180
rect 15092 26124 15372 26180
rect 15428 26124 15438 26180
rect 18722 26124 18732 26180
rect 18788 26124 20524 26180
rect 20580 26124 20590 26180
rect 25666 26124 25676 26180
rect 25732 26124 28812 26180
rect 28868 26124 28878 26180
rect 18274 26012 18284 26068
rect 18340 26012 19180 26068
rect 19236 26012 19246 26068
rect 19590 26012 19628 26068
rect 19684 26012 19694 26068
rect 18722 25900 18732 25956
rect 18788 25900 21980 25956
rect 22036 25900 22046 25956
rect 4466 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4750 25900
rect 35186 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35470 25900
rect 18610 25788 18620 25844
rect 18676 25788 19068 25844
rect 19124 25788 21532 25844
rect 21588 25788 21598 25844
rect 20514 25676 20524 25732
rect 20580 25676 21756 25732
rect 21812 25676 21822 25732
rect 21084 25620 21140 25676
rect 41200 25620 42000 25648
rect 21074 25564 21084 25620
rect 21140 25564 21150 25620
rect 21634 25564 21644 25620
rect 21700 25564 23548 25620
rect 23604 25564 23614 25620
rect 27794 25564 27804 25620
rect 27860 25564 28588 25620
rect 28644 25564 37660 25620
rect 37716 25564 37726 25620
rect 40002 25564 40012 25620
rect 40068 25564 42000 25620
rect 41200 25536 42000 25564
rect 13794 25452 13804 25508
rect 13860 25452 18732 25508
rect 18788 25452 18798 25508
rect 19170 25452 19180 25508
rect 19236 25452 19404 25508
rect 19460 25452 22316 25508
rect 22372 25452 23436 25508
rect 23492 25452 23502 25508
rect 27010 25452 27020 25508
rect 27076 25452 27086 25508
rect 27020 25396 27076 25452
rect 13570 25340 13580 25396
rect 13636 25340 15148 25396
rect 18274 25340 18284 25396
rect 18340 25340 19628 25396
rect 19684 25340 27076 25396
rect 15092 25284 15148 25340
rect 15092 25228 18172 25284
rect 18228 25228 18238 25284
rect 18694 25228 18732 25284
rect 18788 25228 18798 25284
rect 19058 25228 19068 25284
rect 19124 25228 19404 25284
rect 19460 25228 19628 25284
rect 19684 25228 19694 25284
rect 20738 25228 20748 25284
rect 20804 25228 21644 25284
rect 21700 25228 21710 25284
rect 21858 25228 21868 25284
rect 21924 25228 22764 25284
rect 22820 25228 22830 25284
rect 19826 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20110 25116
rect 13458 24892 13468 24948
rect 13524 24892 17388 24948
rect 17444 24892 17454 24948
rect 19366 24892 19404 24948
rect 19460 24892 19470 24948
rect 22082 24892 22092 24948
rect 22148 24892 26236 24948
rect 26292 24892 26302 24948
rect 18274 24780 18284 24836
rect 18340 24780 20468 24836
rect 20412 24724 20468 24780
rect 17938 24668 17948 24724
rect 18004 24668 18396 24724
rect 18452 24668 19068 24724
rect 19124 24668 19134 24724
rect 20402 24668 20412 24724
rect 20468 24668 20478 24724
rect 4466 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4750 24332
rect 35186 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35470 24332
rect 4274 23884 4284 23940
rect 4340 23884 11004 23940
rect 11060 23884 13692 23940
rect 13748 23884 13758 23940
rect 14354 23772 14364 23828
rect 14420 23772 14700 23828
rect 14756 23772 18172 23828
rect 18228 23772 18238 23828
rect 13122 23660 13132 23716
rect 13188 23660 14028 23716
rect 14084 23660 14094 23716
rect 15092 23660 15372 23716
rect 15428 23660 16604 23716
rect 16660 23660 16670 23716
rect 17602 23660 17612 23716
rect 17668 23660 26124 23716
rect 26180 23660 26190 23716
rect 26450 23660 26460 23716
rect 26516 23660 27916 23716
rect 27972 23660 28364 23716
rect 28420 23660 28430 23716
rect 0 23604 800 23632
rect 15092 23604 15148 23660
rect 41200 23604 42000 23632
rect 0 23548 1932 23604
rect 1988 23548 1998 23604
rect 14354 23548 14364 23604
rect 14420 23548 15148 23604
rect 40002 23548 40012 23604
rect 40068 23548 42000 23604
rect 0 23520 800 23548
rect 19826 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20110 23548
rect 41200 23520 42000 23548
rect 20626 23436 20636 23492
rect 20692 23436 21308 23492
rect 21364 23436 21374 23492
rect 21308 23380 21364 23436
rect 21308 23324 21980 23380
rect 22036 23324 22046 23380
rect 15586 23212 15596 23268
rect 15652 23212 17836 23268
rect 17892 23212 17902 23268
rect 14130 23100 14140 23156
rect 14196 23100 15372 23156
rect 15428 23100 16044 23156
rect 16100 23100 16110 23156
rect 18722 23100 18732 23156
rect 18788 23100 20524 23156
rect 20580 23100 20590 23156
rect 16818 22988 16828 23044
rect 16884 22988 17500 23044
rect 17556 22988 19068 23044
rect 19124 22988 19134 23044
rect 24658 22988 24668 23044
rect 24724 22988 37324 23044
rect 37380 22988 37390 23044
rect 41200 22932 42000 22960
rect 4162 22876 4172 22932
rect 4228 22876 8428 22932
rect 18834 22876 18844 22932
rect 18900 22876 19180 22932
rect 19236 22876 21420 22932
rect 21476 22876 21486 22932
rect 40002 22876 40012 22932
rect 40068 22876 42000 22932
rect 4466 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4750 22764
rect 8372 22372 8428 22876
rect 41200 22848 42000 22876
rect 35186 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35470 22764
rect 15250 22652 15260 22708
rect 15316 22652 19628 22708
rect 19684 22652 19694 22708
rect 20178 22652 20188 22708
rect 20244 22652 20748 22708
rect 20804 22652 20814 22708
rect 21298 22652 21308 22708
rect 21364 22652 21644 22708
rect 21700 22652 21710 22708
rect 17266 22540 17276 22596
rect 17332 22540 18284 22596
rect 18340 22540 18350 22596
rect 18834 22540 18844 22596
rect 18900 22540 22316 22596
rect 22372 22540 22382 22596
rect 8372 22316 19068 22372
rect 19124 22316 20748 22372
rect 20804 22316 20814 22372
rect 21410 22316 21420 22372
rect 21476 22316 22540 22372
rect 22596 22316 22606 22372
rect 41200 22260 42000 22288
rect 16930 22204 16940 22260
rect 16996 22204 17612 22260
rect 17668 22204 17678 22260
rect 17826 22204 17836 22260
rect 17892 22204 18844 22260
rect 18900 22204 18910 22260
rect 40002 22204 40012 22260
rect 40068 22204 42000 22260
rect 41200 22176 42000 22204
rect 29586 22092 29596 22148
rect 29652 22092 37884 22148
rect 37940 22092 37950 22148
rect 20178 21980 20188 22036
rect 20244 21980 22316 22036
rect 22372 21980 25452 22036
rect 25508 21980 25518 22036
rect 28242 21980 28252 22036
rect 28308 21980 29372 22036
rect 29428 21980 29932 22036
rect 29988 21980 37660 22036
rect 37716 21980 37726 22036
rect 19826 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20110 21980
rect 18172 21868 19628 21924
rect 19684 21868 19694 21924
rect 21858 21868 21868 21924
rect 21924 21868 23996 21924
rect 24052 21868 25340 21924
rect 25396 21868 26684 21924
rect 26740 21868 26750 21924
rect 18172 21812 18228 21868
rect 11330 21756 11340 21812
rect 11396 21756 14588 21812
rect 14644 21756 15372 21812
rect 15428 21756 15438 21812
rect 15922 21756 15932 21812
rect 15988 21756 17164 21812
rect 17220 21756 17724 21812
rect 17780 21756 18172 21812
rect 18228 21756 18238 21812
rect 20178 21756 20188 21812
rect 20244 21756 21308 21812
rect 21364 21756 21374 21812
rect 22306 21756 22316 21812
rect 22372 21756 24556 21812
rect 24612 21756 24622 21812
rect 25890 21756 25900 21812
rect 25956 21756 26572 21812
rect 26628 21756 31948 21812
rect 14914 21644 14924 21700
rect 14980 21644 15708 21700
rect 15764 21644 15774 21700
rect 16818 21644 16828 21700
rect 16884 21644 17948 21700
rect 18004 21644 19292 21700
rect 19348 21644 19358 21700
rect 24658 21644 24668 21700
rect 24724 21644 25340 21700
rect 25396 21644 25406 21700
rect 31892 21588 31948 21756
rect 41200 21588 42000 21616
rect 12002 21532 12012 21588
rect 12068 21532 20300 21588
rect 20356 21532 20366 21588
rect 22978 21532 22988 21588
rect 23044 21532 25564 21588
rect 25620 21532 25630 21588
rect 31892 21532 37660 21588
rect 37716 21532 37726 21588
rect 40002 21532 40012 21588
rect 40068 21532 42000 21588
rect 41200 21504 42000 21532
rect 17378 21420 17388 21476
rect 17444 21420 18172 21476
rect 18228 21420 18620 21476
rect 18676 21420 25228 21476
rect 25284 21420 25294 21476
rect 25330 21308 25340 21364
rect 25396 21308 27916 21364
rect 27972 21308 27982 21364
rect 4466 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4750 21196
rect 35186 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35470 21196
rect 20066 20748 20076 20804
rect 20132 20748 22876 20804
rect 22932 20748 22942 20804
rect 21522 20524 21532 20580
rect 21588 20524 22316 20580
rect 22372 20524 22382 20580
rect 18946 20412 18956 20468
rect 19012 20412 19404 20468
rect 19460 20412 19470 20468
rect 19826 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20110 20412
rect 18386 20188 18396 20244
rect 18452 20188 25340 20244
rect 25396 20188 25406 20244
rect 19058 20076 19068 20132
rect 19124 20076 21756 20132
rect 21812 20076 23660 20132
rect 23716 20076 23726 20132
rect 18050 19964 18060 20020
rect 18116 19964 19964 20020
rect 20020 19964 20524 20020
rect 20580 19964 20590 20020
rect 20962 19964 20972 20020
rect 21028 19964 21420 20020
rect 21476 19964 21486 20020
rect 22082 19964 22092 20020
rect 22148 19964 23772 20020
rect 23828 19964 25676 20020
rect 25732 19964 25742 20020
rect 31892 19964 37660 20020
rect 37716 19964 37726 20020
rect 31892 19908 31948 19964
rect 19282 19852 19292 19908
rect 19348 19852 21308 19908
rect 21364 19852 21374 19908
rect 29138 19852 29148 19908
rect 29204 19852 31948 19908
rect 17154 19740 17164 19796
rect 17220 19740 20636 19796
rect 20692 19740 21196 19796
rect 21252 19740 21262 19796
rect 4466 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4750 19628
rect 35186 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35470 19628
rect 41200 19572 42000 19600
rect 40002 19516 40012 19572
rect 40068 19516 42000 19572
rect 41200 19488 42000 19516
rect 14690 19404 14700 19460
rect 14756 19404 15148 19460
rect 17602 19404 17612 19460
rect 17668 19404 18620 19460
rect 18676 19404 18686 19460
rect 15092 19348 15148 19404
rect 15092 19292 18172 19348
rect 18228 19292 18238 19348
rect 16930 19180 16940 19236
rect 16996 19180 18508 19236
rect 18564 19180 18574 19236
rect 15922 19068 15932 19124
rect 15988 19068 18732 19124
rect 18788 19068 18798 19124
rect 19394 19068 19404 19124
rect 19460 19068 20076 19124
rect 20132 19068 22428 19124
rect 22484 19068 22494 19124
rect 25890 19068 25900 19124
rect 25956 19068 29148 19124
rect 29204 19068 29214 19124
rect 17714 18956 17724 19012
rect 17780 18956 19292 19012
rect 19348 18956 19358 19012
rect 41200 18900 42000 18928
rect 21746 18844 21756 18900
rect 21812 18844 23548 18900
rect 23604 18844 24892 18900
rect 24948 18844 24958 18900
rect 40002 18844 40012 18900
rect 40068 18844 42000 18900
rect 19826 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20110 18844
rect 41200 18816 42000 18844
rect 20738 18732 20748 18788
rect 20804 18732 22204 18788
rect 22260 18732 22270 18788
rect 22428 18732 26684 18788
rect 26740 18732 26750 18788
rect 22428 18676 22484 18732
rect 17826 18620 17836 18676
rect 17892 18620 19852 18676
rect 19908 18620 20300 18676
rect 20356 18620 20366 18676
rect 20738 18620 20748 18676
rect 20804 18620 22092 18676
rect 22148 18620 22484 18676
rect 23202 18620 23212 18676
rect 23268 18620 24108 18676
rect 24164 18620 24556 18676
rect 24612 18620 25228 18676
rect 25284 18620 25294 18676
rect 18162 18508 18172 18564
rect 18228 18508 23884 18564
rect 23940 18508 23950 18564
rect 16482 18396 16492 18452
rect 16548 18396 17500 18452
rect 17556 18396 17724 18452
rect 17780 18396 17790 18452
rect 18610 18396 18620 18452
rect 18676 18396 19180 18452
rect 19236 18396 20076 18452
rect 20132 18396 20142 18452
rect 20850 18396 20860 18452
rect 20916 18396 22652 18452
rect 22708 18396 22718 18452
rect 23202 18396 23212 18452
rect 23268 18396 23996 18452
rect 24052 18396 24062 18452
rect 25554 18396 25564 18452
rect 25620 18396 26236 18452
rect 26292 18396 28588 18452
rect 28644 18396 29596 18452
rect 29652 18396 29662 18452
rect 15026 18284 15036 18340
rect 15092 18284 16268 18340
rect 16324 18284 16716 18340
rect 16772 18284 16782 18340
rect 19394 18284 19404 18340
rect 19460 18284 21980 18340
rect 22036 18284 23548 18340
rect 23604 18284 24444 18340
rect 24500 18284 24510 18340
rect 24994 18284 25004 18340
rect 25060 18284 26012 18340
rect 26068 18284 26078 18340
rect 41200 18228 42000 18256
rect 14466 18172 14476 18228
rect 14532 18172 15596 18228
rect 15652 18172 15662 18228
rect 19618 18172 19628 18228
rect 19684 18172 20188 18228
rect 20244 18172 21420 18228
rect 21476 18172 21486 18228
rect 25442 18172 25452 18228
rect 25508 18172 28140 18228
rect 28196 18172 37884 18228
rect 37940 18172 37950 18228
rect 40002 18172 40012 18228
rect 40068 18172 42000 18228
rect 41200 18144 42000 18172
rect 21746 18060 21756 18116
rect 21812 18060 26572 18116
rect 26628 18060 26638 18116
rect 4466 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4750 18060
rect 35186 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35470 18060
rect 31892 17836 37660 17892
rect 37716 17836 37726 17892
rect 31892 17780 31948 17836
rect 12898 17724 12908 17780
rect 12964 17724 18732 17780
rect 18788 17724 20300 17780
rect 20356 17724 20366 17780
rect 24098 17724 24108 17780
rect 24164 17724 24892 17780
rect 24948 17724 31948 17780
rect 15138 17612 15148 17668
rect 15204 17612 15596 17668
rect 15652 17612 15662 17668
rect 18834 17612 18844 17668
rect 18900 17612 19404 17668
rect 19460 17612 19470 17668
rect 24770 17612 24780 17668
rect 24836 17612 25788 17668
rect 25844 17612 26460 17668
rect 26516 17612 26526 17668
rect 28466 17612 28476 17668
rect 28532 17612 29484 17668
rect 29540 17612 37660 17668
rect 37716 17612 37726 17668
rect 41200 17556 42000 17584
rect 17042 17500 17052 17556
rect 17108 17500 18060 17556
rect 18116 17500 18508 17556
rect 18564 17500 18574 17556
rect 40002 17500 40012 17556
rect 40068 17500 42000 17556
rect 41200 17472 42000 17500
rect 15362 17388 15372 17444
rect 15428 17388 18956 17444
rect 19012 17388 19022 17444
rect 19826 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20110 17276
rect 21970 17052 21980 17108
rect 22036 17052 25340 17108
rect 25396 17052 26236 17108
rect 26292 17052 26302 17108
rect 12898 16940 12908 16996
rect 12964 16940 14476 16996
rect 14532 16940 14542 16996
rect 12226 16828 12236 16884
rect 12292 16828 15484 16884
rect 15540 16828 15550 16884
rect 4466 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4750 16492
rect 35186 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35470 16492
rect 19826 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20110 15708
rect 24210 15484 24220 15540
rect 24276 15484 25676 15540
rect 25732 15484 25742 15540
rect 26114 15484 26124 15540
rect 26180 15484 26796 15540
rect 26852 15484 26862 15540
rect 26124 15428 26180 15484
rect 16482 15372 16492 15428
rect 16548 15372 17388 15428
rect 17444 15372 21868 15428
rect 21924 15372 26180 15428
rect 18162 15260 18172 15316
rect 18228 15260 18844 15316
rect 18900 15260 18910 15316
rect 13906 15148 13916 15204
rect 13972 15148 16268 15204
rect 16324 15148 16334 15204
rect 18386 15148 18396 15204
rect 18452 15148 19964 15204
rect 20020 15148 20030 15204
rect 25890 14924 25900 14980
rect 25956 14924 26908 14980
rect 26964 14924 26974 14980
rect 4466 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4750 14924
rect 35186 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35470 14924
rect 41200 14868 42000 14896
rect 40002 14812 40012 14868
rect 40068 14812 42000 14868
rect 41200 14784 42000 14812
rect 27010 14700 27020 14756
rect 27076 14700 27804 14756
rect 27860 14700 37660 14756
rect 37716 14700 37726 14756
rect 24994 14588 25004 14644
rect 25060 14588 26572 14644
rect 26628 14588 28252 14644
rect 28308 14588 28318 14644
rect 18274 14476 18284 14532
rect 18340 14476 19852 14532
rect 19908 14476 19918 14532
rect 20178 14476 20188 14532
rect 20244 14476 21868 14532
rect 21924 14476 22204 14532
rect 22260 14476 22270 14532
rect 22418 14476 22428 14532
rect 22484 14476 23660 14532
rect 23716 14476 23726 14532
rect 19954 14364 19964 14420
rect 20020 14364 21252 14420
rect 21410 14364 21420 14420
rect 21476 14364 23212 14420
rect 23268 14364 23278 14420
rect 21196 14308 21252 14364
rect 13346 14252 13356 14308
rect 13412 14252 15484 14308
rect 15540 14252 16268 14308
rect 16324 14252 16828 14308
rect 16884 14252 17612 14308
rect 17668 14252 20636 14308
rect 20692 14252 20702 14308
rect 21196 14252 21756 14308
rect 21812 14252 22652 14308
rect 22708 14252 22718 14308
rect 19826 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20110 14140
rect 21298 13804 21308 13860
rect 21364 13804 24220 13860
rect 24276 13804 24286 13860
rect 23538 13580 23548 13636
rect 23604 13580 24668 13636
rect 24724 13580 25228 13636
rect 25284 13580 25294 13636
rect 21858 13468 21868 13524
rect 21924 13468 21934 13524
rect 21868 13412 21924 13468
rect 21410 13356 21420 13412
rect 21476 13356 21924 13412
rect 4466 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4750 13356
rect 35186 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35470 13356
rect 19618 13132 19628 13188
rect 19684 13132 20524 13188
rect 20580 13132 20590 13188
rect 19826 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20110 12572
rect 16034 12460 16044 12516
rect 16100 12460 17388 12516
rect 17444 12460 17454 12516
rect 4466 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4750 11788
rect 35186 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35470 11788
rect 19826 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20110 11004
rect 4466 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4750 10220
rect 35186 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35470 10220
rect 19826 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20110 9436
rect 4466 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4750 8652
rect 35186 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35470 8652
rect 19826 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20110 7868
rect 4466 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4750 7084
rect 35186 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35470 7084
rect 19826 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20110 6300
rect 4466 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4750 5516
rect 35186 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35470 5516
rect 19826 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20110 4732
rect 16146 4172 16156 4228
rect 16212 4172 18508 4228
rect 18564 4172 18574 4228
rect 20178 4060 20188 4116
rect 20244 4060 21420 4116
rect 21476 4060 21486 4116
rect 24882 4060 24892 4116
rect 24948 4060 26236 4116
rect 26292 4060 26302 4116
rect 4466 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4750 3948
rect 35186 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35470 3948
rect 23762 3612 23772 3668
rect 23828 3612 25564 3668
rect 25620 3612 25630 3668
rect 18050 3500 18060 3556
rect 18116 3500 19180 3556
rect 19236 3500 19246 3556
rect 19826 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20110 3164
<< via3 >>
rect 4476 38388 4532 38444
rect 4580 38388 4636 38444
rect 4684 38388 4740 38444
rect 35196 38388 35252 38444
rect 35300 38388 35356 38444
rect 35404 38388 35460 38444
rect 19836 37604 19892 37660
rect 19940 37604 19996 37660
rect 20044 37604 20100 37660
rect 4476 36820 4532 36876
rect 4580 36820 4636 36876
rect 4684 36820 4740 36876
rect 35196 36820 35252 36876
rect 35300 36820 35356 36876
rect 35404 36820 35460 36876
rect 19836 36036 19892 36092
rect 19940 36036 19996 36092
rect 20044 36036 20100 36092
rect 4476 35252 4532 35308
rect 4580 35252 4636 35308
rect 4684 35252 4740 35308
rect 35196 35252 35252 35308
rect 35300 35252 35356 35308
rect 35404 35252 35460 35308
rect 19836 34468 19892 34524
rect 19940 34468 19996 34524
rect 20044 34468 20100 34524
rect 4476 33684 4532 33740
rect 4580 33684 4636 33740
rect 4684 33684 4740 33740
rect 35196 33684 35252 33740
rect 35300 33684 35356 33740
rect 35404 33684 35460 33740
rect 19836 32900 19892 32956
rect 19940 32900 19996 32956
rect 20044 32900 20100 32956
rect 4476 32116 4532 32172
rect 4580 32116 4636 32172
rect 4684 32116 4740 32172
rect 35196 32116 35252 32172
rect 35300 32116 35356 32172
rect 35404 32116 35460 32172
rect 19836 31332 19892 31388
rect 19940 31332 19996 31388
rect 20044 31332 20100 31388
rect 4476 30548 4532 30604
rect 4580 30548 4636 30604
rect 4684 30548 4740 30604
rect 35196 30548 35252 30604
rect 35300 30548 35356 30604
rect 35404 30548 35460 30604
rect 19836 29764 19892 29820
rect 19940 29764 19996 29820
rect 20044 29764 20100 29820
rect 4476 28980 4532 29036
rect 4580 28980 4636 29036
rect 4684 28980 4740 29036
rect 35196 28980 35252 29036
rect 35300 28980 35356 29036
rect 35404 28980 35460 29036
rect 19836 28196 19892 28252
rect 19940 28196 19996 28252
rect 20044 28196 20100 28252
rect 4476 27412 4532 27468
rect 4580 27412 4636 27468
rect 4684 27412 4740 27468
rect 35196 27412 35252 27468
rect 35300 27412 35356 27468
rect 35404 27412 35460 27468
rect 19836 26628 19892 26684
rect 19940 26628 19996 26684
rect 20044 26628 20100 26684
rect 19628 26012 19684 26068
rect 4476 25844 4532 25900
rect 4580 25844 4636 25900
rect 4684 25844 4740 25900
rect 35196 25844 35252 25900
rect 35300 25844 35356 25900
rect 35404 25844 35460 25900
rect 19404 25452 19460 25508
rect 18732 25228 18788 25284
rect 19628 25228 19684 25284
rect 19836 25060 19892 25116
rect 19940 25060 19996 25116
rect 20044 25060 20100 25116
rect 19404 24892 19460 24948
rect 4476 24276 4532 24332
rect 4580 24276 4636 24332
rect 4684 24276 4740 24332
rect 35196 24276 35252 24332
rect 35300 24276 35356 24332
rect 35404 24276 35460 24332
rect 19836 23492 19892 23548
rect 19940 23492 19996 23548
rect 20044 23492 20100 23548
rect 4476 22708 4532 22764
rect 4580 22708 4636 22764
rect 4684 22708 4740 22764
rect 35196 22708 35252 22764
rect 35300 22708 35356 22764
rect 35404 22708 35460 22764
rect 20748 22652 20804 22708
rect 19836 21924 19892 21980
rect 19940 21924 19996 21980
rect 20044 21924 20100 21980
rect 4476 21140 4532 21196
rect 4580 21140 4636 21196
rect 4684 21140 4740 21196
rect 35196 21140 35252 21196
rect 35300 21140 35356 21196
rect 35404 21140 35460 21196
rect 19836 20356 19892 20412
rect 19940 20356 19996 20412
rect 20044 20356 20100 20412
rect 4476 19572 4532 19628
rect 4580 19572 4636 19628
rect 4684 19572 4740 19628
rect 35196 19572 35252 19628
rect 35300 19572 35356 19628
rect 35404 19572 35460 19628
rect 19836 18788 19892 18844
rect 19940 18788 19996 18844
rect 20044 18788 20100 18844
rect 20748 18620 20804 18676
rect 4476 18004 4532 18060
rect 4580 18004 4636 18060
rect 4684 18004 4740 18060
rect 35196 18004 35252 18060
rect 35300 18004 35356 18060
rect 35404 18004 35460 18060
rect 18732 17724 18788 17780
rect 19836 17220 19892 17276
rect 19940 17220 19996 17276
rect 20044 17220 20100 17276
rect 4476 16436 4532 16492
rect 4580 16436 4636 16492
rect 4684 16436 4740 16492
rect 35196 16436 35252 16492
rect 35300 16436 35356 16492
rect 35404 16436 35460 16492
rect 19836 15652 19892 15708
rect 19940 15652 19996 15708
rect 20044 15652 20100 15708
rect 4476 14868 4532 14924
rect 4580 14868 4636 14924
rect 4684 14868 4740 14924
rect 35196 14868 35252 14924
rect 35300 14868 35356 14924
rect 35404 14868 35460 14924
rect 19836 14084 19892 14140
rect 19940 14084 19996 14140
rect 20044 14084 20100 14140
rect 4476 13300 4532 13356
rect 4580 13300 4636 13356
rect 4684 13300 4740 13356
rect 35196 13300 35252 13356
rect 35300 13300 35356 13356
rect 35404 13300 35460 13356
rect 19836 12516 19892 12572
rect 19940 12516 19996 12572
rect 20044 12516 20100 12572
rect 4476 11732 4532 11788
rect 4580 11732 4636 11788
rect 4684 11732 4740 11788
rect 35196 11732 35252 11788
rect 35300 11732 35356 11788
rect 35404 11732 35460 11788
rect 19836 10948 19892 11004
rect 19940 10948 19996 11004
rect 20044 10948 20100 11004
rect 4476 10164 4532 10220
rect 4580 10164 4636 10220
rect 4684 10164 4740 10220
rect 35196 10164 35252 10220
rect 35300 10164 35356 10220
rect 35404 10164 35460 10220
rect 19836 9380 19892 9436
rect 19940 9380 19996 9436
rect 20044 9380 20100 9436
rect 4476 8596 4532 8652
rect 4580 8596 4636 8652
rect 4684 8596 4740 8652
rect 35196 8596 35252 8652
rect 35300 8596 35356 8652
rect 35404 8596 35460 8652
rect 19836 7812 19892 7868
rect 19940 7812 19996 7868
rect 20044 7812 20100 7868
rect 4476 7028 4532 7084
rect 4580 7028 4636 7084
rect 4684 7028 4740 7084
rect 35196 7028 35252 7084
rect 35300 7028 35356 7084
rect 35404 7028 35460 7084
rect 19836 6244 19892 6300
rect 19940 6244 19996 6300
rect 20044 6244 20100 6300
rect 4476 5460 4532 5516
rect 4580 5460 4636 5516
rect 4684 5460 4740 5516
rect 35196 5460 35252 5516
rect 35300 5460 35356 5516
rect 35404 5460 35460 5516
rect 19836 4676 19892 4732
rect 19940 4676 19996 4732
rect 20044 4676 20100 4732
rect 4476 3892 4532 3948
rect 4580 3892 4636 3948
rect 4684 3892 4740 3948
rect 35196 3892 35252 3948
rect 35300 3892 35356 3948
rect 35404 3892 35460 3948
rect 19836 3108 19892 3164
rect 19940 3108 19996 3164
rect 20044 3108 20100 3164
<< metal4 >>
rect 4448 38444 4768 38476
rect 4448 38388 4476 38444
rect 4532 38388 4580 38444
rect 4636 38388 4684 38444
rect 4740 38388 4768 38444
rect 4448 36876 4768 38388
rect 4448 36820 4476 36876
rect 4532 36820 4580 36876
rect 4636 36820 4684 36876
rect 4740 36820 4768 36876
rect 4448 35308 4768 36820
rect 4448 35252 4476 35308
rect 4532 35252 4580 35308
rect 4636 35252 4684 35308
rect 4740 35252 4768 35308
rect 4448 33740 4768 35252
rect 4448 33684 4476 33740
rect 4532 33684 4580 33740
rect 4636 33684 4684 33740
rect 4740 33684 4768 33740
rect 4448 32172 4768 33684
rect 4448 32116 4476 32172
rect 4532 32116 4580 32172
rect 4636 32116 4684 32172
rect 4740 32116 4768 32172
rect 4448 30604 4768 32116
rect 4448 30548 4476 30604
rect 4532 30548 4580 30604
rect 4636 30548 4684 30604
rect 4740 30548 4768 30604
rect 4448 29036 4768 30548
rect 4448 28980 4476 29036
rect 4532 28980 4580 29036
rect 4636 28980 4684 29036
rect 4740 28980 4768 29036
rect 4448 27468 4768 28980
rect 4448 27412 4476 27468
rect 4532 27412 4580 27468
rect 4636 27412 4684 27468
rect 4740 27412 4768 27468
rect 4448 25900 4768 27412
rect 19808 37660 20128 38476
rect 19808 37604 19836 37660
rect 19892 37604 19940 37660
rect 19996 37604 20044 37660
rect 20100 37604 20128 37660
rect 19808 36092 20128 37604
rect 19808 36036 19836 36092
rect 19892 36036 19940 36092
rect 19996 36036 20044 36092
rect 20100 36036 20128 36092
rect 19808 34524 20128 36036
rect 19808 34468 19836 34524
rect 19892 34468 19940 34524
rect 19996 34468 20044 34524
rect 20100 34468 20128 34524
rect 19808 32956 20128 34468
rect 19808 32900 19836 32956
rect 19892 32900 19940 32956
rect 19996 32900 20044 32956
rect 20100 32900 20128 32956
rect 19808 31388 20128 32900
rect 19808 31332 19836 31388
rect 19892 31332 19940 31388
rect 19996 31332 20044 31388
rect 20100 31332 20128 31388
rect 19808 29820 20128 31332
rect 19808 29764 19836 29820
rect 19892 29764 19940 29820
rect 19996 29764 20044 29820
rect 20100 29764 20128 29820
rect 19808 28252 20128 29764
rect 19808 28196 19836 28252
rect 19892 28196 19940 28252
rect 19996 28196 20044 28252
rect 20100 28196 20128 28252
rect 19808 26684 20128 28196
rect 19808 26628 19836 26684
rect 19892 26628 19940 26684
rect 19996 26628 20044 26684
rect 20100 26628 20128 26684
rect 4448 25844 4476 25900
rect 4532 25844 4580 25900
rect 4636 25844 4684 25900
rect 4740 25844 4768 25900
rect 4448 24332 4768 25844
rect 19628 26068 19684 26078
rect 19404 25508 19460 25518
rect 4448 24276 4476 24332
rect 4532 24276 4580 24332
rect 4636 24276 4684 24332
rect 4740 24276 4768 24332
rect 4448 22764 4768 24276
rect 4448 22708 4476 22764
rect 4532 22708 4580 22764
rect 4636 22708 4684 22764
rect 4740 22708 4768 22764
rect 4448 21196 4768 22708
rect 4448 21140 4476 21196
rect 4532 21140 4580 21196
rect 4636 21140 4684 21196
rect 4740 21140 4768 21196
rect 4448 19628 4768 21140
rect 4448 19572 4476 19628
rect 4532 19572 4580 19628
rect 4636 19572 4684 19628
rect 4740 19572 4768 19628
rect 4448 18060 4768 19572
rect 4448 18004 4476 18060
rect 4532 18004 4580 18060
rect 4636 18004 4684 18060
rect 4740 18004 4768 18060
rect 4448 16492 4768 18004
rect 18732 25284 18788 25294
rect 18732 17780 18788 25228
rect 19404 24948 19460 25452
rect 19628 25284 19684 26012
rect 19628 25218 19684 25228
rect 19404 24882 19460 24892
rect 19808 25116 20128 26628
rect 19808 25060 19836 25116
rect 19892 25060 19940 25116
rect 19996 25060 20044 25116
rect 20100 25060 20128 25116
rect 18732 17714 18788 17724
rect 19808 23548 20128 25060
rect 19808 23492 19836 23548
rect 19892 23492 19940 23548
rect 19996 23492 20044 23548
rect 20100 23492 20128 23548
rect 19808 21980 20128 23492
rect 35168 38444 35488 38476
rect 35168 38388 35196 38444
rect 35252 38388 35300 38444
rect 35356 38388 35404 38444
rect 35460 38388 35488 38444
rect 35168 36876 35488 38388
rect 35168 36820 35196 36876
rect 35252 36820 35300 36876
rect 35356 36820 35404 36876
rect 35460 36820 35488 36876
rect 35168 35308 35488 36820
rect 35168 35252 35196 35308
rect 35252 35252 35300 35308
rect 35356 35252 35404 35308
rect 35460 35252 35488 35308
rect 35168 33740 35488 35252
rect 35168 33684 35196 33740
rect 35252 33684 35300 33740
rect 35356 33684 35404 33740
rect 35460 33684 35488 33740
rect 35168 32172 35488 33684
rect 35168 32116 35196 32172
rect 35252 32116 35300 32172
rect 35356 32116 35404 32172
rect 35460 32116 35488 32172
rect 35168 30604 35488 32116
rect 35168 30548 35196 30604
rect 35252 30548 35300 30604
rect 35356 30548 35404 30604
rect 35460 30548 35488 30604
rect 35168 29036 35488 30548
rect 35168 28980 35196 29036
rect 35252 28980 35300 29036
rect 35356 28980 35404 29036
rect 35460 28980 35488 29036
rect 35168 27468 35488 28980
rect 35168 27412 35196 27468
rect 35252 27412 35300 27468
rect 35356 27412 35404 27468
rect 35460 27412 35488 27468
rect 35168 25900 35488 27412
rect 35168 25844 35196 25900
rect 35252 25844 35300 25900
rect 35356 25844 35404 25900
rect 35460 25844 35488 25900
rect 35168 24332 35488 25844
rect 35168 24276 35196 24332
rect 35252 24276 35300 24332
rect 35356 24276 35404 24332
rect 35460 24276 35488 24332
rect 35168 22764 35488 24276
rect 19808 21924 19836 21980
rect 19892 21924 19940 21980
rect 19996 21924 20044 21980
rect 20100 21924 20128 21980
rect 19808 20412 20128 21924
rect 19808 20356 19836 20412
rect 19892 20356 19940 20412
rect 19996 20356 20044 20412
rect 20100 20356 20128 20412
rect 19808 18844 20128 20356
rect 19808 18788 19836 18844
rect 19892 18788 19940 18844
rect 19996 18788 20044 18844
rect 20100 18788 20128 18844
rect 4448 16436 4476 16492
rect 4532 16436 4580 16492
rect 4636 16436 4684 16492
rect 4740 16436 4768 16492
rect 4448 14924 4768 16436
rect 4448 14868 4476 14924
rect 4532 14868 4580 14924
rect 4636 14868 4684 14924
rect 4740 14868 4768 14924
rect 4448 13356 4768 14868
rect 4448 13300 4476 13356
rect 4532 13300 4580 13356
rect 4636 13300 4684 13356
rect 4740 13300 4768 13356
rect 4448 11788 4768 13300
rect 4448 11732 4476 11788
rect 4532 11732 4580 11788
rect 4636 11732 4684 11788
rect 4740 11732 4768 11788
rect 4448 10220 4768 11732
rect 4448 10164 4476 10220
rect 4532 10164 4580 10220
rect 4636 10164 4684 10220
rect 4740 10164 4768 10220
rect 4448 8652 4768 10164
rect 4448 8596 4476 8652
rect 4532 8596 4580 8652
rect 4636 8596 4684 8652
rect 4740 8596 4768 8652
rect 4448 7084 4768 8596
rect 4448 7028 4476 7084
rect 4532 7028 4580 7084
rect 4636 7028 4684 7084
rect 4740 7028 4768 7084
rect 4448 5516 4768 7028
rect 4448 5460 4476 5516
rect 4532 5460 4580 5516
rect 4636 5460 4684 5516
rect 4740 5460 4768 5516
rect 4448 3948 4768 5460
rect 4448 3892 4476 3948
rect 4532 3892 4580 3948
rect 4636 3892 4684 3948
rect 4740 3892 4768 3948
rect 4448 3076 4768 3892
rect 19808 17276 20128 18788
rect 20748 22708 20804 22718
rect 20748 18676 20804 22652
rect 20748 18610 20804 18620
rect 35168 22708 35196 22764
rect 35252 22708 35300 22764
rect 35356 22708 35404 22764
rect 35460 22708 35488 22764
rect 35168 21196 35488 22708
rect 35168 21140 35196 21196
rect 35252 21140 35300 21196
rect 35356 21140 35404 21196
rect 35460 21140 35488 21196
rect 35168 19628 35488 21140
rect 35168 19572 35196 19628
rect 35252 19572 35300 19628
rect 35356 19572 35404 19628
rect 35460 19572 35488 19628
rect 19808 17220 19836 17276
rect 19892 17220 19940 17276
rect 19996 17220 20044 17276
rect 20100 17220 20128 17276
rect 19808 15708 20128 17220
rect 19808 15652 19836 15708
rect 19892 15652 19940 15708
rect 19996 15652 20044 15708
rect 20100 15652 20128 15708
rect 19808 14140 20128 15652
rect 19808 14084 19836 14140
rect 19892 14084 19940 14140
rect 19996 14084 20044 14140
rect 20100 14084 20128 14140
rect 19808 12572 20128 14084
rect 19808 12516 19836 12572
rect 19892 12516 19940 12572
rect 19996 12516 20044 12572
rect 20100 12516 20128 12572
rect 19808 11004 20128 12516
rect 19808 10948 19836 11004
rect 19892 10948 19940 11004
rect 19996 10948 20044 11004
rect 20100 10948 20128 11004
rect 19808 9436 20128 10948
rect 19808 9380 19836 9436
rect 19892 9380 19940 9436
rect 19996 9380 20044 9436
rect 20100 9380 20128 9436
rect 19808 7868 20128 9380
rect 19808 7812 19836 7868
rect 19892 7812 19940 7868
rect 19996 7812 20044 7868
rect 20100 7812 20128 7868
rect 19808 6300 20128 7812
rect 19808 6244 19836 6300
rect 19892 6244 19940 6300
rect 19996 6244 20044 6300
rect 20100 6244 20128 6300
rect 19808 4732 20128 6244
rect 19808 4676 19836 4732
rect 19892 4676 19940 4732
rect 19996 4676 20044 4732
rect 20100 4676 20128 4732
rect 19808 3164 20128 4676
rect 19808 3108 19836 3164
rect 19892 3108 19940 3164
rect 19996 3108 20044 3164
rect 20100 3108 20128 3164
rect 19808 3076 20128 3108
rect 35168 18060 35488 19572
rect 35168 18004 35196 18060
rect 35252 18004 35300 18060
rect 35356 18004 35404 18060
rect 35460 18004 35488 18060
rect 35168 16492 35488 18004
rect 35168 16436 35196 16492
rect 35252 16436 35300 16492
rect 35356 16436 35404 16492
rect 35460 16436 35488 16492
rect 35168 14924 35488 16436
rect 35168 14868 35196 14924
rect 35252 14868 35300 14924
rect 35356 14868 35404 14924
rect 35460 14868 35488 14924
rect 35168 13356 35488 14868
rect 35168 13300 35196 13356
rect 35252 13300 35300 13356
rect 35356 13300 35404 13356
rect 35460 13300 35488 13356
rect 35168 11788 35488 13300
rect 35168 11732 35196 11788
rect 35252 11732 35300 11788
rect 35356 11732 35404 11788
rect 35460 11732 35488 11788
rect 35168 10220 35488 11732
rect 35168 10164 35196 10220
rect 35252 10164 35300 10220
rect 35356 10164 35404 10220
rect 35460 10164 35488 10220
rect 35168 8652 35488 10164
rect 35168 8596 35196 8652
rect 35252 8596 35300 8652
rect 35356 8596 35404 8652
rect 35460 8596 35488 8652
rect 35168 7084 35488 8596
rect 35168 7028 35196 7084
rect 35252 7028 35300 7084
rect 35356 7028 35404 7084
rect 35460 7028 35488 7084
rect 35168 5516 35488 7028
rect 35168 5460 35196 5516
rect 35252 5460 35300 5516
rect 35356 5460 35404 5516
rect 35460 5460 35488 5516
rect 35168 3948 35488 5460
rect 35168 3892 35196 3948
rect 35252 3892 35300 3948
rect 35356 3892 35404 3948
rect 35460 3892 35488 3948
rect 35168 3076 35488 3892
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _111_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 15456 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__inv_1  _112_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19152 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _113_
timestamp 1698175906
transform 1 0 19600 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _114_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 16240 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _115_
timestamp 1698175906
transform 1 0 14784 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _116_
timestamp 1698175906
transform 1 0 16576 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _117_
timestamp 1698175906
transform -1 0 19376 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _118_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18816 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _119_
timestamp 1698175906
transform 1 0 16576 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _120_
timestamp 1698175906
transform 1 0 18368 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _121_
timestamp 1698175906
transform 1 0 17360 0 -1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _122_
timestamp 1698175906
transform 1 0 15456 0 -1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _123_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16128 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _124_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19488 0 1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor3_2  _125_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 19488 0 -1 18816
box -86 -86 1654 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _126_
timestamp 1698175906
transform 1 0 18592 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _127_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 22064 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _128_
timestamp 1698175906
transform -1 0 22736 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _129_
timestamp 1698175906
transform -1 0 18592 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _130_
timestamp 1698175906
transform 1 0 17360 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _131_
timestamp 1698175906
transform -1 0 17920 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _132_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 14000 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _133_
timestamp 1698175906
transform 1 0 16800 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _134_
timestamp 1698175906
transform 1 0 18032 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _135_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16128 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _136_
timestamp 1698175906
transform 1 0 16688 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _137_
timestamp 1698175906
transform -1 0 18704 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _138_
timestamp 1698175906
transform -1 0 14560 0 1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _139_
timestamp 1698175906
transform 1 0 19824 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _140_
timestamp 1698175906
transform 1 0 20160 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _141_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 19488 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _142_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21392 0 -1 26656
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _143_
timestamp 1698175906
transform 1 0 25984 0 1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _144_
timestamp 1698175906
transform -1 0 27888 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _145_
timestamp 1698175906
transform -1 0 26544 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _146_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 15456 0 1 17248
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _147_
timestamp 1698175906
transform -1 0 15008 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _148_
timestamp 1698175906
transform 1 0 19376 0 -1 23520
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _149_
timestamp 1698175906
transform 1 0 20272 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _150_
timestamp 1698175906
transform 1 0 15120 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _151_
timestamp 1698175906
transform -1 0 21952 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _152_
timestamp 1698175906
transform 1 0 20496 0 -1 20384
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _153_
timestamp 1698175906
transform 1 0 20048 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _154_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18928 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _155_
timestamp 1698175906
transform -1 0 14896 0 1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _156_
timestamp 1698175906
transform -1 0 19152 0 1 21952
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _157_
timestamp 1698175906
transform 1 0 21168 0 1 26656
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _158_
timestamp 1698175906
transform 1 0 18368 0 1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _159_
timestamp 1698175906
transform 1 0 19600 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _160_
timestamp 1698175906
transform -1 0 21616 0 -1 23520
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _161_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20160 0 -1 26656
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_2  _162_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18480 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _163_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 17584 0 1 26656
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _164_
timestamp 1698175906
transform -1 0 16240 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _165_
timestamp 1698175906
transform 1 0 17472 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _166_
timestamp 1698175906
transform -1 0 18592 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _167_
timestamp 1698175906
transform -1 0 15120 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _168_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13440 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _169_
timestamp 1698175906
transform 1 0 20272 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _170_
timestamp 1698175906
transform 1 0 21168 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _171_
timestamp 1698175906
transform -1 0 23968 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _172_
timestamp 1698175906
transform -1 0 24304 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _173_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 22176 0 -1 18816
box -86 -86 1430 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _174_
timestamp 1698175906
transform 1 0 18032 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _175_
timestamp 1698175906
transform 1 0 18928 0 -1 25088
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _176_
timestamp 1698175906
transform 1 0 17808 0 1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _177_
timestamp 1698175906
transform -1 0 20048 0 1 25088
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__nor4_1  _178_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 19600 0 -1 26656
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _179_
timestamp 1698175906
transform -1 0 18480 0 -1 28224
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _180_
timestamp 1698175906
transform -1 0 28112 0 -1 25088
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _181_
timestamp 1698175906
transform -1 0 27328 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _182_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21616 0 1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _183_
timestamp 1698175906
transform 1 0 19712 0 -1 20384
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_2  _184_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 21168 0 1 21952
box -86 -86 2102 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _185_
timestamp 1698175906
transform 1 0 22288 0 -1 20384
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _186_
timestamp 1698175906
transform 1 0 18928 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _187_
timestamp 1698175906
transform 1 0 24304 0 -1 18816
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _188_
timestamp 1698175906
transform 1 0 25088 0 1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _189_
timestamp 1698175906
transform -1 0 25312 0 1 18816
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _190_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 18928 0 -1 21952
box -86 -86 1542 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _191_
timestamp 1698175906
transform 1 0 28000 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _192_
timestamp 1698175906
transform -1 0 28000 0 1 21952
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _193_
timestamp 1698175906
transform 1 0 25312 0 -1 20384
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _194_
timestamp 1698175906
transform 1 0 25088 0 -1 21952
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _195_
timestamp 1698175906
transform 1 0 25312 0 1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _196_
timestamp 1698175906
transform 1 0 26096 0 1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _197_
timestamp 1698175906
transform 1 0 13664 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _198_
timestamp 1698175906
transform 1 0 14896 0 1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _199_
timestamp 1698175906
transform 1 0 23184 0 -1 26656
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _200_
timestamp 1698175906
transform -1 0 22400 0 1 25088
box -86 -86 1318 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _201_
timestamp 1698175906
transform 1 0 22624 0 -1 26656
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _202_
timestamp 1698175906
transform 1 0 18480 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _203_
timestamp 1698175906
transform -1 0 17920 0 1 17248
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _204_
timestamp 1698175906
transform -1 0 22064 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _205_
timestamp 1698175906
transform 1 0 23072 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _206_
timestamp 1698175906
transform 1 0 22176 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _207_
timestamp 1698175906
transform 1 0 15344 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _208_
timestamp 1698175906
transform 1 0 16016 0 -1 15680
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _209_
timestamp 1698175906
transform -1 0 20832 0 1 12544
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _210_
timestamp 1698175906
transform 1 0 15232 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand4_2  _211_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17360 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _212_
timestamp 1698175906
transform 1 0 19376 0 1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _213_
timestamp 1698175906
transform -1 0 28672 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__aoi211_1  _214_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 22176 0 -1 18816
box -86 -86 1206 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _215_
timestamp 1698175906
transform 1 0 26432 0 1 17248
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _216_
timestamp 1698175906
transform -1 0 27216 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _217_
timestamp 1698175906
transform 1 0 23520 0 -1 18816
box -86 -86 870 870
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _218_
timestamp 1698175906
transform -1 0 26320 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _219_
timestamp 1698175906
transform 1 0 21056 0 -1 14112
box -86 -86 646 870
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _220_
timestamp 1698175906
transform 1 0 19488 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _221_
timestamp 1698175906
transform 1 0 21168 0 1 14112
box -86 -86 1094 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _222_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16128 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _223_
timestamp 1698175906
transform -1 0 14112 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _224_
timestamp 1698175906
transform 1 0 25312 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _225_
timestamp 1698175906
transform 1 0 11984 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _226_
timestamp 1698175906
transform 1 0 11984 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _227_
timestamp 1698175906
transform 1 0 11088 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _228_
timestamp 1698175906
transform 1 0 13328 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _229_
timestamp 1698175906
transform 1 0 19936 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _230_
timestamp 1698175906
transform 1 0 13776 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _231_
timestamp 1698175906
transform -1 0 14560 0 -1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _232_
timestamp 1698175906
transform 1 0 21840 0 1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _233_
timestamp 1698175906
transform 1 0 16464 0 1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _234_
timestamp 1698175906
transform 1 0 25536 0 1 25088
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _235_
timestamp 1698175906
transform 1 0 21616 0 -1 23520
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _236_
timestamp 1698175906
transform 1 0 25088 0 -1 18816
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _237_
timestamp 1698175906
transform 1 0 26880 0 -1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _238_
timestamp 1698175906
transform 1 0 23744 0 1 21952
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _239_
timestamp 1698175906
transform 1 0 26096 0 -1 20384
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _240_
timestamp 1698175906
transform 1 0 10528 0 -1 28224
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _241_
timestamp 1698175906
transform 1 0 22512 0 1 26656
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _242_
timestamp 1698175906
transform 1 0 21616 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _243_
timestamp 1698175906
transform 1 0 12992 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _244_
timestamp 1698175906
transform 1 0 17360 0 -1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _245_
timestamp 1698175906
transform 1 0 26432 0 -1 17248
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _246_
timestamp 1698175906
transform 1 0 24752 0 1 14112
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _247_
timestamp 1698175906
transform 1 0 21168 0 1 12544
box -86 -86 3334 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _249_
timestamp 1698175906
transform -1 0 14896 0 1 26656
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _250_
timestamp 1698175906
transform 1 0 29120 0 1 21952
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _251_
timestamp 1698175906
transform 1 0 25088 0 -1 14112
box -86 -86 758 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__182__C dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 21616 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__222__CLK
timestamp 1698175906
transform 1 0 20608 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__223__CLK
timestamp 1698175906
transform 1 0 14336 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__224__CLK
timestamp 1698175906
transform 1 0 28784 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__225__CLK
timestamp 1698175906
transform 1 0 15232 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__226__CLK
timestamp 1698175906
transform 1 0 15456 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__227__CLK
timestamp 1698175906
transform 1 0 14560 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__228__CLK
timestamp 1698175906
transform 1 0 16576 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__229__CLK
timestamp 1698175906
transform -1 0 23632 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__230__CLK
timestamp 1698175906
transform 1 0 17472 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__231__CLK
timestamp 1698175906
transform 1 0 15344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__232__CLK
timestamp 1698175906
transform 1 0 25312 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__233__CLK
timestamp 1698175906
transform 1 0 19936 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__234__CLK
timestamp 1698175906
transform 1 0 29232 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__235__CLK
timestamp 1698175906
transform 1 0 25312 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__236__CLK
timestamp 1698175906
transform 1 0 28560 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__237__CLK
timestamp 1698175906
transform 1 0 26656 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__238__CLK
timestamp 1698175906
transform 1 0 27216 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__239__CLK
timestamp 1698175906
transform 1 0 29568 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__240__CLK
timestamp 1698175906
transform 1 0 13776 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__241__CLK
timestamp 1698175906
transform 1 0 25984 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__242__CLK
timestamp 1698175906
transform -1 0 25088 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__243__CLK
timestamp 1698175906
transform -1 0 16464 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__244__CLK
timestamp 1698175906
transform 1 0 16800 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__245__CLK
timestamp 1698175906
transform 1 0 26208 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__246__CLK
timestamp 1698175906
transform 1 0 28224 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__247__CLK
timestamp 1698175906
transform -1 0 25536 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform 1 0 20720 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_output10_I
timestamp 1698175906
transform 1 0 37296 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 18928 0 -1 21952
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform -1 0 20944 0 1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 22736 0 1 20384
box -86 -86 5686 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 5376 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 9184 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 12992 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 16800 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 17248 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_172
timestamp 1698175906
transform 1 0 20608 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_176
timestamp 1698175906
transform 1 0 21056 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_232
timestamp 1698175906
transform 1 0 27328 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_236
timestamp 1698175906
transform 1 0 27776 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 28224 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 32032 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 35840 0 1 3136
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 39648 0 1 3136
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 40096 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 40320 0 1 3136
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1568 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 8736 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 9408 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 16576 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_168
timestamp 1698175906
transform 1 0 20160 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_195 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 23184 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_203
timestamp 1698175906
transform 1 0 24080 0 -1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_207
timestamp 1698175906
transform 1 0 24528 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_209
timestamp 1698175906
transform 1 0 24752 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_238
timestamp 1698175906
transform 1 0 28000 0 -1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_270
timestamp 1698175906
transform 1 0 31584 0 -1 4704
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_278
timestamp 1698175906
transform 1 0 32480 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 32928 0 -1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 40096 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 40320 0 -1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 1568 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 5152 0 1 4704
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 5488 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 12656 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 13328 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 20496 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_177
timestamp 1698175906
transform 1 0 21168 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 28336 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 29008 0 1 4704
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 36176 0 1 4704
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 36848 0 1 4704
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 1568 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 8736 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 9408 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 16576 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 17248 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 24416 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 25088 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 32256 0 -1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 32928 0 -1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 40096 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 40320 0 -1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 1568 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 5152 0 1 6272
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 5488 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 12656 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 13328 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 20496 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 21168 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 28336 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 29008 0 1 6272
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 36176 0 1 6272
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 36848 0 1 6272
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 1568 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 8736 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 9408 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 16576 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 17248 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 24416 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 25088 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 32256 0 -1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 32928 0 -1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 40096 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 40320 0 -1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 1568 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 5152 0 1 7840
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 5488 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 12656 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 13328 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 20496 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 21168 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 28336 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 29008 0 1 7840
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 36176 0 1 7840
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 36848 0 1 7840
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 1568 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 8736 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 9408 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 16576 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 17248 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 24416 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 25088 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 32256 0 -1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 32928 0 -1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 40096 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 40320 0 -1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 1568 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 5152 0 1 9408
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 5488 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 12656 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 13328 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 20496 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 21168 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 28336 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 29008 0 1 9408
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 36176 0 1 9408
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 36848 0 1 9408
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 1568 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 8736 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 9408 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 16576 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 17248 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 24416 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 25088 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 32256 0 -1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 32928 0 -1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 40096 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 40320 0 -1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 1568 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 5152 0 1 10976
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 5488 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 12656 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 13328 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 20496 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 21168 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 28336 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 29008 0 1 10976
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 36176 0 1 10976
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 36848 0 1 10976
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 1568 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 8736 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 9408 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 16576 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 17248 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 24416 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 25088 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 32256 0 -1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 32928 0 -1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 40096 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 40320 0 -1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 1568 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 5152 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 5488 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 12656 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_107 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13328 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_123
timestamp 1698175906
transform 1 0 15120 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_131
timestamp 1698175906
transform 1 0 16016 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_135
timestamp 1698175906
transform 1 0 16464 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_167
timestamp 1698175906
transform 1 0 20048 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_174
timestamp 1698175906
transform 1 0 20832 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_206
timestamp 1698175906
transform 1 0 24416 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_212
timestamp 1698175906
transform 1 0 25088 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_216
timestamp 1698175906
transform 1 0 25536 0 1 12544
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_12_232
timestamp 1698175906
transform 1 0 27328 0 1 12544
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_240
timestamp 1698175906
transform 1 0 28224 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_244
timestamp 1698175906
transform 1 0 28672 0 1 12544
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 29008 0 1 12544
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 36176 0 1 12544
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 36848 0 1 12544
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 1568 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 8736 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_72
timestamp 1698175906
transform 1 0 9408 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_133
timestamp 1698175906
transform 1 0 16240 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_137
timestamp 1698175906
transform 1 0 16688 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_142
timestamp 1698175906
transform 1 0 17248 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_172
timestamp 1698175906
transform 1 0 20608 0 -1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_13_218
timestamp 1698175906
transform 1 0 25760 0 -1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_226
timestamp 1698175906
transform 1 0 26656 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_231
timestamp 1698175906
transform 1 0 27216 0 -1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_13_263
timestamp 1698175906
transform 1 0 30800 0 -1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_279
timestamp 1698175906
transform 1 0 32592 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 32928 0 -1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 40096 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 40320 0 -1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 1568 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 5152 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 5488 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 12656 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_107
timestamp 1698175906
transform 1 0 13328 0 1 14112
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_123
timestamp 1698175906
transform 1 0 15120 0 1 14112
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_131
timestamp 1698175906
transform 1 0 16016 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_170
timestamp 1698175906
transform 1 0 20384 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_174
timestamp 1698175906
transform 1 0 20832 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_202
timestamp 1698175906
transform 1 0 23968 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_206
timestamp 1698175906
transform 1 0 24416 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_208
timestamp 1698175906
transform 1 0 24640 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_238
timestamp 1698175906
transform 1 0 28000 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_242
timestamp 1698175906
transform 1 0 28448 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_244
timestamp 1698175906
transform 1 0 28672 0 1 14112
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 29008 0 1 14112
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 36176 0 1 14112
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 36848 0 1 14112
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 1568 0 -1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 8736 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_72
timestamp 1698175906
transform 1 0 9408 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_104
timestamp 1698175906
transform 1 0 12992 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_120
timestamp 1698175906
transform 1 0 14784 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_124
timestamp 1698175906
transform 1 0 15232 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_137
timestamp 1698175906
transform 1 0 16688 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_139
timestamp 1698175906
transform 1 0 16912 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_142
timestamp 1698175906
transform 1 0 17248 0 -1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_146
timestamp 1698175906
transform 1 0 17696 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_170
timestamp 1698175906
transform 1 0 20384 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_178
timestamp 1698175906
transform 1 0 21280 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_180
timestamp 1698175906
transform 1 0 21504 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_191
timestamp 1698175906
transform 1 0 22736 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_207
timestamp 1698175906
transform 1 0 24528 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_209
timestamp 1698175906
transform 1 0 24752 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_212
timestamp 1698175906
transform 1 0 25088 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_214
timestamp 1698175906
transform 1 0 25312 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_223
timestamp 1698175906
transform 1 0 26320 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_255
timestamp 1698175906
transform 1 0 29904 0 -1 15680
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_271
timestamp 1698175906
transform 1 0 31696 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_279
timestamp 1698175906
transform 1 0 32592 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_282
timestamp 1698175906
transform 1 0 32928 0 -1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_314
timestamp 1698175906
transform 1 0 36512 0 -1 15680
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_322
timestamp 1698175906
transform 1 0 37408 0 -1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 1568 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 5152 0 1 15680
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 5488 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 12656 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_107
timestamp 1698175906
transform 1 0 13328 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_171
timestamp 1698175906
transform 1 0 20496 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_177
timestamp 1698175906
transform 1 0 21168 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_241
timestamp 1698175906
transform 1 0 28336 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 29008 0 1 15680
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 36176 0 1 15680
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_317
timestamp 1698175906
transform 1 0 36848 0 1 15680
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_2
timestamp 1698175906
transform 1 0 1568 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_66
timestamp 1698175906
transform 1 0 8736 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_72
timestamp 1698175906
transform 1 0 9408 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_88
timestamp 1698175906
transform 1 0 11200 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_92
timestamp 1698175906
transform 1 0 11648 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_94
timestamp 1698175906
transform 1 0 11872 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_124
timestamp 1698175906
transform 1 0 15232 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_128
timestamp 1698175906
transform 1 0 15680 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_136
timestamp 1698175906
transform 1 0 16576 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_142
timestamp 1698175906
transform 1 0 17248 0 -1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_174
timestamp 1698175906
transform 1 0 20832 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_190
timestamp 1698175906
transform 1 0 22624 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_198
timestamp 1698175906
transform 1 0 23520 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_200
timestamp 1698175906
transform 1 0 23744 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_205
timestamp 1698175906
transform 1 0 24304 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1698175906
transform 1 0 24752 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_212
timestamp 1698175906
transform 1 0 25088 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_216
timestamp 1698175906
transform 1 0 25536 0 -1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_220
timestamp 1698175906
transform 1 0 25984 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_17_253
timestamp 1698175906
transform 1 0 29680 0 -1 17248
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_269
timestamp 1698175906
transform 1 0 31472 0 -1 17248
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_277
timestamp 1698175906
transform 1 0 32368 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_279
timestamp 1698175906
transform 1 0 32592 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_17_282
timestamp 1698175906
transform 1 0 32928 0 -1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_346
timestamp 1698175906
transform 1 0 40096 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_348
timestamp 1698175906
transform 1 0 40320 0 -1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_2
timestamp 1698175906
transform 1 0 1568 0 1 17248
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 5152 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698175906
transform 1 0 5488 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698175906
transform 1 0 12656 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_107
timestamp 1698175906
transform 1 0 13328 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_111
timestamp 1698175906
transform 1 0 13776 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_113
timestamp 1698175906
transform 1 0 14000 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_132
timestamp 1698175906
transform 1 0 16128 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_148
timestamp 1698175906
transform 1 0 17920 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_164
timestamp 1698175906
transform 1 0 19712 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_171
timestamp 1698175906
transform 1 0 20496 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_177
timestamp 1698175906
transform 1 0 21168 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_181
timestamp 1698175906
transform 1 0 21616 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_220
timestamp 1698175906
transform 1 0 25984 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_233
timestamp 1698175906
transform 1 0 27440 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_237
timestamp 1698175906
transform 1 0 27888 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_239
timestamp 1698175906
transform 1 0 28112 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_244
timestamp 1698175906
transform 1 0 28672 0 1 17248
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698175906
transform 1 0 29008 0 1 17248
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698175906
transform 1 0 36176 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_317
timestamp 1698175906
transform 1 0 36848 0 1 17248
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_321
timestamp 1698175906
transform 1 0 37296 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698175906
transform 1 0 1568 0 -1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698175906
transform 1 0 8736 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_72
timestamp 1698175906
transform 1 0 9408 0 -1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_88
timestamp 1698175906
transform 1 0 11200 0 -1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_92
timestamp 1698175906
transform 1 0 11648 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_94
timestamp 1698175906
transform 1 0 11872 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_142
timestamp 1698175906
transform 1 0 17248 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_241
timestamp 1698175906
transform 1 0 28336 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_245
timestamp 1698175906
transform 1 0 28784 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_277
timestamp 1698175906
transform 1 0 32368 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_279
timestamp 1698175906
transform 1 0 32592 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_19_282
timestamp 1698175906
transform 1 0 32928 0 -1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_314
timestamp 1698175906
transform 1 0 36512 0 -1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_322
timestamp 1698175906
transform 1 0 37408 0 -1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 1568 0 1 18816
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 5152 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_37
timestamp 1698175906
transform 1 0 5488 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_101
timestamp 1698175906
transform 1 0 12656 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_107
timestamp 1698175906
transform 1 0 13328 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_115
timestamp 1698175906
transform 1 0 14224 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_122
timestamp 1698175906
transform 1 0 15008 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_126
timestamp 1698175906
transform 1 0 15456 0 1 18816
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_134
timestamp 1698175906
transform 1 0 16352 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_136
timestamp 1698175906
transform 1 0 16576 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_183
timestamp 1698175906
transform 1 0 21840 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_191
timestamp 1698175906
transform 1 0 22736 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_207
timestamp 1698175906
transform 1 0 24528 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_228
timestamp 1698175906
transform 1 0 26880 0 1 18816
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_244
timestamp 1698175906
transform 1 0 28672 0 1 18816
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_20_247
timestamp 1698175906
transform 1 0 29008 0 1 18816
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_311
timestamp 1698175906
transform 1 0 36176 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_317
timestamp 1698175906
transform 1 0 36848 0 1 18816
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_321
timestamp 1698175906
transform 1 0 37296 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_2
timestamp 1698175906
transform 1 0 1568 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_66
timestamp 1698175906
transform 1 0 8736 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_21_72
timestamp 1698175906
transform 1 0 9408 0 -1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_136
timestamp 1698175906
transform 1 0 16576 0 -1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_142
timestamp 1698175906
transform 1 0 17248 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_161
timestamp 1698175906
transform 1 0 19376 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_163
timestamp 1698175906
transform 1 0 19600 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_169
timestamp 1698175906
transform 1 0 20272 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_177
timestamp 1698175906
transform 1 0 21168 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_184
timestamp 1698175906
transform 1 0 21952 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_186
timestamp 1698175906
transform 1 0 22176 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_202
timestamp 1698175906
transform 1 0 23968 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_212
timestamp 1698175906
transform 1 0 25088 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_250
timestamp 1698175906
transform 1 0 29344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_254
timestamp 1698175906
transform 1 0 29792 0 -1 20384
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_270
timestamp 1698175906
transform 1 0 31584 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_278
timestamp 1698175906
transform 1 0 32480 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_282
timestamp 1698175906
transform 1 0 32928 0 -1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_314
timestamp 1698175906
transform 1 0 36512 0 -1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_322
timestamp 1698175906
transform 1 0 37408 0 -1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 1568 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 5152 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698175906
transform 1 0 5488 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698175906
transform 1 0 12656 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_107
timestamp 1698175906
transform 1 0 13328 0 1 20384
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_115
timestamp 1698175906
transform 1 0 14224 0 1 20384
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_121
timestamp 1698175906
transform 1 0 14896 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_177
timestamp 1698175906
transform 1 0 21168 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_241
timestamp 1698175906
transform 1 0 28336 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698175906
transform 1 0 29008 0 1 20384
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698175906
transform 1 0 36176 0 1 20384
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_317
timestamp 1698175906
transform 1 0 36848 0 1 20384
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698175906
transform 1 0 1568 0 -1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698175906
transform 1 0 8736 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_72
timestamp 1698175906
transform 1 0 9408 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_80
timestamp 1698175906
transform 1 0 10304 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_84
timestamp 1698175906
transform 1 0 10752 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_86
timestamp 1698175906
transform 1 0 10976 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_116
timestamp 1698175906
transform 1 0 14336 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_142
timestamp 1698175906
transform 1 0 17248 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_207
timestamp 1698175906
transform 1 0 24528 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_209
timestamp 1698175906
transform 1 0 24752 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_222
timestamp 1698175906
transform 1 0 26208 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_257
timestamp 1698175906
transform 1 0 30128 0 -1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_273
timestamp 1698175906
transform 1 0 31920 0 -1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_277
timestamp 1698175906
transform 1 0 32368 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_279
timestamp 1698175906
transform 1 0 32592 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_23_282
timestamp 1698175906
transform 1 0 32928 0 -1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_314
timestamp 1698175906
transform 1 0 36512 0 -1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_322
timestamp 1698175906
transform 1 0 37408 0 -1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698175906
transform 1 0 1568 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 5152 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698175906
transform 1 0 5488 0 1 21952
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698175906
transform 1 0 12656 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_136
timestamp 1698175906
transform 1 0 16576 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_159
timestamp 1698175906
transform 1 0 19152 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_161
timestamp 1698175906
transform 1 0 19376 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_171
timestamp 1698175906
transform 1 0 20496 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_195
timestamp 1698175906
transform 1 0 23184 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_199
timestamp 1698175906
transform 1 0 23632 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_229
timestamp 1698175906
transform 1 0 26992 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_243
timestamp 1698175906
transform 1 0 28560 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_247
timestamp 1698175906
transform 1 0 29008 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_254
timestamp 1698175906
transform 1 0 29792 0 1 21952
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_286
timestamp 1698175906
transform 1 0 33376 0 1 21952
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_302
timestamp 1698175906
transform 1 0 35168 0 1 21952
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_310
timestamp 1698175906
transform 1 0 36064 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_314
timestamp 1698175906
transform 1 0 36512 0 1 21952
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_317
timestamp 1698175906
transform 1 0 36848 0 1 21952
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698175906
transform 1 0 37296 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2
timestamp 1698175906
transform 1 0 1568 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_66
timestamp 1698175906
transform 1 0 8736 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_72
timestamp 1698175906
transform 1 0 9408 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_80
timestamp 1698175906
transform 1 0 10304 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_84
timestamp 1698175906
transform 1 0 10752 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_114
timestamp 1698175906
transform 1 0 14112 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_118
timestamp 1698175906
transform 1 0 14560 0 -1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_122
timestamp 1698175906
transform 1 0 15008 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_133
timestamp 1698175906
transform 1 0 16240 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_135
timestamp 1698175906
transform 1 0 16464 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_142
timestamp 1698175906
transform 1 0 17248 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_166
timestamp 1698175906
transform 1 0 19936 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_212
timestamp 1698175906
transform 1 0 25088 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_216
timestamp 1698175906
transform 1 0 25536 0 -1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_282
timestamp 1698175906
transform 1 0 32928 0 -1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_314
timestamp 1698175906
transform 1 0 36512 0 -1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_322
timestamp 1698175906
transform 1 0 37408 0 -1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_28
timestamp 1698175906
transform 1 0 4480 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_32
timestamp 1698175906
transform 1 0 4928 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 5152 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698175906
transform 1 0 5488 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698175906
transform 1 0 12656 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_107
timestamp 1698175906
transform 1 0 13328 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_118
timestamp 1698175906
transform 1 0 14560 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_134
timestamp 1698175906
transform 1 0 16352 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_138
timestamp 1698175906
transform 1 0 16800 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_146
timestamp 1698175906
transform 1 0 17696 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_155
timestamp 1698175906
transform 1 0 18704 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_171
timestamp 1698175906
transform 1 0 20496 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_177
timestamp 1698175906
transform 1 0 21168 0 1 23520
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_209
timestamp 1698175906
transform 1 0 24752 0 1 23520
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_217
timestamp 1698175906
transform 1 0 25648 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_219
timestamp 1698175906
transform 1 0 25872 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_26_226
timestamp 1698175906
transform 1 0 26656 0 1 23520
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_242
timestamp 1698175906
transform 1 0 28448 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_244
timestamp 1698175906
transform 1 0 28672 0 1 23520
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 29008 0 1 23520
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 36176 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_317
timestamp 1698175906
transform 1 0 36848 0 1 23520
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698175906
transform 1 0 1568 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698175906
transform 1 0 8736 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_72
timestamp 1698175906
transform 1 0 9408 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_136
timestamp 1698175906
transform 1 0 16576 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_148
timestamp 1698175906
transform 1 0 17920 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_154
timestamp 1698175906
transform 1 0 18592 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_156
timestamp 1698175906
transform 1 0 18816 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_163
timestamp 1698175906
transform 1 0 19600 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_167
timestamp 1698175906
transform 1 0 20048 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_174
timestamp 1698175906
transform 1 0 20832 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_206
timestamp 1698175906
transform 1 0 24416 0 -1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_212
timestamp 1698175906
transform 1 0 25088 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_225
timestamp 1698175906
transform 1 0 26544 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_233
timestamp 1698175906
transform 1 0 27440 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_239
timestamp 1698175906
transform 1 0 28112 0 -1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_271
timestamp 1698175906
transform 1 0 31696 0 -1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_279
timestamp 1698175906
transform 1 0 32592 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_282
timestamp 1698175906
transform 1 0 32928 0 -1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_346
timestamp 1698175906
transform 1 0 40096 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_348
timestamp 1698175906
transform 1 0 40320 0 -1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698175906
transform 1 0 1568 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 5152 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 5488 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 12656 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_107
timestamp 1698175906
transform 1 0 13328 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_116
timestamp 1698175906
transform 1 0 14336 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_132
timestamp 1698175906
transform 1 0 16128 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_140
timestamp 1698175906
transform 1 0 17024 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_144
timestamp 1698175906
transform 1 0 17472 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_146
timestamp 1698175906
transform 1 0 17696 0 1 25088
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_167
timestamp 1698175906
transform 1 0 20048 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_188
timestamp 1698175906
transform 1 0 22400 0 1 25088
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_204
timestamp 1698175906
transform 1 0 24192 0 1 25088
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_212
timestamp 1698175906
transform 1 0 25088 0 1 25088
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_247
timestamp 1698175906
transform 1 0 29008 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_251
timestamp 1698175906
transform 1 0 29456 0 1 25088
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_317
timestamp 1698175906
transform 1 0 36848 0 1 25088
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2
timestamp 1698175906
transform 1 0 1568 0 -1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_66
timestamp 1698175906
transform 1 0 8736 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_72
timestamp 1698175906
transform 1 0 9408 0 -1 26656
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_88
timestamp 1698175906
transform 1 0 11200 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_123
timestamp 1698175906
transform 1 0 15120 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_127
timestamp 1698175906
transform 1 0 15568 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_135
timestamp 1698175906
transform 1 0 16464 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_139
timestamp 1698175906
transform 1 0 16912 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_142
timestamp 1698175906
transform 1 0 17248 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_146
timestamp 1698175906
transform 1 0 17696 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_148
timestamp 1698175906
transform 1 0 17920 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_186
timestamp 1698175906
transform 1 0 22176 0 -1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_202
timestamp 1698175906
transform 1 0 23968 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_212
timestamp 1698175906
transform 1 0 25088 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_243
timestamp 1698175906
transform 1 0 28560 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_247
timestamp 1698175906
transform 1 0 29008 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_279
timestamp 1698175906
transform 1 0 32592 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_282
timestamp 1698175906
transform 1 0 32928 0 -1 26656
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_314
timestamp 1698175906
transform 1 0 36512 0 -1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_322
timestamp 1698175906
transform 1 0 37408 0 -1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_28
timestamp 1698175906
transform 1 0 4480 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_32
timestamp 1698175906
transform 1 0 4928 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 5152 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 5488 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 12656 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_107
timestamp 1698175906
transform 1 0 13328 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_109
timestamp 1698175906
transform 1 0 13552 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_126
timestamp 1698175906
transform 1 0 15456 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_128
timestamp 1698175906
transform 1 0 15680 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_133
timestamp 1698175906
transform 1 0 16240 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_135
timestamp 1698175906
transform 1 0 16464 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_145
timestamp 1698175906
transform 1 0 17584 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_153
timestamp 1698175906
transform 1 0 18480 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_155
timestamp 1698175906
transform 1 0 18704 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_162
timestamp 1698175906
transform 1 0 19488 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_170
timestamp 1698175906
transform 1 0 20384 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_174
timestamp 1698175906
transform 1 0 20832 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_184
timestamp 1698175906
transform 1 0 21952 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_188
timestamp 1698175906
transform 1 0 22400 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_218
timestamp 1698175906
transform 1 0 25760 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_222
timestamp 1698175906
transform 1 0 26208 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_226
timestamp 1698175906
transform 1 0 26656 0 1 26656
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_237
timestamp 1698175906
transform 1 0 27888 0 1 26656
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 29008 0 1 26656
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 36176 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_317
timestamp 1698175906
transform 1 0 36848 0 1 26656
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_321
timestamp 1698175906
transform 1 0 37296 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 1568 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 8736 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_72
timestamp 1698175906
transform 1 0 9408 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_80
timestamp 1698175906
transform 1 0 10304 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_142
timestamp 1698175906
transform 1 0 17248 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_146
timestamp 1698175906
transform 1 0 17696 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_153
timestamp 1698175906
transform 1 0 18480 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_161
timestamp 1698175906
transform 1 0 19376 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_165
timestamp 1698175906
transform 1 0 19824 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_195
timestamp 1698175906
transform 1 0 23184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_31_199
timestamp 1698175906
transform 1 0 23632 0 -1 28224
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_207
timestamp 1698175906
transform 1 0 24528 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_209
timestamp 1698175906
transform 1 0 24752 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698175906
transform 1 0 25088 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698175906
transform 1 0 32256 0 -1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 32928 0 -1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 40096 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 40320 0 -1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 1568 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 5152 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 5488 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 12656 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_107
timestamp 1698175906
transform 1 0 13328 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_32_113
timestamp 1698175906
transform 1 0 14000 0 1 28224
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_129
timestamp 1698175906
transform 1 0 15792 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_133
timestamp 1698175906
transform 1 0 16240 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_164
timestamp 1698175906
transform 1 0 19712 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_168
timestamp 1698175906
transform 1 0 20160 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_32_172
timestamp 1698175906
transform 1 0 20608 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_174
timestamp 1698175906
transform 1 0 20832 0 1 28224
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698175906
transform 1 0 21168 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698175906
transform 1 0 28336 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 29008 0 1 28224
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 36176 0 1 28224
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 36848 0 1 28224
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 1568 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 8736 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 9408 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 16576 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_142
timestamp 1698175906
transform 1 0 17248 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_206
timestamp 1698175906
transform 1 0 24416 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 25088 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 32256 0 -1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 32928 0 -1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 40096 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 40320 0 -1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 1568 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 5152 0 1 29792
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 5488 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 12656 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 13328 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 20496 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 21168 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 28336 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 29008 0 1 29792
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 36176 0 1 29792
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 36848 0 1 29792
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 1568 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 8736 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 9408 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 16576 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 17248 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 24416 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 25088 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 32256 0 -1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 32928 0 -1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 40096 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 40320 0 -1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 1568 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 5152 0 1 31360
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 5488 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 12656 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 13328 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 20496 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 21168 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 28336 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 29008 0 1 31360
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 36176 0 1 31360
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 36848 0 1 31360
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 1568 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 8736 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 9408 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 16576 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 17248 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 24416 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 25088 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 32256 0 -1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 32928 0 -1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 40096 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 40320 0 -1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 1568 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 5152 0 1 32928
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 5488 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 12656 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 13328 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 20496 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 21168 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 28336 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 29008 0 1 32928
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 36176 0 1 32928
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 36848 0 1 32928
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 1568 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 8736 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 9408 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 16576 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 17248 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 24416 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 25088 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 32256 0 -1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 32928 0 -1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 40096 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 40320 0 -1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 1568 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 5152 0 1 34496
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 5488 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 12656 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 13328 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 20496 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 21168 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 28336 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 29008 0 1 34496
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 36176 0 1 34496
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 36848 0 1 34496
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 1568 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 8736 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 9408 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 16576 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 17248 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 24416 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 25088 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 32256 0 -1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 32928 0 -1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 40096 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 40320 0 -1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 1568 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 5152 0 1 36064
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 5488 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 12656 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_107
timestamp 1698175906
transform 1 0 13328 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_171
timestamp 1698175906
transform 1 0 20496 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698175906
transform 1 0 21168 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 28336 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 29008 0 1 36064
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 36176 0 1 36064
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 36848 0 1 36064
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 1568 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 8736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_72
timestamp 1698175906
transform 1 0 9408 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_104
timestamp 1698175906
transform 1 0 12992 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_112
timestamp 1698175906
transform 1 0 13888 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_142
timestamp 1698175906
transform 1 0 17248 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_174
timestamp 1698175906
transform 1 0 20832 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_182
timestamp 1698175906
transform 1 0 21728 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_186
timestamp 1698175906
transform 1 0 22176 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_43_191
timestamp 1698175906
transform 1 0 22736 0 -1 37632
box -86 -86 1878 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_207
timestamp 1698175906
transform 1 0 24528 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 24752 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_43_238
timestamp 1698175906
transform 1 0 28000 0 -1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_270
timestamp 1698175906
transform 1 0 31584 0 -1 37632
box -86 -86 982 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_278
timestamp 1698175906
transform 1 0 32480 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 32928 0 -1 37632
box -86 -86 7254 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 40096 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 40320 0 -1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 1568 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 5376 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 9184 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_104
timestamp 1698175906
transform 1 0 12992 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_108
timestamp 1698175906
transform 1 0 13440 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_138
timestamp 1698175906
transform 1 0 16800 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_142
timestamp 1698175906
transform 1 0 17248 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_198
timestamp 1698175906
transform 1 0 23520 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_202
timestamp 1698175906
transform 1 0 23968 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_232
timestamp 1698175906
transform 1 0 27328 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_236
timestamp 1698175906
transform 1 0 27776 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_240
timestamp 1698175906
transform 1 0 28224 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 32032 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 35840 0 1 37632
box -86 -86 3670 870
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 39648 0 1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 40096 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 40320 0 1 37632
box -86 -86 198 870
use gf180mcu_fd_sc_mcu7t5v0__tiel  ita35_26 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 22736 0 -1 37632
box -86 -86 534 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 37520 0 1 17248
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform 1 0 37520 0 -1 15680
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform -1 0 24192 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform 1 0 25088 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform 1 0 37520 0 1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform 1 0 24416 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform 1 0 13664 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform 1 0 37520 0 1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform 1 0 14112 0 -1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform 1 0 37520 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform 1 0 37520 0 -1 21952
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform 1 0 37520 0 -1 20384
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform 1 0 20272 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform 1 0 37520 0 -1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform 1 0 25088 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform 1 0 17248 0 -1 4704
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform 1 0 20608 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform 1 0 37520 0 -1 18816
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform -1 0 4480 0 1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform 1 0 17472 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform 1 0 24416 0 1 37632
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform 1 0 37520 0 1 26656
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform -1 0 4480 0 1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698175906
transform 1 0 37520 0 -1 23520
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output25
timestamp 1698175906
transform 1 0 17472 0 1 3136
box -86 -86 2998 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 1344 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 40656 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 1344 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 40656 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 1344 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 40656 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 1344 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 40656 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 1344 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 40656 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 1344 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 40656 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 1344 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 40656 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 1344 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 40656 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 1344 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 40656 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 1344 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 40656 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 1344 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 40656 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 1344 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 40656 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 1344 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 40656 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 1344 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 40656 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 1344 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 40656 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 1344 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 40656 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 1344 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 40656 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 1344 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 40656 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 1344 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 40656 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 1344 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 40656 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 1344 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 40656 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 1344 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 40656 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 1344 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 40656 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 1344 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 40656 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 1344 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 40656 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 1344 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 40656 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 1344 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 40656 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 1344 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 40656 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 1344 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 40656 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 1344 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 40656 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 1344 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 40656 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 1344 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 40656 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 1344 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 40656 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 1344 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 40656 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 1344 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 40656 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 1344 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 40656 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 1344 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 40656 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 1344 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 40656 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 1344 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 40656 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 1344 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 40656 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 1344 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 40656 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 1344 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 40656 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 1344 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 40656 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 1344 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 40656 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 1344 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 40656 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 5152 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 8960 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 12768 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 16576 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 20384 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 24192 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 28000 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 31808 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 35616 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 39424 0 1 3136
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 9184 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 17024 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 24864 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 32704 0 -1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 5264 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 13104 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 20944 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 28784 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 36624 0 1 4704
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 9184 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 17024 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 24864 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 32704 0 -1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 5264 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 13104 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 20944 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 28784 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 36624 0 1 6272
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 9184 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 17024 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 24864 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 32704 0 -1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 5264 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 13104 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 20944 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 28784 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 36624 0 1 7840
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 9184 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 17024 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 24864 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 32704 0 -1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 5264 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 13104 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 20944 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 28784 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 36624 0 1 9408
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 9184 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 17024 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 24864 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 32704 0 -1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 5264 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 13104 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 20944 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 28784 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 36624 0 1 10976
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 9184 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 17024 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 24864 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 32704 0 -1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 5264 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 13104 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 20944 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 28784 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 36624 0 1 12544
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 9184 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 17024 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 24864 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 32704 0 -1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 5264 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 13104 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 20944 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 28784 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 36624 0 1 14112
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 9184 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 17024 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 24864 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 32704 0 -1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 5264 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 13104 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 20944 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 28784 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 36624 0 1 15680
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 9184 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 17024 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 24864 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 32704 0 -1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 5264 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 13104 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 20944 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 28784 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 36624 0 1 17248
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 9184 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 17024 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 24864 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 32704 0 -1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 5264 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 13104 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 20944 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 28784 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 36624 0 1 18816
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 9184 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 17024 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 24864 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 32704 0 -1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 5264 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 13104 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 20944 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 28784 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 36624 0 1 20384
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 9184 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 17024 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 24864 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 32704 0 -1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 5264 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 13104 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 20944 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 28784 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 36624 0 1 21952
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 9184 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 17024 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 24864 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 32704 0 -1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 5264 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 13104 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 20944 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 28784 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 36624 0 1 23520
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 9184 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 17024 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 24864 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 32704 0 -1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 5264 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 13104 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 20944 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 28784 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 36624 0 1 25088
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 9184 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 17024 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 24864 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 32704 0 -1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 5264 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 13104 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 20944 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 28784 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 36624 0 1 26656
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 9184 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 17024 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 24864 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 32704 0 -1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 5264 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 13104 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 20944 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 28784 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 36624 0 1 28224
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 9184 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 17024 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 24864 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 32704 0 -1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 5264 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 13104 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 20944 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 28784 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 36624 0 1 29792
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 9184 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 17024 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 24864 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 32704 0 -1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 5264 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 13104 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 20944 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 28784 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 36624 0 1 31360
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 9184 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 17024 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 24864 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 32704 0 -1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 5264 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 13104 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 20944 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 28784 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 36624 0 1 32928
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 9184 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 17024 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 24864 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 32704 0 -1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 5264 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 13104 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 20944 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 28784 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 36624 0 1 34496
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 9184 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 17024 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 24864 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 32704 0 -1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 5264 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 13104 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 20944 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 28784 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 36624 0 1 36064
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 9184 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 17024 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 24864 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 32704 0 -1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 5152 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 8960 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 12768 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 16576 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 20384 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 24192 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 28000 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 31808 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 35616 0 1 37632
box -86 -86 310 870
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 39424 0 1 37632
box -86 -86 310 870
<< labels >>
flabel metal3 s 0 27552 800 27664 0 FreeSans 448 0 0 0 clk
port 0 nsew signal input
flabel metal2 s 22176 41200 22288 42000 0 FreeSans 448 90 0 0 segm[0]
port 1 nsew signal tristate
flabel metal3 s 41200 17472 42000 17584 0 FreeSans 448 0 0 0 segm[10]
port 2 nsew signal tristate
flabel metal3 s 41200 14784 42000 14896 0 FreeSans 448 0 0 0 segm[11]
port 3 nsew signal tristate
flabel metal2 s 22176 0 22288 800 0 FreeSans 448 90 0 0 segm[12]
port 4 nsew signal tristate
flabel metal2 s 24864 41200 24976 42000 0 FreeSans 448 90 0 0 segm[13]
port 5 nsew signal tristate
flabel metal3 s 41200 18816 42000 18928 0 FreeSans 448 0 0 0 segm[1]
port 6 nsew signal tristate
flabel metal2 s 23520 0 23632 800 0 FreeSans 448 90 0 0 segm[2]
port 7 nsew signal tristate
flabel metal2 s 14784 41200 14896 42000 0 FreeSans 448 90 0 0 segm[3]
port 8 nsew signal tristate
flabel metal3 s 41200 22176 42000 22288 0 FreeSans 448 0 0 0 segm[4]
port 9 nsew signal tristate
flabel metal2 s 14112 41200 14224 42000 0 FreeSans 448 90 0 0 segm[5]
port 10 nsew signal tristate
flabel metal3 s 41200 23520 42000 23632 0 FreeSans 448 0 0 0 segm[6]
port 11 nsew signal tristate
flabel metal3 s 41200 21504 42000 21616 0 FreeSans 448 0 0 0 segm[7]
port 12 nsew signal tristate
flabel metal3 s 41200 19488 42000 19600 0 FreeSans 448 0 0 0 segm[8]
port 13 nsew signal tristate
flabel metal2 s 20160 0 20272 800 0 FreeSans 448 90 0 0 segm[9]
port 14 nsew signal tristate
flabel metal3 s 41200 25536 42000 25648 0 FreeSans 448 0 0 0 sel[0]
port 15 nsew signal tristate
flabel metal2 s 24864 0 24976 800 0 FreeSans 448 90 0 0 sel[10]
port 16 nsew signal tristate
flabel metal2 s 16128 0 16240 800 0 FreeSans 448 90 0 0 sel[11]
port 17 nsew signal tristate
flabel metal2 s 19488 41200 19600 42000 0 FreeSans 448 90 0 0 sel[1]
port 18 nsew signal tristate
flabel metal3 s 41200 18144 42000 18256 0 FreeSans 448 0 0 0 sel[2]
port 19 nsew signal tristate
flabel metal3 s 0 26208 800 26320 0 FreeSans 448 0 0 0 sel[3]
port 20 nsew signal tristate
flabel metal2 s 17472 41200 17584 42000 0 FreeSans 448 90 0 0 sel[4]
port 21 nsew signal tristate
flabel metal2 s 22848 41200 22960 42000 0 FreeSans 448 90 0 0 sel[5]
port 22 nsew signal tristate
flabel metal3 s 41200 26208 42000 26320 0 FreeSans 448 0 0 0 sel[6]
port 23 nsew signal tristate
flabel metal3 s 0 23520 800 23632 0 FreeSans 448 0 0 0 sel[7]
port 24 nsew signal tristate
flabel metal3 s 41200 22848 42000 22960 0 FreeSans 448 0 0 0 sel[8]
port 25 nsew signal tristate
flabel metal2 s 19488 0 19600 800 0 FreeSans 448 90 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 4448 3076 4768 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 35168 3076 35488 38476 0 FreeSans 1280 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 19808 3076 20128 38476 0 FreeSans 1280 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 21000 38416 21000 38416 0 vdd
rlabel metal1 21000 37632 21000 37632 0 vss
rlabel metal2 13664 25592 13664 25592 0 _000_
rlabel metal2 22792 17808 22792 17808 0 _001_
rlabel metal2 17976 27888 17976 27888 0 _002_
rlabel metal2 26824 26208 26824 26208 0 _003_
rlabel metal2 22512 23016 22512 23016 0 _004_
rlabel metal3 25536 18312 25536 18312 0 _005_
rlabel metal2 27832 21728 27832 21728 0 _006_
rlabel metal2 24696 21952 24696 21952 0 _007_
rlabel metal2 26824 19656 26824 19656 0 _008_
rlabel metal3 13328 27272 13328 27272 0 _009_
rlabel metal2 23128 26432 23128 26432 0 _010_
rlabel metal2 22568 14056 22568 14056 0 _011_
rlabel metal2 13944 14504 13944 14504 0 _012_
rlabel metal2 18312 14168 18312 14168 0 _013_
rlabel metal2 27384 17024 27384 17024 0 _014_
rlabel metal2 25704 14672 25704 14672 0 _015_
rlabel metal2 22120 13160 22120 13160 0 _016_
rlabel metal2 17080 14840 17080 14840 0 _017_
rlabel metal2 13160 23464 13160 23464 0 _018_
rlabel metal2 26040 25536 26040 25536 0 _019_
rlabel metal2 12936 18032 12936 18032 0 _020_
rlabel metal2 14504 17976 14504 17976 0 _021_
rlabel metal2 20328 22288 20328 22288 0 _022_
rlabel metal2 14392 21504 14392 21504 0 _023_
rlabel metal2 20832 27720 20832 27720 0 _024_
rlabel metal2 15960 27496 15960 27496 0 _025_
rlabel metal3 19544 25256 19544 25256 0 _026_
rlabel metal2 20160 26376 20160 26376 0 _027_
rlabel metal2 20664 26040 20664 26040 0 _028_
rlabel metal2 17696 26936 17696 26936 0 _029_
rlabel metal3 16520 27160 16520 27160 0 _030_
rlabel metal3 18200 24696 18200 24696 0 _031_
rlabel metal3 14364 25368 14364 25368 0 _032_
rlabel metal2 14336 25480 14336 25480 0 _033_
rlabel metal3 22232 14280 22232 14280 0 _034_
rlabel metal2 22120 19880 22120 19880 0 _035_
rlabel metal2 23128 18648 23128 18648 0 _036_
rlabel metal2 24024 17752 24024 17752 0 _037_
rlabel metal3 18760 26040 18760 26040 0 _038_
rlabel metal2 21784 18648 21784 18648 0 _039_
rlabel metal3 27048 25424 27048 25424 0 _040_
rlabel metal2 19320 25816 19320 25816 0 _041_
rlabel metal2 18312 27356 18312 27356 0 _042_
rlabel metal2 27608 25312 27608 25312 0 _043_
rlabel metal2 22792 20496 22792 20496 0 _044_
rlabel metal2 21336 22008 21336 22008 0 _045_
rlabel metal2 23016 21280 23016 21280 0 _046_
rlabel metal2 22008 18424 22008 18424 0 _047_
rlabel metal3 26152 17640 26152 17640 0 _048_
rlabel metal2 25368 17360 25368 17360 0 _049_
rlabel metal2 27832 22120 27832 22120 0 _050_
rlabel metal2 28168 22568 28168 22568 0 _051_
rlabel metal2 26040 20888 26040 20888 0 _052_
rlabel metal2 26152 19096 26152 19096 0 _053_
rlabel metal2 15064 26992 15064 26992 0 _054_
rlabel metal2 22904 26208 22904 26208 0 _055_
rlabel metal2 22792 25760 22792 25760 0 _056_
rlabel metal2 17640 19264 17640 19264 0 _057_
rlabel metal3 26488 15512 26488 15512 0 _058_
rlabel metal2 21224 13328 21224 13328 0 _059_
rlabel metal2 23240 14616 23240 14616 0 _060_
rlabel metal2 16016 15176 16016 15176 0 _061_
rlabel metal2 19656 13720 19656 13720 0 _062_
rlabel metal2 15960 18872 15960 18872 0 _063_
rlabel metal2 19712 14504 19712 14504 0 _064_
rlabel metal2 27720 17640 27720 17640 0 _065_
rlabel metal2 21672 18368 21672 18368 0 _066_
rlabel metal2 26936 14448 26936 14448 0 _067_
rlabel metal2 24248 16856 24248 16856 0 _068_
rlabel metal2 21560 14112 21560 14112 0 _069_
rlabel metal2 21336 14784 21336 14784 0 _070_
rlabel metal2 16520 17864 16520 17864 0 _071_
rlabel metal2 19768 20104 19768 20104 0 _072_
rlabel metal3 19768 19096 19768 19096 0 _073_
rlabel metal2 15736 22232 15736 22232 0 _074_
rlabel metal2 15288 22232 15288 22232 0 _075_
rlabel metal3 17192 23016 17192 23016 0 _076_
rlabel metal2 21448 22624 21448 22624 0 _077_
rlabel metal2 18760 15848 18760 15848 0 _078_
rlabel metal3 17808 17528 17808 17528 0 _079_
rlabel metal2 19208 18480 19208 18480 0 _080_
rlabel metal3 18872 18648 18872 18648 0 _081_
rlabel metal2 17192 21952 17192 21952 0 _082_
rlabel metal2 19320 19936 19320 19936 0 _083_
rlabel metal2 22400 19992 22400 19992 0 _084_
rlabel metal3 20832 18200 20832 18200 0 _085_
rlabel metal2 18200 15344 18200 15344 0 _086_
rlabel metal3 23072 14504 23072 14504 0 _087_
rlabel metal3 22064 14504 22064 14504 0 _088_
rlabel metal2 17640 23520 17640 23520 0 _089_
rlabel metal2 13832 26656 13832 26656 0 _090_
rlabel metal2 14280 23912 14280 23912 0 _091_
rlabel metal2 18312 22736 18312 22736 0 _092_
rlabel metal2 19320 26908 19320 26908 0 _093_
rlabel metal2 18536 19264 18536 19264 0 _094_
rlabel metal3 18928 19768 18928 19768 0 _095_
rlabel metal2 14616 21112 14616 21112 0 _096_
rlabel metal2 21336 24416 21336 24416 0 _097_
rlabel metal3 18088 26936 18088 26936 0 _098_
rlabel metal3 24192 24920 24192 24920 0 _099_
rlabel metal2 28392 23016 28392 23016 0 _100_
rlabel metal2 26376 25816 26376 25816 0 _101_
rlabel metal2 14280 18480 14280 18480 0 _102_
rlabel metal2 20440 25144 20440 25144 0 _103_
rlabel metal2 26712 18872 26712 18872 0 _104_
rlabel metal2 17864 22736 17864 22736 0 _105_
rlabel metal2 21560 22792 21560 22792 0 _106_
rlabel metal2 20720 20104 20720 20104 0 _107_
rlabel metal2 14728 20048 14728 20048 0 _108_
rlabel metal2 21336 26908 21336 26908 0 _109_
rlabel metal2 21168 27160 21168 27160 0 _110_
rlabel metal3 2478 27608 2478 27608 0 clk
rlabel metal2 22904 21112 22904 21112 0 clknet_0_clk
rlabel metal2 17528 28336 17528 28336 0 clknet_1_0__leaf_clk
rlabel metal2 22680 27440 22680 27440 0 clknet_1_1__leaf_clk
rlabel metal2 14952 17976 14952 17976 0 dut35.count\[0\]
rlabel metal2 15064 17192 15064 17192 0 dut35.count\[1\]
rlabel metal2 14168 22288 14168 22288 0 dut35.count\[2\]
rlabel metal2 16408 22008 16408 22008 0 dut35.count\[3\]
rlabel metal2 29512 17192 29512 17192 0 net1
rlabel metal2 37352 23352 37352 23352 0 net10
rlabel metal3 31920 21672 31920 21672 0 net11
rlabel metal2 29176 19488 29176 19488 0 net12
rlabel metal2 20496 12712 20496 12712 0 net13
rlabel metal2 27832 25256 27832 25256 0 net14
rlabel metal2 25368 6356 25368 6356 0 net15
rlabel metal2 16072 13048 16072 13048 0 net16
rlabel metal3 20216 38024 20216 38024 0 net17
rlabel metal3 31920 17808 31920 17808 0 net18
rlabel metal2 4312 26600 4312 26600 0 net19
rlabel metal2 27832 14672 27832 14672 0 net2
rlabel metal2 16912 26936 16912 26936 0 net20
rlabel metal3 23800 27720 23800 27720 0 net21
rlabel metal2 27608 26992 27608 26992 0 net22
rlabel metal2 11032 23464 11032 23464 0 net23
rlabel metal2 37912 22624 37912 22624 0 net24
rlabel metal3 18648 3528 18648 3528 0 net25
rlabel metal2 22344 37464 22344 37464 0 net26
rlabel metal2 23576 5964 23576 5964 0 net3
rlabel metal2 25592 32200 25592 32200 0 net4
rlabel metal2 28168 18256 28168 18256 0 net5
rlabel metal2 24584 5964 24584 5964 0 net6
rlabel metal2 14336 38024 14336 38024 0 net7
rlabel metal2 29960 21728 29960 21728 0 net8
rlabel metal2 13944 27328 13944 27328 0 net9
rlabel metal2 40040 17640 40040 17640 0 segm[10]
rlabel metal2 40040 15008 40040 15008 0 segm[11]
rlabel metal2 22232 2086 22232 2086 0 segm[12]
rlabel metal2 24920 39354 24920 39354 0 segm[13]
rlabel metal2 40040 19096 40040 19096 0 segm[1]
rlabel metal2 23576 854 23576 854 0 segm[2]
rlabel metal2 14840 39746 14840 39746 0 segm[3]
rlabel metal2 40040 22344 40040 22344 0 segm[4]
rlabel metal2 14168 39354 14168 39354 0 segm[5]
rlabel metal2 40040 23800 40040 23800 0 segm[6]
rlabel metal2 40040 21504 40040 21504 0 segm[7]
rlabel metal2 40040 19656 40040 19656 0 segm[8]
rlabel metal2 20216 2422 20216 2422 0 segm[9]
rlabel metal2 40040 25816 40040 25816 0 sel[0]
rlabel metal2 24920 2422 24920 2422 0 sel[10]
rlabel metal2 16184 2478 16184 2478 0 sel[11]
rlabel metal2 19544 39690 19544 39690 0 sel[1]
rlabel metal3 40642 18200 40642 18200 0 sel[2]
rlabel metal3 1358 26264 1358 26264 0 sel[3]
rlabel metal2 17528 39746 17528 39746 0 sel[4]
rlabel metal2 22904 39746 22904 39746 0 sel[5]
rlabel metal2 40040 26712 40040 26712 0 sel[6]
rlabel metal3 1358 23576 1358 23576 0 sel[7]
rlabel metal3 40642 22904 40642 22904 0 sel[8]
rlabel metal2 19544 2086 19544 2086 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 42000 42000
<< end >>
