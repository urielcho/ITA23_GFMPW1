VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO ita6
  CLASS BLOCK ;
  FOREIGN ita6 ;
  ORIGIN 0.000 0.000 ;
  SIZE 210.000 BY 210.000 ;
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 4.738000 ;
    ANTENNADIFFAREA 0.410400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 137.760 4.000 138.320 ;
    END
  END clk
  PIN segm[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal3 ;
        RECT 206.000 131.040 210.000 131.600 ;
    END
  END segm[0]
  PIN segm[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 94.080 4.000 94.640 ;
    END
  END segm[10]
  PIN segm[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 110.880 206.000 111.440 210.000 ;
    END
  END segm[11]
  PIN segm[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 120.960 206.000 121.520 210.000 ;
    END
  END segm[12]
  PIN segm[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 114.240 0.000 114.800 4.000 ;
    END
  END segm[13]
  PIN segm[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 206.000 120.960 210.000 121.520 ;
    END
  END segm[1]
  PIN segm[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 206.000 110.880 210.000 111.440 ;
    END
  END segm[2]
  PIN segm[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.360800 ;
    PORT
      LAYER Metal2 ;
        RECT 100.800 0.000 101.360 4.000 ;
    END
  END segm[3]
  PIN segm[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 206.000 117.600 210.000 118.160 ;
    END
  END segm[4]
  PIN segm[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 206.000 104.160 210.000 104.720 ;
    END
  END segm[5]
  PIN segm[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 131.040 4.000 131.600 ;
    END
  END segm[6]
  PIN segm[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 114.240 4.000 114.800 ;
    END
  END segm[7]
  PIN segm[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 206.000 127.680 210.000 128.240 ;
    END
  END segm[8]
  PIN segm[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 206.000 124.320 210.000 124.880 ;
    END
  END segm[9]
  PIN sel[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 206.000 87.360 210.000 87.920 ;
    END
  END sel[0]
  PIN sel[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 94.080 0.000 94.640 4.000 ;
    END
  END sel[10]
  PIN sel[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 97.440 206.000 98.000 210.000 ;
    END
  END sel[11]
  PIN sel[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 206.000 107.520 210.000 108.080 ;
    END
  END sel[1]
  PIN sel[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 127.680 4.000 128.240 ;
    END
  END sel[2]
  PIN sel[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 206.000 100.800 210.000 101.360 ;
    END
  END sel[3]
  PIN sel[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 206.000 94.080 210.000 94.640 ;
    END
  END sel[4]
  PIN sel[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 117.600 4.000 118.160 ;
    END
  END sel[5]
  PIN sel[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 90.720 206.000 91.280 210.000 ;
    END
  END sel[6]
  PIN sel[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal3 ;
        RECT 206.000 114.240 210.000 114.800 ;
    END
  END sel[7]
  PIN sel[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 124.320 0.000 124.880 4.000 ;
    END
  END sel[8]
  PIN sel[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    ANTENNADIFFAREA 4.731200 ;
    PORT
      LAYER Metal2 ;
        RECT 104.160 0.000 104.720 4.000 ;
    END
  END sel[9]
  PIN vdd
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal4 ;
        RECT 22.240 15.380 23.840 192.380 ;
    END
    PORT
      LAYER Metal4 ;
        RECT 175.840 15.380 177.440 192.380 ;
    END
  END vdd
  PIN vss
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal4 ;
        RECT 99.040 15.380 100.640 192.380 ;
    END
  END vss
  OBS
      LAYER Metal1 ;
        RECT 6.720 15.380 203.280 192.380 ;
      LAYER Metal2 ;
        RECT 9.660 205.700 90.420 206.000 ;
        RECT 91.580 205.700 97.140 206.000 ;
        RECT 98.300 205.700 110.580 206.000 ;
        RECT 111.740 205.700 120.660 206.000 ;
        RECT 121.820 205.700 201.460 206.000 ;
        RECT 9.660 4.300 201.460 205.700 ;
        RECT 9.660 4.000 93.780 4.300 ;
        RECT 94.940 4.000 100.500 4.300 ;
        RECT 101.660 4.000 103.860 4.300 ;
        RECT 105.020 4.000 113.940 4.300 ;
        RECT 115.100 4.000 124.020 4.300 ;
        RECT 125.180 4.000 201.460 4.300 ;
      LAYER Metal3 ;
        RECT 4.000 138.620 206.000 192.220 ;
        RECT 4.300 137.460 206.000 138.620 ;
        RECT 4.000 131.900 206.000 137.460 ;
        RECT 4.300 130.740 205.700 131.900 ;
        RECT 4.000 128.540 206.000 130.740 ;
        RECT 4.300 127.380 205.700 128.540 ;
        RECT 4.000 125.180 206.000 127.380 ;
        RECT 4.000 124.020 205.700 125.180 ;
        RECT 4.000 121.820 206.000 124.020 ;
        RECT 4.000 120.660 205.700 121.820 ;
        RECT 4.000 118.460 206.000 120.660 ;
        RECT 4.300 117.300 205.700 118.460 ;
        RECT 4.000 115.100 206.000 117.300 ;
        RECT 4.300 113.940 205.700 115.100 ;
        RECT 4.000 111.740 206.000 113.940 ;
        RECT 4.000 110.580 205.700 111.740 ;
        RECT 4.000 108.380 206.000 110.580 ;
        RECT 4.000 107.220 205.700 108.380 ;
        RECT 4.000 105.020 206.000 107.220 ;
        RECT 4.000 103.860 205.700 105.020 ;
        RECT 4.000 101.660 206.000 103.860 ;
        RECT 4.000 100.500 205.700 101.660 ;
        RECT 4.000 94.940 206.000 100.500 ;
        RECT 4.300 93.780 205.700 94.940 ;
        RECT 4.000 88.220 206.000 93.780 ;
        RECT 4.000 87.060 205.700 88.220 ;
        RECT 4.000 15.540 206.000 87.060 ;
      LAYER Metal4 ;
        RECT 108.780 93.050 109.060 111.910 ;
  END
END ita6
END LIBRARY

