magic
tech gf180mcuD
magscale 1 5
timestamp 1699642890
<< metal1 >>
rect 672 19221 20328 19238
rect 672 19195 2239 19221
rect 2265 19195 2291 19221
rect 2317 19195 2343 19221
rect 2369 19195 17599 19221
rect 17625 19195 17651 19221
rect 17677 19195 17703 19221
rect 17729 19195 20328 19221
rect 672 19178 20328 19195
rect 9311 19137 9337 19143
rect 9311 19105 9337 19111
rect 11215 19137 11241 19143
rect 11215 19105 11241 19111
rect 13063 19137 13089 19143
rect 13063 19105 13089 19111
rect 8969 18999 8975 19025
rect 9001 18999 9007 19025
rect 10705 18999 10711 19025
rect 10737 18999 10743 19025
rect 12665 18999 12671 19025
rect 12697 18999 12703 19025
rect 672 18829 20328 18846
rect 672 18803 9919 18829
rect 9945 18803 9971 18829
rect 9997 18803 10023 18829
rect 10049 18803 20328 18829
rect 672 18786 20328 18803
rect 9367 18745 9393 18751
rect 9367 18713 9393 18719
rect 11383 18745 11409 18751
rect 11383 18713 11409 18719
rect 9025 18607 9031 18633
rect 9057 18607 9063 18633
rect 10985 18607 10991 18633
rect 11017 18607 11023 18633
rect 672 18437 20328 18454
rect 672 18411 2239 18437
rect 2265 18411 2291 18437
rect 2317 18411 2343 18437
rect 2369 18411 17599 18437
rect 17625 18411 17651 18437
rect 17677 18411 17703 18437
rect 17729 18411 20328 18437
rect 672 18394 20328 18411
rect 8639 18353 8665 18359
rect 8639 18321 8665 18327
rect 9585 18215 9591 18241
rect 9617 18215 9623 18241
rect 672 18045 20328 18062
rect 672 18019 9919 18045
rect 9945 18019 9971 18045
rect 9997 18019 10023 18045
rect 10049 18019 20328 18045
rect 672 18002 20328 18019
rect 672 17653 20328 17670
rect 672 17627 2239 17653
rect 2265 17627 2291 17653
rect 2317 17627 2343 17653
rect 2369 17627 17599 17653
rect 17625 17627 17651 17653
rect 17677 17627 17703 17653
rect 17729 17627 20328 17653
rect 672 17610 20328 17627
rect 672 17261 20328 17278
rect 672 17235 9919 17261
rect 9945 17235 9971 17261
rect 9997 17235 10023 17261
rect 10049 17235 20328 17261
rect 672 17218 20328 17235
rect 672 16869 20328 16886
rect 672 16843 2239 16869
rect 2265 16843 2291 16869
rect 2317 16843 2343 16869
rect 2369 16843 17599 16869
rect 17625 16843 17651 16869
rect 17677 16843 17703 16869
rect 17729 16843 20328 16869
rect 672 16826 20328 16843
rect 672 16477 20328 16494
rect 672 16451 9919 16477
rect 9945 16451 9971 16477
rect 9997 16451 10023 16477
rect 10049 16451 20328 16477
rect 672 16434 20328 16451
rect 672 16085 20328 16102
rect 672 16059 2239 16085
rect 2265 16059 2291 16085
rect 2317 16059 2343 16085
rect 2369 16059 17599 16085
rect 17625 16059 17651 16085
rect 17677 16059 17703 16085
rect 17729 16059 20328 16085
rect 672 16042 20328 16059
rect 672 15693 20328 15710
rect 672 15667 9919 15693
rect 9945 15667 9971 15693
rect 9997 15667 10023 15693
rect 10049 15667 20328 15693
rect 672 15650 20328 15667
rect 672 15301 20328 15318
rect 672 15275 2239 15301
rect 2265 15275 2291 15301
rect 2317 15275 2343 15301
rect 2369 15275 17599 15301
rect 17625 15275 17651 15301
rect 17677 15275 17703 15301
rect 17729 15275 20328 15301
rect 672 15258 20328 15275
rect 672 14909 20328 14926
rect 672 14883 9919 14909
rect 9945 14883 9971 14909
rect 9997 14883 10023 14909
rect 10049 14883 20328 14909
rect 672 14866 20328 14883
rect 9585 14687 9591 14713
rect 9617 14687 9623 14713
rect 11327 14657 11353 14663
rect 9977 14631 9983 14657
rect 10009 14631 10015 14657
rect 11041 14631 11047 14657
rect 11073 14631 11079 14657
rect 11327 14625 11353 14631
rect 672 14517 20328 14534
rect 672 14491 2239 14517
rect 2265 14491 2291 14517
rect 2317 14491 2343 14517
rect 2369 14491 17599 14517
rect 17625 14491 17651 14517
rect 17677 14491 17703 14517
rect 17729 14491 20328 14517
rect 672 14474 20328 14491
rect 8527 14321 8553 14327
rect 8527 14289 8553 14295
rect 672 14125 20328 14142
rect 672 14099 9919 14125
rect 9945 14099 9971 14125
rect 9997 14099 10023 14125
rect 10049 14099 20328 14125
rect 672 14082 20328 14099
rect 9031 14041 9057 14047
rect 8857 14015 8863 14041
rect 8889 14015 8895 14041
rect 9031 14009 9057 14015
rect 11215 14041 11241 14047
rect 11215 14009 11241 14015
rect 7009 13903 7015 13929
rect 7041 13903 7047 13929
rect 9585 13903 9591 13929
rect 9617 13903 9623 13929
rect 7345 13847 7351 13873
rect 7377 13847 7383 13873
rect 8409 13847 8415 13873
rect 8441 13847 8447 13873
rect 9921 13847 9927 13873
rect 9953 13847 9959 13873
rect 10985 13847 10991 13873
rect 11017 13847 11023 13873
rect 672 13733 20328 13750
rect 672 13707 2239 13733
rect 2265 13707 2291 13733
rect 2317 13707 2343 13733
rect 2369 13707 17599 13733
rect 17625 13707 17651 13733
rect 17677 13707 17703 13733
rect 17729 13707 20328 13733
rect 672 13690 20328 13707
rect 10711 13649 10737 13655
rect 10711 13617 10737 13623
rect 967 13593 993 13599
rect 9591 13593 9617 13599
rect 9081 13567 9087 13593
rect 9113 13567 9119 13593
rect 967 13561 993 13567
rect 9591 13561 9617 13567
rect 20007 13593 20033 13599
rect 20007 13561 20033 13567
rect 10151 13537 10177 13543
rect 2137 13511 2143 13537
rect 2169 13511 2175 13537
rect 7681 13511 7687 13537
rect 7713 13511 7719 13537
rect 10151 13505 10177 13511
rect 10319 13537 10345 13543
rect 18937 13511 18943 13537
rect 18969 13511 18975 13537
rect 10319 13505 10345 13511
rect 9199 13481 9225 13487
rect 8017 13455 8023 13481
rect 8049 13455 8055 13481
rect 9199 13449 9225 13455
rect 9311 13481 9337 13487
rect 9311 13449 9337 13455
rect 9367 13481 9393 13487
rect 9367 13449 9393 13455
rect 10655 13481 10681 13487
rect 10655 13449 10681 13455
rect 10711 13481 10737 13487
rect 10711 13449 10737 13455
rect 10263 13425 10289 13431
rect 10263 13393 10289 13399
rect 672 13341 20328 13358
rect 672 13315 9919 13341
rect 9945 13315 9971 13341
rect 9997 13315 10023 13341
rect 10049 13315 20328 13341
rect 672 13298 20328 13315
rect 7967 13257 7993 13263
rect 7967 13225 7993 13231
rect 8247 13257 8273 13263
rect 8247 13225 8273 13231
rect 8751 13257 8777 13263
rect 8751 13225 8777 13231
rect 10655 13257 10681 13263
rect 10655 13225 10681 13231
rect 8079 13201 8105 13207
rect 8079 13169 8105 13175
rect 8135 13201 8161 13207
rect 8135 13169 8161 13175
rect 8359 13201 8385 13207
rect 8359 13169 8385 13175
rect 9927 13201 9953 13207
rect 9927 13169 9953 13175
rect 10543 13201 10569 13207
rect 10543 13169 10569 13175
rect 12671 13201 12697 13207
rect 12671 13169 12697 13175
rect 13567 13201 13593 13207
rect 13567 13169 13593 13175
rect 8415 13145 8441 13151
rect 7681 13119 7687 13145
rect 7713 13119 7719 13145
rect 8415 13113 8441 13119
rect 8639 13145 8665 13151
rect 8639 13113 8665 13119
rect 8807 13145 8833 13151
rect 8807 13113 8833 13119
rect 9871 13145 9897 13151
rect 9871 13113 9897 13119
rect 10711 13145 10737 13151
rect 12727 13145 12753 13151
rect 10929 13119 10935 13145
rect 10961 13119 10967 13145
rect 10711 13113 10737 13119
rect 12727 13113 12753 13119
rect 13511 13145 13537 13151
rect 18825 13119 18831 13145
rect 18857 13119 18863 13145
rect 13511 13113 13537 13119
rect 12951 13089 12977 13095
rect 6281 13063 6287 13089
rect 6313 13063 6319 13089
rect 7345 13063 7351 13089
rect 7377 13063 7383 13089
rect 11265 13063 11271 13089
rect 11297 13063 11303 13089
rect 12329 13063 12335 13089
rect 12361 13063 12367 13089
rect 12951 13057 12977 13063
rect 14519 13089 14545 13095
rect 14519 13057 14545 13063
rect 9927 13033 9953 13039
rect 9927 13001 9953 13007
rect 12671 13033 12697 13039
rect 12671 13001 12697 13007
rect 13567 13033 13593 13039
rect 13567 13001 13593 13007
rect 14463 13033 14489 13039
rect 14463 13001 14489 13007
rect 20007 13033 20033 13039
rect 20007 13001 20033 13007
rect 672 12949 20328 12966
rect 672 12923 2239 12949
rect 2265 12923 2291 12949
rect 2317 12923 2343 12949
rect 2369 12923 17599 12949
rect 17625 12923 17651 12949
rect 17677 12923 17703 12949
rect 17729 12923 20328 12949
rect 672 12906 20328 12923
rect 7687 12809 7713 12815
rect 7687 12777 7713 12783
rect 7855 12809 7881 12815
rect 7855 12777 7881 12783
rect 8247 12809 8273 12815
rect 8247 12777 8273 12783
rect 11775 12809 11801 12815
rect 14065 12783 14071 12809
rect 14097 12783 14103 12809
rect 11775 12777 11801 12783
rect 7911 12753 7937 12759
rect 7911 12721 7937 12727
rect 8191 12753 8217 12759
rect 8191 12721 8217 12727
rect 8359 12753 8385 12759
rect 8359 12721 8385 12727
rect 12055 12753 12081 12759
rect 12055 12721 12081 12727
rect 12447 12753 12473 12759
rect 12665 12727 12671 12753
rect 12697 12727 12703 12753
rect 12447 12721 12473 12727
rect 10201 12671 10207 12697
rect 10233 12671 10239 12697
rect 13001 12671 13007 12697
rect 13033 12671 13039 12697
rect 8135 12641 8161 12647
rect 8135 12609 8161 12615
rect 8303 12641 8329 12647
rect 8303 12609 8329 12615
rect 10375 12641 10401 12647
rect 10375 12609 10401 12615
rect 10767 12641 10793 12647
rect 11719 12641 11745 12647
rect 10929 12615 10935 12641
rect 10961 12615 10967 12641
rect 10767 12609 10793 12615
rect 11719 12609 11745 12615
rect 11831 12641 11857 12647
rect 11831 12609 11857 12615
rect 672 12557 20328 12574
rect 672 12531 9919 12557
rect 9945 12531 9971 12557
rect 9997 12531 10023 12557
rect 10049 12531 20328 12557
rect 672 12514 20328 12531
rect 12895 12473 12921 12479
rect 8353 12447 8359 12473
rect 8385 12447 8391 12473
rect 12895 12441 12921 12447
rect 13343 12473 13369 12479
rect 13343 12441 13369 12447
rect 8191 12361 8217 12367
rect 12839 12361 12865 12367
rect 9809 12335 9815 12361
rect 9841 12335 9847 12361
rect 8191 12329 8217 12335
rect 12839 12329 12865 12335
rect 12951 12361 12977 12367
rect 12951 12329 12977 12335
rect 13175 12361 13201 12367
rect 13505 12335 13511 12361
rect 13537 12335 13543 12361
rect 13175 12329 13201 12335
rect 8079 12305 8105 12311
rect 8079 12273 8105 12279
rect 8807 12305 8833 12311
rect 10481 12279 10487 12305
rect 10513 12279 10519 12305
rect 13897 12279 13903 12305
rect 13929 12279 13935 12305
rect 14961 12279 14967 12305
rect 14993 12279 14999 12305
rect 8807 12273 8833 12279
rect 672 12165 20328 12182
rect 672 12139 2239 12165
rect 2265 12139 2291 12165
rect 2317 12139 2343 12165
rect 2369 12139 17599 12165
rect 17625 12139 17651 12165
rect 17677 12139 17703 12165
rect 17729 12139 20328 12165
rect 672 12122 20328 12139
rect 8863 12081 8889 12087
rect 8863 12049 8889 12055
rect 967 12025 993 12031
rect 10823 12025 10849 12031
rect 6729 11999 6735 12025
rect 6761 11999 6767 12025
rect 9137 11999 9143 12025
rect 9169 11999 9175 12025
rect 967 11993 993 11999
rect 10823 11993 10849 11999
rect 8751 11969 8777 11975
rect 2137 11943 2143 11969
rect 2169 11943 2175 11969
rect 8185 11943 8191 11969
rect 8217 11943 8223 11969
rect 8577 11943 8583 11969
rect 8609 11943 8615 11969
rect 8751 11937 8777 11943
rect 9367 11969 9393 11975
rect 9367 11937 9393 11943
rect 10151 11969 10177 11975
rect 10151 11937 10177 11943
rect 13343 11969 13369 11975
rect 13343 11937 13369 11943
rect 13623 11969 13649 11975
rect 13623 11937 13649 11943
rect 13735 11969 13761 11975
rect 13897 11943 13903 11969
rect 13929 11943 13935 11969
rect 14177 11943 14183 11969
rect 14209 11943 14215 11969
rect 13735 11937 13761 11943
rect 8471 11913 8497 11919
rect 7793 11887 7799 11913
rect 7825 11887 7831 11913
rect 8471 11881 8497 11887
rect 9983 11913 10009 11919
rect 9983 11881 10009 11887
rect 13399 11913 13425 11919
rect 13399 11881 13425 11887
rect 8415 11857 8441 11863
rect 8415 11825 8441 11831
rect 8527 11857 8553 11863
rect 8527 11825 8553 11831
rect 9087 11857 9113 11863
rect 9087 11825 9113 11831
rect 9199 11857 9225 11863
rect 9199 11825 9225 11831
rect 10039 11857 10065 11863
rect 10039 11825 10065 11831
rect 13511 11857 13537 11863
rect 13511 11825 13537 11831
rect 14071 11857 14097 11863
rect 14071 11825 14097 11831
rect 672 11773 20328 11790
rect 672 11747 9919 11773
rect 9945 11747 9971 11773
rect 9997 11747 10023 11773
rect 10049 11747 20328 11773
rect 672 11730 20328 11747
rect 8079 11689 8105 11695
rect 8079 11657 8105 11663
rect 12671 11689 12697 11695
rect 12671 11657 12697 11663
rect 8975 11633 9001 11639
rect 5889 11607 5895 11633
rect 5921 11607 5927 11633
rect 8975 11601 9001 11607
rect 9031 11633 9057 11639
rect 9031 11601 9057 11607
rect 7183 11577 7209 11583
rect 5553 11551 5559 11577
rect 5585 11551 5591 11577
rect 7183 11545 7209 11551
rect 8023 11577 8049 11583
rect 8023 11545 8049 11551
rect 8359 11577 8385 11583
rect 9249 11551 9255 11577
rect 9281 11551 9287 11577
rect 10929 11551 10935 11577
rect 10961 11551 10967 11577
rect 13617 11551 13623 11577
rect 13649 11551 13655 11577
rect 8359 11545 8385 11551
rect 13735 11521 13761 11527
rect 6953 11495 6959 11521
rect 6985 11495 6991 11521
rect 9641 11495 9647 11521
rect 9673 11495 9679 11521
rect 10705 11495 10711 11521
rect 10737 11495 10743 11521
rect 11265 11495 11271 11521
rect 11297 11495 11303 11521
rect 12329 11495 12335 11521
rect 12361 11495 12367 11521
rect 13735 11489 13761 11495
rect 8079 11465 8105 11471
rect 8079 11433 8105 11439
rect 8975 11465 9001 11471
rect 8975 11433 9001 11439
rect 13791 11465 13817 11471
rect 13791 11433 13817 11439
rect 672 11381 20328 11398
rect 672 11355 2239 11381
rect 2265 11355 2291 11381
rect 2317 11355 2343 11381
rect 2369 11355 17599 11381
rect 17625 11355 17651 11381
rect 17677 11355 17703 11381
rect 17729 11355 20328 11381
rect 672 11338 20328 11355
rect 9479 11297 9505 11303
rect 9479 11265 9505 11271
rect 10879 11241 10905 11247
rect 10879 11209 10905 11215
rect 11495 11241 11521 11247
rect 13959 11241 13985 11247
rect 12889 11215 12895 11241
rect 12921 11215 12927 11241
rect 11495 11209 11521 11215
rect 13959 11209 13985 11215
rect 20007 11241 20033 11247
rect 20007 11209 20033 11215
rect 8471 11185 8497 11191
rect 7737 11159 7743 11185
rect 7769 11159 7775 11185
rect 8241 11159 8247 11185
rect 8273 11159 8279 11185
rect 8471 11153 8497 11159
rect 8807 11185 8833 11191
rect 8807 11153 8833 11159
rect 8919 11185 8945 11191
rect 8919 11153 8945 11159
rect 9423 11185 9449 11191
rect 9423 11153 9449 11159
rect 10599 11185 10625 11191
rect 10599 11153 10625 11159
rect 10935 11185 10961 11191
rect 10935 11153 10961 11159
rect 11103 11185 11129 11191
rect 11103 11153 11129 11159
rect 11439 11185 11465 11191
rect 11439 11153 11465 11159
rect 11607 11185 11633 11191
rect 11607 11153 11633 11159
rect 12055 11185 12081 11191
rect 12055 11153 12081 11159
rect 12727 11185 12753 11191
rect 14065 11159 14071 11185
rect 14097 11159 14103 11185
rect 18825 11159 18831 11185
rect 18857 11159 18863 11185
rect 12727 11153 12753 11159
rect 10151 11129 10177 11135
rect 7849 11103 7855 11129
rect 7881 11103 7887 11129
rect 9921 11103 9927 11129
rect 9953 11103 9959 11129
rect 10151 11097 10177 11103
rect 10319 11129 10345 11135
rect 10319 11097 10345 11103
rect 11215 11129 11241 11135
rect 11215 11097 11241 11103
rect 11719 11129 11745 11135
rect 12895 11129 12921 11135
rect 13903 11129 13929 11135
rect 11881 11103 11887 11129
rect 11913 11103 11919 11129
rect 12945 11103 12951 11129
rect 12977 11103 12983 11129
rect 11719 11097 11745 11103
rect 12895 11097 12921 11103
rect 13903 11097 13929 11103
rect 9479 11073 9505 11079
rect 9081 11047 9087 11073
rect 9113 11047 9119 11073
rect 9479 11041 9505 11047
rect 9759 11073 9785 11079
rect 9759 11041 9785 11047
rect 10095 11073 10121 11079
rect 10095 11041 10121 11047
rect 10207 11073 10233 11079
rect 10207 11041 10233 11047
rect 10823 11073 10849 11079
rect 10823 11041 10849 11047
rect 11159 11073 11185 11079
rect 11159 11041 11185 11047
rect 12839 11073 12865 11079
rect 12839 11041 12865 11047
rect 672 10989 20328 11006
rect 672 10963 9919 10989
rect 9945 10963 9971 10989
rect 9997 10963 10023 10989
rect 10049 10963 20328 10989
rect 672 10946 20328 10963
rect 12783 10905 12809 10911
rect 12783 10873 12809 10879
rect 13175 10905 13201 10911
rect 13175 10873 13201 10879
rect 8695 10849 8721 10855
rect 8409 10823 8415 10849
rect 8441 10823 8447 10849
rect 8695 10817 8721 10823
rect 12671 10849 12697 10855
rect 13729 10823 13735 10849
rect 13761 10823 13767 10849
rect 12671 10817 12697 10823
rect 7855 10793 7881 10799
rect 8807 10793 8833 10799
rect 5833 10767 5839 10793
rect 5865 10767 5871 10793
rect 7681 10767 7687 10793
rect 7713 10767 7719 10793
rect 8297 10767 8303 10793
rect 8329 10767 8335 10793
rect 7855 10761 7881 10767
rect 8807 10761 8833 10767
rect 9479 10793 9505 10799
rect 12615 10793 12641 10799
rect 9697 10767 9703 10793
rect 9729 10767 9735 10793
rect 13337 10767 13343 10793
rect 13369 10767 13375 10793
rect 9479 10761 9505 10767
rect 12615 10761 12641 10767
rect 7407 10737 7433 10743
rect 6169 10711 6175 10737
rect 6201 10711 6207 10737
rect 7233 10711 7239 10737
rect 7265 10711 7271 10737
rect 10929 10711 10935 10737
rect 10961 10711 10967 10737
rect 14793 10711 14799 10737
rect 14825 10711 14831 10737
rect 7407 10705 7433 10711
rect 8975 10681 9001 10687
rect 8975 10649 9001 10655
rect 672 10597 20328 10614
rect 672 10571 2239 10597
rect 2265 10571 2291 10597
rect 2317 10571 2343 10597
rect 2369 10571 17599 10597
rect 17625 10571 17651 10597
rect 17677 10571 17703 10597
rect 17729 10571 20328 10597
rect 672 10554 20328 10571
rect 7407 10457 7433 10463
rect 11383 10457 11409 10463
rect 20007 10457 20033 10463
rect 8857 10431 8863 10457
rect 8889 10431 8895 10457
rect 12889 10431 12895 10457
rect 12921 10431 12927 10457
rect 7407 10425 7433 10431
rect 11383 10425 11409 10431
rect 20007 10425 20033 10431
rect 7015 10401 7041 10407
rect 7015 10369 7041 10375
rect 9143 10401 9169 10407
rect 9927 10401 9953 10407
rect 9305 10375 9311 10401
rect 9337 10375 9343 10401
rect 9143 10369 9169 10375
rect 9927 10369 9953 10375
rect 11103 10401 11129 10407
rect 12727 10401 12753 10407
rect 11881 10375 11887 10401
rect 11913 10375 11919 10401
rect 12945 10375 12951 10401
rect 12977 10375 12983 10401
rect 13113 10375 13119 10401
rect 13145 10375 13151 10401
rect 18937 10375 18943 10401
rect 18969 10375 18975 10401
rect 11103 10369 11129 10375
rect 12727 10369 12753 10375
rect 6847 10345 6873 10351
rect 6847 10313 6873 10319
rect 8863 10345 8889 10351
rect 12839 10345 12865 10351
rect 9417 10319 9423 10345
rect 9449 10319 9455 10345
rect 8863 10313 8889 10319
rect 12839 10313 12865 10319
rect 8975 10289 9001 10295
rect 10089 10263 10095 10289
rect 10121 10263 10127 10289
rect 11769 10263 11775 10289
rect 11801 10263 11807 10289
rect 8975 10257 9001 10263
rect 672 10205 20328 10222
rect 672 10179 9919 10205
rect 9945 10179 9971 10205
rect 9997 10179 10023 10205
rect 10049 10179 20328 10205
rect 672 10162 20328 10179
rect 8415 10121 8441 10127
rect 8415 10089 8441 10095
rect 7631 10065 7657 10071
rect 11383 10065 11409 10071
rect 8241 10039 8247 10065
rect 8273 10039 8279 10065
rect 9809 10039 9815 10065
rect 9841 10039 9847 10065
rect 10257 10039 10263 10065
rect 10289 10039 10295 10065
rect 11657 10039 11663 10065
rect 11689 10039 11695 10065
rect 11937 10039 11943 10065
rect 11969 10039 11975 10065
rect 13281 10039 13287 10065
rect 13313 10039 13319 10065
rect 14681 10039 14687 10065
rect 14713 10039 14719 10065
rect 7631 10033 7657 10039
rect 11383 10033 11409 10039
rect 7071 10009 7097 10015
rect 2137 9983 2143 10009
rect 2169 9983 2175 10009
rect 7071 9977 7097 9983
rect 7183 10009 7209 10015
rect 7183 9977 7209 9983
rect 7295 10009 7321 10015
rect 7295 9977 7321 9983
rect 7407 10009 7433 10015
rect 7407 9977 7433 9983
rect 7519 10009 7545 10015
rect 7519 9977 7545 9983
rect 7687 10009 7713 10015
rect 11047 10009 11073 10015
rect 8913 9983 8919 10009
rect 8945 9983 8951 10009
rect 9473 9983 9479 10009
rect 9505 9983 9511 10009
rect 11265 9983 11271 10009
rect 11297 9983 11303 10009
rect 11601 9983 11607 10009
rect 11633 9983 11639 10009
rect 12945 9983 12951 10009
rect 12977 9983 12983 10009
rect 14569 9983 14575 10009
rect 14601 9983 14607 10009
rect 18825 9983 18831 10009
rect 18857 9983 18863 10009
rect 7687 9977 7713 9983
rect 11047 9977 11073 9983
rect 7015 9953 7041 9959
rect 7015 9921 7041 9927
rect 7911 9953 7937 9959
rect 12783 9953 12809 9959
rect 9025 9927 9031 9953
rect 9057 9927 9063 9953
rect 10873 9927 10879 9953
rect 10905 9927 10911 9953
rect 14345 9927 14351 9953
rect 14377 9927 14383 9953
rect 7911 9921 7937 9927
rect 12783 9921 12809 9927
rect 967 9897 993 9903
rect 967 9865 993 9871
rect 11439 9897 11465 9903
rect 11439 9865 11465 9871
rect 20007 9897 20033 9903
rect 20007 9865 20033 9871
rect 672 9813 20328 9830
rect 672 9787 2239 9813
rect 2265 9787 2291 9813
rect 2317 9787 2343 9813
rect 2369 9787 17599 9813
rect 17625 9787 17651 9813
rect 17677 9787 17703 9813
rect 17729 9787 20328 9813
rect 672 9770 20328 9787
rect 7295 9729 7321 9735
rect 7295 9697 7321 9703
rect 9759 9729 9785 9735
rect 9759 9697 9785 9703
rect 10655 9729 10681 9735
rect 10655 9697 10681 9703
rect 8695 9673 8721 9679
rect 12055 9673 12081 9679
rect 4993 9647 4999 9673
rect 5025 9647 5031 9673
rect 6057 9647 6063 9673
rect 6089 9647 6095 9673
rect 10761 9647 10767 9673
rect 10793 9647 10799 9673
rect 8695 9641 8721 9647
rect 12055 9641 12081 9647
rect 13455 9673 13481 9679
rect 13455 9641 13481 9647
rect 20007 9673 20033 9679
rect 20007 9641 20033 9647
rect 7071 9617 7097 9623
rect 6449 9591 6455 9617
rect 6481 9591 6487 9617
rect 7071 9585 7097 9591
rect 8023 9617 8049 9623
rect 8023 9585 8049 9591
rect 8303 9617 8329 9623
rect 8303 9585 8329 9591
rect 8583 9617 8609 9623
rect 8583 9585 8609 9591
rect 9031 9617 9057 9623
rect 11607 9617 11633 9623
rect 10817 9591 10823 9617
rect 10849 9591 10855 9617
rect 9031 9585 9057 9591
rect 11607 9585 11633 9591
rect 11831 9617 11857 9623
rect 11831 9585 11857 9591
rect 13231 9617 13257 9623
rect 13231 9585 13257 9591
rect 13399 9617 13425 9623
rect 13399 9585 13425 9591
rect 13511 9617 13537 9623
rect 13511 9585 13537 9591
rect 13791 9617 13817 9623
rect 13791 9585 13817 9591
rect 14071 9617 14097 9623
rect 18825 9591 18831 9617
rect 18857 9591 18863 9617
rect 14071 9585 14097 9591
rect 7015 9561 7041 9567
rect 7015 9529 7041 9535
rect 7295 9561 7321 9567
rect 7295 9529 7321 9535
rect 7351 9561 7377 9567
rect 8863 9561 8889 9567
rect 14015 9561 14041 9567
rect 7849 9535 7855 9561
rect 7881 9535 7887 9561
rect 9305 9535 9311 9561
rect 9337 9535 9343 9561
rect 9473 9535 9479 9561
rect 9505 9535 9511 9561
rect 7351 9529 7377 9535
rect 8863 9529 8889 9535
rect 14015 9529 14041 9535
rect 14575 9561 14601 9567
rect 14575 9529 14601 9535
rect 14743 9561 14769 9567
rect 14743 9529 14769 9535
rect 6791 9505 6817 9511
rect 6791 9473 6817 9479
rect 6903 9505 6929 9511
rect 6903 9473 6929 9479
rect 8135 9505 8161 9511
rect 8135 9473 8161 9479
rect 8247 9505 8273 9511
rect 8247 9473 8273 9479
rect 8751 9505 8777 9511
rect 9815 9505 9841 9511
rect 9081 9479 9087 9505
rect 9113 9479 9119 9505
rect 8751 9473 8777 9479
rect 9815 9473 9841 9479
rect 9871 9505 9897 9511
rect 11159 9505 11185 9511
rect 11775 9505 11801 9511
rect 10985 9479 10991 9505
rect 11017 9479 11023 9505
rect 11433 9479 11439 9505
rect 11465 9479 11471 9505
rect 9871 9473 9897 9479
rect 11159 9473 11185 9479
rect 11775 9473 11801 9479
rect 11999 9505 12025 9511
rect 11999 9473 12025 9479
rect 13623 9505 13649 9511
rect 13623 9473 13649 9479
rect 13903 9505 13929 9511
rect 13903 9473 13929 9479
rect 14631 9505 14657 9511
rect 14631 9473 14657 9479
rect 672 9421 20328 9438
rect 672 9395 9919 9421
rect 9945 9395 9971 9421
rect 9997 9395 10023 9421
rect 10049 9395 20328 9421
rect 672 9378 20328 9395
rect 9143 9337 9169 9343
rect 7233 9311 7239 9337
rect 7265 9311 7271 9337
rect 8801 9311 8807 9337
rect 8833 9311 8839 9337
rect 9143 9305 9169 9311
rect 9255 9337 9281 9343
rect 9255 9305 9281 9311
rect 11215 9337 11241 9343
rect 11215 9305 11241 9311
rect 9759 9281 9785 9287
rect 9585 9255 9591 9281
rect 9617 9255 9623 9281
rect 9921 9255 9927 9281
rect 9953 9255 9959 9281
rect 10705 9255 10711 9281
rect 10737 9255 10743 9281
rect 11041 9255 11047 9281
rect 11073 9255 11079 9281
rect 11993 9255 11999 9281
rect 12025 9255 12031 9281
rect 13505 9255 13511 9281
rect 13537 9255 13543 9281
rect 9759 9249 9785 9255
rect 7015 9225 7041 9231
rect 6505 9199 6511 9225
rect 6537 9199 6543 9225
rect 6897 9199 6903 9225
rect 6929 9199 6935 9225
rect 7015 9193 7041 9199
rect 7239 9225 7265 9231
rect 7239 9193 7265 9199
rect 7295 9225 7321 9231
rect 7295 9193 7321 9199
rect 7519 9225 7545 9231
rect 7519 9193 7545 9199
rect 8975 9225 9001 9231
rect 10095 9225 10121 9231
rect 11383 9225 11409 9231
rect 11831 9225 11857 9231
rect 9417 9199 9423 9225
rect 9449 9199 9455 9225
rect 10817 9199 10823 9225
rect 10849 9199 10855 9225
rect 11601 9199 11607 9225
rect 11633 9199 11639 9225
rect 13113 9199 13119 9225
rect 13145 9199 13151 9225
rect 8975 9193 9001 9199
rect 10095 9193 10121 9199
rect 11383 9193 11409 9199
rect 11831 9193 11857 9199
rect 7407 9169 7433 9175
rect 5441 9143 5447 9169
rect 5473 9143 5479 9169
rect 7407 9137 7433 9143
rect 7743 9169 7769 9175
rect 7743 9137 7769 9143
rect 9199 9169 9225 9175
rect 9199 9137 9225 9143
rect 12951 9169 12977 9175
rect 14569 9143 14575 9169
rect 14601 9143 14607 9169
rect 12951 9137 12977 9143
rect 672 9029 20328 9046
rect 672 9003 2239 9029
rect 2265 9003 2291 9029
rect 2317 9003 2343 9029
rect 2369 9003 17599 9029
rect 17625 9003 17651 9029
rect 17677 9003 17703 9029
rect 17729 9003 20328 9029
rect 672 8986 20328 9003
rect 6791 8945 6817 8951
rect 6791 8913 6817 8919
rect 7519 8945 7545 8951
rect 7519 8913 7545 8919
rect 8975 8945 9001 8951
rect 8975 8913 9001 8919
rect 967 8889 993 8895
rect 20007 8889 20033 8895
rect 8409 8863 8415 8889
rect 8441 8863 8447 8889
rect 8857 8863 8863 8889
rect 8889 8863 8895 8889
rect 9361 8863 9367 8889
rect 9393 8863 9399 8889
rect 11097 8863 11103 8889
rect 11129 8863 11135 8889
rect 967 8857 993 8863
rect 20007 8857 20033 8863
rect 6847 8833 6873 8839
rect 2137 8807 2143 8833
rect 2169 8807 2175 8833
rect 6847 8801 6873 8807
rect 7015 8833 7041 8839
rect 7015 8801 7041 8807
rect 7127 8833 7153 8839
rect 7127 8801 7153 8807
rect 7239 8833 7265 8839
rect 7239 8801 7265 8807
rect 7351 8833 7377 8839
rect 7351 8801 7377 8807
rect 8695 8833 8721 8839
rect 11999 8833 12025 8839
rect 8801 8807 8807 8833
rect 8833 8807 8839 8833
rect 9249 8807 9255 8833
rect 9281 8807 9287 8833
rect 9697 8807 9703 8833
rect 9729 8807 9735 8833
rect 10985 8807 10991 8833
rect 11017 8807 11023 8833
rect 11657 8807 11663 8833
rect 11689 8807 11695 8833
rect 18937 8807 18943 8833
rect 18969 8807 18975 8833
rect 8695 8801 8721 8807
rect 11999 8801 12025 8807
rect 6791 8777 6817 8783
rect 6791 8745 6817 8751
rect 7575 8777 7601 8783
rect 10655 8777 10681 8783
rect 11943 8777 11969 8783
rect 9473 8751 9479 8777
rect 9505 8751 9511 8777
rect 11545 8751 11551 8777
rect 11577 8751 11583 8777
rect 7575 8745 7601 8751
rect 10655 8745 10681 8751
rect 11943 8745 11969 8751
rect 7407 8721 7433 8727
rect 7407 8689 7433 8695
rect 8415 8721 8441 8727
rect 8415 8689 8441 8695
rect 8527 8721 8553 8727
rect 8527 8689 8553 8695
rect 11831 8721 11857 8727
rect 11831 8689 11857 8695
rect 672 8637 20328 8654
rect 672 8611 9919 8637
rect 9945 8611 9971 8637
rect 9997 8611 10023 8637
rect 10049 8611 20328 8637
rect 672 8594 20328 8611
rect 7743 8553 7769 8559
rect 7743 8521 7769 8527
rect 7855 8553 7881 8559
rect 7855 8521 7881 8527
rect 9087 8553 9113 8559
rect 9087 8521 9113 8527
rect 9199 8553 9225 8559
rect 9199 8521 9225 8527
rect 12615 8553 12641 8559
rect 12615 8521 12641 8527
rect 12839 8553 12865 8559
rect 12839 8521 12865 8527
rect 12727 8497 12753 8503
rect 6505 8471 6511 8497
rect 6537 8471 6543 8497
rect 13673 8471 13679 8497
rect 13705 8471 13711 8497
rect 12727 8465 12753 8471
rect 8079 8441 8105 8447
rect 2137 8415 2143 8441
rect 2169 8415 2175 8441
rect 6897 8415 6903 8441
rect 6929 8415 6935 8441
rect 8079 8409 8105 8415
rect 8863 8441 8889 8447
rect 13119 8441 13145 8447
rect 9585 8415 9591 8441
rect 9617 8415 9623 8441
rect 13561 8415 13567 8441
rect 13593 8415 13599 8441
rect 18825 8415 18831 8441
rect 18857 8415 18863 8441
rect 8863 8409 8889 8415
rect 13119 8409 13145 8415
rect 967 8385 993 8391
rect 7127 8385 7153 8391
rect 5441 8359 5447 8385
rect 5473 8359 5479 8385
rect 967 8353 993 8359
rect 7127 8353 7153 8359
rect 7799 8385 7825 8391
rect 7799 8353 7825 8359
rect 8975 8385 9001 8391
rect 8975 8353 9001 8359
rect 9143 8385 9169 8391
rect 12671 8385 12697 8391
rect 10649 8359 10655 8385
rect 10681 8359 10687 8385
rect 19945 8359 19951 8385
rect 19977 8359 19983 8385
rect 9143 8353 9169 8359
rect 12671 8353 12697 8359
rect 13063 8329 13089 8335
rect 13063 8297 13089 8303
rect 672 8245 20328 8262
rect 672 8219 2239 8245
rect 2265 8219 2291 8245
rect 2317 8219 2343 8245
rect 2369 8219 17599 8245
rect 17625 8219 17651 8245
rect 17677 8219 17703 8245
rect 17729 8219 20328 8245
rect 672 8202 20328 8219
rect 9423 8161 9449 8167
rect 9423 8129 9449 8135
rect 9591 8161 9617 8167
rect 9591 8129 9617 8135
rect 10711 8161 10737 8167
rect 10711 8129 10737 8135
rect 10823 8161 10849 8167
rect 10823 8129 10849 8135
rect 12167 8161 12193 8167
rect 12167 8129 12193 8135
rect 12335 8161 12361 8167
rect 12335 8129 12361 8135
rect 10935 8105 10961 8111
rect 8409 8079 8415 8105
rect 8441 8079 8447 8105
rect 10935 8073 10961 8079
rect 11887 8105 11913 8111
rect 11887 8073 11913 8079
rect 12055 8105 12081 8111
rect 20007 8105 20033 8111
rect 14065 8079 14071 8105
rect 14097 8079 14103 8105
rect 12055 8073 12081 8079
rect 20007 8073 20033 8079
rect 8695 8049 8721 8055
rect 8521 8023 8527 8049
rect 8553 8023 8559 8049
rect 8695 8017 8721 8023
rect 11383 8049 11409 8055
rect 12553 8023 12559 8049
rect 12585 8023 12591 8049
rect 18825 8023 18831 8049
rect 18857 8023 18863 8049
rect 11383 8017 11409 8023
rect 11439 7993 11465 7999
rect 11439 7961 11465 7967
rect 11551 7993 11577 7999
rect 12945 7967 12951 7993
rect 12977 7967 12983 7993
rect 11551 7961 11577 7967
rect 8415 7937 8441 7943
rect 8415 7905 8441 7911
rect 8863 7937 8889 7943
rect 8863 7905 8889 7911
rect 9479 7937 9505 7943
rect 9479 7905 9505 7911
rect 11047 7937 11073 7943
rect 11047 7905 11073 7911
rect 11103 7937 11129 7943
rect 11103 7905 11129 7911
rect 11159 7937 11185 7943
rect 11159 7905 11185 7911
rect 672 7853 20328 7870
rect 672 7827 9919 7853
rect 9945 7827 9971 7853
rect 9997 7827 10023 7853
rect 10049 7827 20328 7853
rect 672 7810 20328 7827
rect 11327 7769 11353 7775
rect 11327 7737 11353 7743
rect 12223 7769 12249 7775
rect 12223 7737 12249 7743
rect 11607 7713 11633 7719
rect 7345 7687 7351 7713
rect 7377 7687 7383 7713
rect 9081 7687 9087 7713
rect 9113 7687 9119 7713
rect 13673 7687 13679 7713
rect 13705 7687 13711 7713
rect 11607 7681 11633 7687
rect 7009 7631 7015 7657
rect 7041 7631 7047 7657
rect 8745 7631 8751 7657
rect 8777 7631 8783 7657
rect 11433 7631 11439 7657
rect 11465 7631 11471 7657
rect 11769 7631 11775 7657
rect 11801 7631 11807 7657
rect 13561 7631 13567 7657
rect 13593 7631 13599 7657
rect 10375 7601 10401 7607
rect 8409 7575 8415 7601
rect 8441 7575 8447 7601
rect 10145 7575 10151 7601
rect 10177 7575 10183 7601
rect 10375 7569 10401 7575
rect 11271 7601 11297 7607
rect 11271 7569 11297 7575
rect 11663 7601 11689 7607
rect 11663 7569 11689 7575
rect 672 7461 20328 7478
rect 672 7435 2239 7461
rect 2265 7435 2291 7461
rect 2317 7435 2343 7461
rect 2369 7435 17599 7461
rect 17625 7435 17651 7461
rect 17677 7435 17703 7461
rect 17729 7435 20328 7461
rect 672 7418 20328 7435
rect 12279 7377 12305 7383
rect 12279 7345 12305 7351
rect 8639 7321 8665 7327
rect 12335 7321 12361 7327
rect 8857 7295 8863 7321
rect 8889 7295 8895 7321
rect 11041 7295 11047 7321
rect 11073 7295 11079 7321
rect 12105 7295 12111 7321
rect 12137 7295 12143 7321
rect 8639 7289 8665 7295
rect 12335 7289 12361 7295
rect 9255 7265 9281 7271
rect 8913 7239 8919 7265
rect 8945 7239 8951 7265
rect 9025 7239 9031 7265
rect 9057 7239 9063 7265
rect 10649 7239 10655 7265
rect 10681 7239 10687 7265
rect 9255 7233 9281 7239
rect 8583 7153 8609 7159
rect 8583 7121 8609 7127
rect 9143 7153 9169 7159
rect 9143 7121 9169 7127
rect 12391 7153 12417 7159
rect 12391 7121 12417 7127
rect 12615 7153 12641 7159
rect 12777 7127 12783 7153
rect 12809 7127 12815 7153
rect 12615 7121 12641 7127
rect 672 7069 20328 7086
rect 672 7043 9919 7069
rect 9945 7043 9971 7069
rect 9997 7043 10023 7069
rect 10049 7043 20328 7069
rect 672 7026 20328 7043
rect 12671 6985 12697 6991
rect 12671 6953 12697 6959
rect 11265 6903 11271 6929
rect 11297 6903 11303 6929
rect 10873 6847 10879 6873
rect 10905 6847 10911 6873
rect 12329 6791 12335 6817
rect 12361 6791 12367 6817
rect 672 6677 20328 6694
rect 672 6651 2239 6677
rect 2265 6651 2291 6677
rect 2317 6651 2343 6677
rect 2369 6651 17599 6677
rect 17625 6651 17651 6677
rect 17677 6651 17703 6677
rect 17729 6651 20328 6677
rect 672 6634 20328 6651
rect 8129 6511 8135 6537
rect 8161 6511 8167 6537
rect 9193 6511 9199 6537
rect 9225 6511 9231 6537
rect 9479 6481 9505 6487
rect 7793 6455 7799 6481
rect 7825 6455 7831 6481
rect 9479 6449 9505 6455
rect 672 6285 20328 6302
rect 672 6259 9919 6285
rect 9945 6259 9971 6285
rect 9997 6259 10023 6285
rect 10049 6259 20328 6285
rect 672 6242 20328 6259
rect 672 5893 20328 5910
rect 672 5867 2239 5893
rect 2265 5867 2291 5893
rect 2317 5867 2343 5893
rect 2369 5867 17599 5893
rect 17625 5867 17651 5893
rect 17677 5867 17703 5893
rect 17729 5867 20328 5893
rect 672 5850 20328 5867
rect 672 5501 20328 5518
rect 672 5475 9919 5501
rect 9945 5475 9971 5501
rect 9997 5475 10023 5501
rect 10049 5475 20328 5501
rect 672 5458 20328 5475
rect 672 5109 20328 5126
rect 672 5083 2239 5109
rect 2265 5083 2291 5109
rect 2317 5083 2343 5109
rect 2369 5083 17599 5109
rect 17625 5083 17651 5109
rect 17677 5083 17703 5109
rect 17729 5083 20328 5109
rect 672 5066 20328 5083
rect 672 4717 20328 4734
rect 672 4691 9919 4717
rect 9945 4691 9971 4717
rect 9997 4691 10023 4717
rect 10049 4691 20328 4717
rect 672 4674 20328 4691
rect 672 4325 20328 4342
rect 672 4299 2239 4325
rect 2265 4299 2291 4325
rect 2317 4299 2343 4325
rect 2369 4299 17599 4325
rect 17625 4299 17651 4325
rect 17677 4299 17703 4325
rect 17729 4299 20328 4325
rect 672 4282 20328 4299
rect 672 3933 20328 3950
rect 672 3907 9919 3933
rect 9945 3907 9971 3933
rect 9997 3907 10023 3933
rect 10049 3907 20328 3933
rect 672 3890 20328 3907
rect 672 3541 20328 3558
rect 672 3515 2239 3541
rect 2265 3515 2291 3541
rect 2317 3515 2343 3541
rect 2369 3515 17599 3541
rect 17625 3515 17651 3541
rect 17677 3515 17703 3541
rect 17729 3515 20328 3541
rect 672 3498 20328 3515
rect 672 3149 20328 3166
rect 672 3123 9919 3149
rect 9945 3123 9971 3149
rect 9997 3123 10023 3149
rect 10049 3123 20328 3149
rect 672 3106 20328 3123
rect 672 2757 20328 2774
rect 672 2731 2239 2757
rect 2265 2731 2291 2757
rect 2317 2731 2343 2757
rect 2369 2731 17599 2757
rect 17625 2731 17651 2757
rect 17677 2731 17703 2757
rect 17729 2731 20328 2757
rect 672 2714 20328 2731
rect 11999 2617 12025 2623
rect 11999 2585 12025 2591
rect 12945 2535 12951 2561
rect 12977 2535 12983 2561
rect 672 2365 20328 2382
rect 672 2339 9919 2365
rect 9945 2339 9971 2365
rect 9997 2339 10023 2365
rect 10049 2339 20328 2365
rect 672 2322 20328 2339
rect 8689 2143 8695 2169
rect 8721 2143 8727 2169
rect 12609 2143 12615 2169
rect 12641 2143 12647 2169
rect 9199 2057 9225 2063
rect 9199 2025 9225 2031
rect 13119 2057 13145 2063
rect 13119 2025 13145 2031
rect 672 1973 20328 1990
rect 672 1947 2239 1973
rect 2265 1947 2291 1973
rect 2317 1947 2343 1973
rect 2369 1947 17599 1973
rect 17625 1947 17651 1973
rect 17677 1947 17703 1973
rect 17729 1947 20328 1973
rect 672 1930 20328 1947
rect 9311 1833 9337 1839
rect 12783 1833 12809 1839
rect 10929 1807 10935 1833
rect 10961 1807 10967 1833
rect 9311 1801 9337 1807
rect 12783 1801 12809 1807
rect 8801 1751 8807 1777
rect 8833 1751 8839 1777
rect 10369 1751 10375 1777
rect 10401 1751 10407 1777
rect 12273 1751 12279 1777
rect 12305 1751 12311 1777
rect 672 1581 20328 1598
rect 672 1555 9919 1581
rect 9945 1555 9971 1581
rect 9997 1555 10023 1581
rect 10049 1555 20328 1581
rect 672 1538 20328 1555
<< via1 >>
rect 2239 19195 2265 19221
rect 2291 19195 2317 19221
rect 2343 19195 2369 19221
rect 17599 19195 17625 19221
rect 17651 19195 17677 19221
rect 17703 19195 17729 19221
rect 9311 19111 9337 19137
rect 11215 19111 11241 19137
rect 13063 19111 13089 19137
rect 8975 18999 9001 19025
rect 10711 18999 10737 19025
rect 12671 18999 12697 19025
rect 9919 18803 9945 18829
rect 9971 18803 9997 18829
rect 10023 18803 10049 18829
rect 9367 18719 9393 18745
rect 11383 18719 11409 18745
rect 9031 18607 9057 18633
rect 10991 18607 11017 18633
rect 2239 18411 2265 18437
rect 2291 18411 2317 18437
rect 2343 18411 2369 18437
rect 17599 18411 17625 18437
rect 17651 18411 17677 18437
rect 17703 18411 17729 18437
rect 8639 18327 8665 18353
rect 9591 18215 9617 18241
rect 9919 18019 9945 18045
rect 9971 18019 9997 18045
rect 10023 18019 10049 18045
rect 2239 17627 2265 17653
rect 2291 17627 2317 17653
rect 2343 17627 2369 17653
rect 17599 17627 17625 17653
rect 17651 17627 17677 17653
rect 17703 17627 17729 17653
rect 9919 17235 9945 17261
rect 9971 17235 9997 17261
rect 10023 17235 10049 17261
rect 2239 16843 2265 16869
rect 2291 16843 2317 16869
rect 2343 16843 2369 16869
rect 17599 16843 17625 16869
rect 17651 16843 17677 16869
rect 17703 16843 17729 16869
rect 9919 16451 9945 16477
rect 9971 16451 9997 16477
rect 10023 16451 10049 16477
rect 2239 16059 2265 16085
rect 2291 16059 2317 16085
rect 2343 16059 2369 16085
rect 17599 16059 17625 16085
rect 17651 16059 17677 16085
rect 17703 16059 17729 16085
rect 9919 15667 9945 15693
rect 9971 15667 9997 15693
rect 10023 15667 10049 15693
rect 2239 15275 2265 15301
rect 2291 15275 2317 15301
rect 2343 15275 2369 15301
rect 17599 15275 17625 15301
rect 17651 15275 17677 15301
rect 17703 15275 17729 15301
rect 9919 14883 9945 14909
rect 9971 14883 9997 14909
rect 10023 14883 10049 14909
rect 9591 14687 9617 14713
rect 9983 14631 10009 14657
rect 11047 14631 11073 14657
rect 11327 14631 11353 14657
rect 2239 14491 2265 14517
rect 2291 14491 2317 14517
rect 2343 14491 2369 14517
rect 17599 14491 17625 14517
rect 17651 14491 17677 14517
rect 17703 14491 17729 14517
rect 8527 14295 8553 14321
rect 9919 14099 9945 14125
rect 9971 14099 9997 14125
rect 10023 14099 10049 14125
rect 8863 14015 8889 14041
rect 9031 14015 9057 14041
rect 11215 14015 11241 14041
rect 7015 13903 7041 13929
rect 9591 13903 9617 13929
rect 7351 13847 7377 13873
rect 8415 13847 8441 13873
rect 9927 13847 9953 13873
rect 10991 13847 11017 13873
rect 2239 13707 2265 13733
rect 2291 13707 2317 13733
rect 2343 13707 2369 13733
rect 17599 13707 17625 13733
rect 17651 13707 17677 13733
rect 17703 13707 17729 13733
rect 10711 13623 10737 13649
rect 967 13567 993 13593
rect 9087 13567 9113 13593
rect 9591 13567 9617 13593
rect 20007 13567 20033 13593
rect 2143 13511 2169 13537
rect 7687 13511 7713 13537
rect 10151 13511 10177 13537
rect 10319 13511 10345 13537
rect 18943 13511 18969 13537
rect 8023 13455 8049 13481
rect 9199 13455 9225 13481
rect 9311 13455 9337 13481
rect 9367 13455 9393 13481
rect 10655 13455 10681 13481
rect 10711 13455 10737 13481
rect 10263 13399 10289 13425
rect 9919 13315 9945 13341
rect 9971 13315 9997 13341
rect 10023 13315 10049 13341
rect 7967 13231 7993 13257
rect 8247 13231 8273 13257
rect 8751 13231 8777 13257
rect 10655 13231 10681 13257
rect 8079 13175 8105 13201
rect 8135 13175 8161 13201
rect 8359 13175 8385 13201
rect 9927 13175 9953 13201
rect 10543 13175 10569 13201
rect 12671 13175 12697 13201
rect 13567 13175 13593 13201
rect 7687 13119 7713 13145
rect 8415 13119 8441 13145
rect 8639 13119 8665 13145
rect 8807 13119 8833 13145
rect 9871 13119 9897 13145
rect 10711 13119 10737 13145
rect 10935 13119 10961 13145
rect 12727 13119 12753 13145
rect 13511 13119 13537 13145
rect 18831 13119 18857 13145
rect 6287 13063 6313 13089
rect 7351 13063 7377 13089
rect 11271 13063 11297 13089
rect 12335 13063 12361 13089
rect 12951 13063 12977 13089
rect 14519 13063 14545 13089
rect 9927 13007 9953 13033
rect 12671 13007 12697 13033
rect 13567 13007 13593 13033
rect 14463 13007 14489 13033
rect 20007 13007 20033 13033
rect 2239 12923 2265 12949
rect 2291 12923 2317 12949
rect 2343 12923 2369 12949
rect 17599 12923 17625 12949
rect 17651 12923 17677 12949
rect 17703 12923 17729 12949
rect 7687 12783 7713 12809
rect 7855 12783 7881 12809
rect 8247 12783 8273 12809
rect 11775 12783 11801 12809
rect 14071 12783 14097 12809
rect 7911 12727 7937 12753
rect 8191 12727 8217 12753
rect 8359 12727 8385 12753
rect 12055 12727 12081 12753
rect 12447 12727 12473 12753
rect 12671 12727 12697 12753
rect 10207 12671 10233 12697
rect 13007 12671 13033 12697
rect 8135 12615 8161 12641
rect 8303 12615 8329 12641
rect 10375 12615 10401 12641
rect 10767 12615 10793 12641
rect 10935 12615 10961 12641
rect 11719 12615 11745 12641
rect 11831 12615 11857 12641
rect 9919 12531 9945 12557
rect 9971 12531 9997 12557
rect 10023 12531 10049 12557
rect 8359 12447 8385 12473
rect 12895 12447 12921 12473
rect 13343 12447 13369 12473
rect 8191 12335 8217 12361
rect 9815 12335 9841 12361
rect 12839 12335 12865 12361
rect 12951 12335 12977 12361
rect 13175 12335 13201 12361
rect 13511 12335 13537 12361
rect 8079 12279 8105 12305
rect 8807 12279 8833 12305
rect 10487 12279 10513 12305
rect 13903 12279 13929 12305
rect 14967 12279 14993 12305
rect 2239 12139 2265 12165
rect 2291 12139 2317 12165
rect 2343 12139 2369 12165
rect 17599 12139 17625 12165
rect 17651 12139 17677 12165
rect 17703 12139 17729 12165
rect 8863 12055 8889 12081
rect 967 11999 993 12025
rect 6735 11999 6761 12025
rect 9143 11999 9169 12025
rect 10823 11999 10849 12025
rect 2143 11943 2169 11969
rect 8191 11943 8217 11969
rect 8583 11943 8609 11969
rect 8751 11943 8777 11969
rect 9367 11943 9393 11969
rect 10151 11943 10177 11969
rect 13343 11943 13369 11969
rect 13623 11943 13649 11969
rect 13735 11943 13761 11969
rect 13903 11943 13929 11969
rect 14183 11943 14209 11969
rect 7799 11887 7825 11913
rect 8471 11887 8497 11913
rect 9983 11887 10009 11913
rect 13399 11887 13425 11913
rect 8415 11831 8441 11857
rect 8527 11831 8553 11857
rect 9087 11831 9113 11857
rect 9199 11831 9225 11857
rect 10039 11831 10065 11857
rect 13511 11831 13537 11857
rect 14071 11831 14097 11857
rect 9919 11747 9945 11773
rect 9971 11747 9997 11773
rect 10023 11747 10049 11773
rect 8079 11663 8105 11689
rect 12671 11663 12697 11689
rect 5895 11607 5921 11633
rect 8975 11607 9001 11633
rect 9031 11607 9057 11633
rect 5559 11551 5585 11577
rect 7183 11551 7209 11577
rect 8023 11551 8049 11577
rect 8359 11551 8385 11577
rect 9255 11551 9281 11577
rect 10935 11551 10961 11577
rect 13623 11551 13649 11577
rect 6959 11495 6985 11521
rect 9647 11495 9673 11521
rect 10711 11495 10737 11521
rect 11271 11495 11297 11521
rect 12335 11495 12361 11521
rect 13735 11495 13761 11521
rect 8079 11439 8105 11465
rect 8975 11439 9001 11465
rect 13791 11439 13817 11465
rect 2239 11355 2265 11381
rect 2291 11355 2317 11381
rect 2343 11355 2369 11381
rect 17599 11355 17625 11381
rect 17651 11355 17677 11381
rect 17703 11355 17729 11381
rect 9479 11271 9505 11297
rect 10879 11215 10905 11241
rect 11495 11215 11521 11241
rect 12895 11215 12921 11241
rect 13959 11215 13985 11241
rect 20007 11215 20033 11241
rect 7743 11159 7769 11185
rect 8247 11159 8273 11185
rect 8471 11159 8497 11185
rect 8807 11159 8833 11185
rect 8919 11159 8945 11185
rect 9423 11159 9449 11185
rect 10599 11159 10625 11185
rect 10935 11159 10961 11185
rect 11103 11159 11129 11185
rect 11439 11159 11465 11185
rect 11607 11159 11633 11185
rect 12055 11159 12081 11185
rect 12727 11159 12753 11185
rect 14071 11159 14097 11185
rect 18831 11159 18857 11185
rect 7855 11103 7881 11129
rect 9927 11103 9953 11129
rect 10151 11103 10177 11129
rect 10319 11103 10345 11129
rect 11215 11103 11241 11129
rect 11719 11103 11745 11129
rect 11887 11103 11913 11129
rect 12895 11103 12921 11129
rect 12951 11103 12977 11129
rect 13903 11103 13929 11129
rect 9087 11047 9113 11073
rect 9479 11047 9505 11073
rect 9759 11047 9785 11073
rect 10095 11047 10121 11073
rect 10207 11047 10233 11073
rect 10823 11047 10849 11073
rect 11159 11047 11185 11073
rect 12839 11047 12865 11073
rect 9919 10963 9945 10989
rect 9971 10963 9997 10989
rect 10023 10963 10049 10989
rect 12783 10879 12809 10905
rect 13175 10879 13201 10905
rect 8415 10823 8441 10849
rect 8695 10823 8721 10849
rect 12671 10823 12697 10849
rect 13735 10823 13761 10849
rect 5839 10767 5865 10793
rect 7687 10767 7713 10793
rect 7855 10767 7881 10793
rect 8303 10767 8329 10793
rect 8807 10767 8833 10793
rect 9479 10767 9505 10793
rect 9703 10767 9729 10793
rect 12615 10767 12641 10793
rect 13343 10767 13369 10793
rect 6175 10711 6201 10737
rect 7239 10711 7265 10737
rect 7407 10711 7433 10737
rect 10935 10711 10961 10737
rect 14799 10711 14825 10737
rect 8975 10655 9001 10681
rect 2239 10571 2265 10597
rect 2291 10571 2317 10597
rect 2343 10571 2369 10597
rect 17599 10571 17625 10597
rect 17651 10571 17677 10597
rect 17703 10571 17729 10597
rect 7407 10431 7433 10457
rect 8863 10431 8889 10457
rect 11383 10431 11409 10457
rect 12895 10431 12921 10457
rect 20007 10431 20033 10457
rect 7015 10375 7041 10401
rect 9143 10375 9169 10401
rect 9311 10375 9337 10401
rect 9927 10375 9953 10401
rect 11103 10375 11129 10401
rect 11887 10375 11913 10401
rect 12727 10375 12753 10401
rect 12951 10375 12977 10401
rect 13119 10375 13145 10401
rect 18943 10375 18969 10401
rect 6847 10319 6873 10345
rect 8863 10319 8889 10345
rect 9423 10319 9449 10345
rect 12839 10319 12865 10345
rect 8975 10263 9001 10289
rect 10095 10263 10121 10289
rect 11775 10263 11801 10289
rect 9919 10179 9945 10205
rect 9971 10179 9997 10205
rect 10023 10179 10049 10205
rect 8415 10095 8441 10121
rect 7631 10039 7657 10065
rect 8247 10039 8273 10065
rect 9815 10039 9841 10065
rect 10263 10039 10289 10065
rect 11383 10039 11409 10065
rect 11663 10039 11689 10065
rect 11943 10039 11969 10065
rect 13287 10039 13313 10065
rect 14687 10039 14713 10065
rect 2143 9983 2169 10009
rect 7071 9983 7097 10009
rect 7183 9983 7209 10009
rect 7295 9983 7321 10009
rect 7407 9983 7433 10009
rect 7519 9983 7545 10009
rect 7687 9983 7713 10009
rect 8919 9983 8945 10009
rect 9479 9983 9505 10009
rect 11047 9983 11073 10009
rect 11271 9983 11297 10009
rect 11607 9983 11633 10009
rect 12951 9983 12977 10009
rect 14575 9983 14601 10009
rect 18831 9983 18857 10009
rect 7015 9927 7041 9953
rect 7911 9927 7937 9953
rect 9031 9927 9057 9953
rect 10879 9927 10905 9953
rect 12783 9927 12809 9953
rect 14351 9927 14377 9953
rect 967 9871 993 9897
rect 11439 9871 11465 9897
rect 20007 9871 20033 9897
rect 2239 9787 2265 9813
rect 2291 9787 2317 9813
rect 2343 9787 2369 9813
rect 17599 9787 17625 9813
rect 17651 9787 17677 9813
rect 17703 9787 17729 9813
rect 7295 9703 7321 9729
rect 9759 9703 9785 9729
rect 10655 9703 10681 9729
rect 4999 9647 5025 9673
rect 6063 9647 6089 9673
rect 8695 9647 8721 9673
rect 10767 9647 10793 9673
rect 12055 9647 12081 9673
rect 13455 9647 13481 9673
rect 20007 9647 20033 9673
rect 6455 9591 6481 9617
rect 7071 9591 7097 9617
rect 8023 9591 8049 9617
rect 8303 9591 8329 9617
rect 8583 9591 8609 9617
rect 9031 9591 9057 9617
rect 10823 9591 10849 9617
rect 11607 9591 11633 9617
rect 11831 9591 11857 9617
rect 13231 9591 13257 9617
rect 13399 9591 13425 9617
rect 13511 9591 13537 9617
rect 13791 9591 13817 9617
rect 14071 9591 14097 9617
rect 18831 9591 18857 9617
rect 7015 9535 7041 9561
rect 7295 9535 7321 9561
rect 7351 9535 7377 9561
rect 7855 9535 7881 9561
rect 8863 9535 8889 9561
rect 9311 9535 9337 9561
rect 9479 9535 9505 9561
rect 14015 9535 14041 9561
rect 14575 9535 14601 9561
rect 14743 9535 14769 9561
rect 6791 9479 6817 9505
rect 6903 9479 6929 9505
rect 8135 9479 8161 9505
rect 8247 9479 8273 9505
rect 8751 9479 8777 9505
rect 9087 9479 9113 9505
rect 9815 9479 9841 9505
rect 9871 9479 9897 9505
rect 10991 9479 11017 9505
rect 11159 9479 11185 9505
rect 11439 9479 11465 9505
rect 11775 9479 11801 9505
rect 11999 9479 12025 9505
rect 13623 9479 13649 9505
rect 13903 9479 13929 9505
rect 14631 9479 14657 9505
rect 9919 9395 9945 9421
rect 9971 9395 9997 9421
rect 10023 9395 10049 9421
rect 7239 9311 7265 9337
rect 8807 9311 8833 9337
rect 9143 9311 9169 9337
rect 9255 9311 9281 9337
rect 11215 9311 11241 9337
rect 9591 9255 9617 9281
rect 9759 9255 9785 9281
rect 9927 9255 9953 9281
rect 10711 9255 10737 9281
rect 11047 9255 11073 9281
rect 11999 9255 12025 9281
rect 13511 9255 13537 9281
rect 6511 9199 6537 9225
rect 6903 9199 6929 9225
rect 7015 9199 7041 9225
rect 7239 9199 7265 9225
rect 7295 9199 7321 9225
rect 7519 9199 7545 9225
rect 8975 9199 9001 9225
rect 9423 9199 9449 9225
rect 10095 9199 10121 9225
rect 10823 9199 10849 9225
rect 11383 9199 11409 9225
rect 11607 9199 11633 9225
rect 11831 9199 11857 9225
rect 13119 9199 13145 9225
rect 5447 9143 5473 9169
rect 7407 9143 7433 9169
rect 7743 9143 7769 9169
rect 9199 9143 9225 9169
rect 12951 9143 12977 9169
rect 14575 9143 14601 9169
rect 2239 9003 2265 9029
rect 2291 9003 2317 9029
rect 2343 9003 2369 9029
rect 17599 9003 17625 9029
rect 17651 9003 17677 9029
rect 17703 9003 17729 9029
rect 6791 8919 6817 8945
rect 7519 8919 7545 8945
rect 8975 8919 9001 8945
rect 967 8863 993 8889
rect 8415 8863 8441 8889
rect 8863 8863 8889 8889
rect 9367 8863 9393 8889
rect 11103 8863 11129 8889
rect 20007 8863 20033 8889
rect 2143 8807 2169 8833
rect 6847 8807 6873 8833
rect 7015 8807 7041 8833
rect 7127 8807 7153 8833
rect 7239 8807 7265 8833
rect 7351 8807 7377 8833
rect 8695 8807 8721 8833
rect 8807 8807 8833 8833
rect 9255 8807 9281 8833
rect 9703 8807 9729 8833
rect 10991 8807 11017 8833
rect 11663 8807 11689 8833
rect 11999 8807 12025 8833
rect 18943 8807 18969 8833
rect 6791 8751 6817 8777
rect 7575 8751 7601 8777
rect 9479 8751 9505 8777
rect 10655 8751 10681 8777
rect 11551 8751 11577 8777
rect 11943 8751 11969 8777
rect 7407 8695 7433 8721
rect 8415 8695 8441 8721
rect 8527 8695 8553 8721
rect 11831 8695 11857 8721
rect 9919 8611 9945 8637
rect 9971 8611 9997 8637
rect 10023 8611 10049 8637
rect 7743 8527 7769 8553
rect 7855 8527 7881 8553
rect 9087 8527 9113 8553
rect 9199 8527 9225 8553
rect 12615 8527 12641 8553
rect 12839 8527 12865 8553
rect 6511 8471 6537 8497
rect 12727 8471 12753 8497
rect 13679 8471 13705 8497
rect 2143 8415 2169 8441
rect 6903 8415 6929 8441
rect 8079 8415 8105 8441
rect 8863 8415 8889 8441
rect 9591 8415 9617 8441
rect 13119 8415 13145 8441
rect 13567 8415 13593 8441
rect 18831 8415 18857 8441
rect 967 8359 993 8385
rect 5447 8359 5473 8385
rect 7127 8359 7153 8385
rect 7799 8359 7825 8385
rect 8975 8359 9001 8385
rect 9143 8359 9169 8385
rect 10655 8359 10681 8385
rect 12671 8359 12697 8385
rect 19951 8359 19977 8385
rect 13063 8303 13089 8329
rect 2239 8219 2265 8245
rect 2291 8219 2317 8245
rect 2343 8219 2369 8245
rect 17599 8219 17625 8245
rect 17651 8219 17677 8245
rect 17703 8219 17729 8245
rect 9423 8135 9449 8161
rect 9591 8135 9617 8161
rect 10711 8135 10737 8161
rect 10823 8135 10849 8161
rect 12167 8135 12193 8161
rect 12335 8135 12361 8161
rect 8415 8079 8441 8105
rect 10935 8079 10961 8105
rect 11887 8079 11913 8105
rect 12055 8079 12081 8105
rect 14071 8079 14097 8105
rect 20007 8079 20033 8105
rect 8527 8023 8553 8049
rect 8695 8023 8721 8049
rect 11383 8023 11409 8049
rect 12559 8023 12585 8049
rect 18831 8023 18857 8049
rect 11439 7967 11465 7993
rect 11551 7967 11577 7993
rect 12951 7967 12977 7993
rect 8415 7911 8441 7937
rect 8863 7911 8889 7937
rect 9479 7911 9505 7937
rect 11047 7911 11073 7937
rect 11103 7911 11129 7937
rect 11159 7911 11185 7937
rect 9919 7827 9945 7853
rect 9971 7827 9997 7853
rect 10023 7827 10049 7853
rect 11327 7743 11353 7769
rect 12223 7743 12249 7769
rect 7351 7687 7377 7713
rect 9087 7687 9113 7713
rect 11607 7687 11633 7713
rect 13679 7687 13705 7713
rect 7015 7631 7041 7657
rect 8751 7631 8777 7657
rect 11439 7631 11465 7657
rect 11775 7631 11801 7657
rect 13567 7631 13593 7657
rect 8415 7575 8441 7601
rect 10151 7575 10177 7601
rect 10375 7575 10401 7601
rect 11271 7575 11297 7601
rect 11663 7575 11689 7601
rect 2239 7435 2265 7461
rect 2291 7435 2317 7461
rect 2343 7435 2369 7461
rect 17599 7435 17625 7461
rect 17651 7435 17677 7461
rect 17703 7435 17729 7461
rect 12279 7351 12305 7377
rect 8639 7295 8665 7321
rect 8863 7295 8889 7321
rect 11047 7295 11073 7321
rect 12111 7295 12137 7321
rect 12335 7295 12361 7321
rect 8919 7239 8945 7265
rect 9031 7239 9057 7265
rect 9255 7239 9281 7265
rect 10655 7239 10681 7265
rect 8583 7127 8609 7153
rect 9143 7127 9169 7153
rect 12391 7127 12417 7153
rect 12615 7127 12641 7153
rect 12783 7127 12809 7153
rect 9919 7043 9945 7069
rect 9971 7043 9997 7069
rect 10023 7043 10049 7069
rect 12671 6959 12697 6985
rect 11271 6903 11297 6929
rect 10879 6847 10905 6873
rect 12335 6791 12361 6817
rect 2239 6651 2265 6677
rect 2291 6651 2317 6677
rect 2343 6651 2369 6677
rect 17599 6651 17625 6677
rect 17651 6651 17677 6677
rect 17703 6651 17729 6677
rect 8135 6511 8161 6537
rect 9199 6511 9225 6537
rect 7799 6455 7825 6481
rect 9479 6455 9505 6481
rect 9919 6259 9945 6285
rect 9971 6259 9997 6285
rect 10023 6259 10049 6285
rect 2239 5867 2265 5893
rect 2291 5867 2317 5893
rect 2343 5867 2369 5893
rect 17599 5867 17625 5893
rect 17651 5867 17677 5893
rect 17703 5867 17729 5893
rect 9919 5475 9945 5501
rect 9971 5475 9997 5501
rect 10023 5475 10049 5501
rect 2239 5083 2265 5109
rect 2291 5083 2317 5109
rect 2343 5083 2369 5109
rect 17599 5083 17625 5109
rect 17651 5083 17677 5109
rect 17703 5083 17729 5109
rect 9919 4691 9945 4717
rect 9971 4691 9997 4717
rect 10023 4691 10049 4717
rect 2239 4299 2265 4325
rect 2291 4299 2317 4325
rect 2343 4299 2369 4325
rect 17599 4299 17625 4325
rect 17651 4299 17677 4325
rect 17703 4299 17729 4325
rect 9919 3907 9945 3933
rect 9971 3907 9997 3933
rect 10023 3907 10049 3933
rect 2239 3515 2265 3541
rect 2291 3515 2317 3541
rect 2343 3515 2369 3541
rect 17599 3515 17625 3541
rect 17651 3515 17677 3541
rect 17703 3515 17729 3541
rect 9919 3123 9945 3149
rect 9971 3123 9997 3149
rect 10023 3123 10049 3149
rect 2239 2731 2265 2757
rect 2291 2731 2317 2757
rect 2343 2731 2369 2757
rect 17599 2731 17625 2757
rect 17651 2731 17677 2757
rect 17703 2731 17729 2757
rect 11999 2591 12025 2617
rect 12951 2535 12977 2561
rect 9919 2339 9945 2365
rect 9971 2339 9997 2365
rect 10023 2339 10049 2365
rect 8695 2143 8721 2169
rect 12615 2143 12641 2169
rect 9199 2031 9225 2057
rect 13119 2031 13145 2057
rect 2239 1947 2265 1973
rect 2291 1947 2317 1973
rect 2343 1947 2369 1973
rect 17599 1947 17625 1973
rect 17651 1947 17677 1973
rect 17703 1947 17729 1973
rect 9311 1807 9337 1833
rect 10935 1807 10961 1833
rect 12783 1807 12809 1833
rect 8807 1751 8833 1777
rect 10375 1751 10401 1777
rect 12279 1751 12305 1777
rect 9919 1555 9945 1581
rect 9971 1555 9997 1581
rect 10023 1555 10049 1581
<< metal2 >>
rect 8400 20600 8456 21000
rect 8736 20600 8792 21000
rect 9072 20600 9128 21000
rect 10752 20600 10808 21000
rect 11088 20600 11144 21000
rect 12432 20600 12488 21000
rect 8414 19418 8442 20600
rect 8414 19390 8666 19418
rect 2238 19222 2370 19227
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2238 19189 2370 19194
rect 2238 18438 2370 18443
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2238 18405 2370 18410
rect 8638 18353 8666 19390
rect 8750 18746 8778 20600
rect 9086 19138 9114 20600
rect 9310 19138 9338 19143
rect 9086 19137 9338 19138
rect 9086 19111 9311 19137
rect 9337 19111 9338 19137
rect 9086 19110 9338 19111
rect 9310 19105 9338 19110
rect 8750 18713 8778 18718
rect 8974 19025 9002 19031
rect 8974 18999 8975 19025
rect 9001 18999 9002 19025
rect 8638 18327 8639 18353
rect 8665 18327 8666 18353
rect 8638 18321 8666 18327
rect 2238 17654 2370 17659
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2238 17621 2370 17626
rect 2238 16870 2370 16875
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2238 16837 2370 16842
rect 2238 16086 2370 16091
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2238 16053 2370 16058
rect 8974 15974 9002 18999
rect 10710 19025 10738 19031
rect 10710 18999 10711 19025
rect 10737 18999 10738 19025
rect 9918 18830 10050 18835
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 9918 18797 10050 18802
rect 9366 18746 9394 18751
rect 9366 18699 9394 18718
rect 8862 15946 9002 15974
rect 9030 18633 9058 18639
rect 9030 18607 9031 18633
rect 9057 18607 9058 18633
rect 2238 15302 2370 15307
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2238 15269 2370 15274
rect 2238 14518 2370 14523
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2238 14485 2370 14490
rect 8526 14322 8554 14327
rect 8526 14275 8554 14294
rect 7686 14266 7714 14271
rect 7014 13930 7042 13935
rect 7014 13883 7042 13902
rect 7686 13930 7714 14238
rect 8862 14041 8890 15946
rect 8862 14015 8863 14041
rect 8889 14015 8890 14041
rect 8862 14009 8890 14015
rect 9030 14042 9058 18607
rect 9590 18241 9618 18247
rect 9590 18215 9591 18241
rect 9617 18215 9618 18241
rect 9590 15974 9618 18215
rect 9918 18046 10050 18051
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 9918 18013 10050 18018
rect 9918 17262 10050 17267
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 9918 17229 10050 17234
rect 9918 16478 10050 16483
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 9918 16445 10050 16450
rect 9254 15946 9618 15974
rect 9030 14041 9114 14042
rect 9030 14015 9031 14041
rect 9057 14015 9114 14041
rect 9030 14014 9114 14015
rect 9030 14009 9058 14014
rect 7350 13873 7378 13879
rect 7350 13847 7351 13873
rect 7377 13847 7378 13873
rect 2086 13818 2114 13823
rect 966 13593 994 13599
rect 966 13567 967 13593
rect 993 13567 994 13593
rect 966 13146 994 13567
rect 966 13113 994 13118
rect 966 12025 994 12031
rect 966 11999 967 12025
rect 993 11999 994 12025
rect 966 11802 994 11999
rect 966 11769 994 11774
rect 2086 10794 2114 13790
rect 2238 13734 2370 13739
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2238 13701 2370 13706
rect 2142 13538 2170 13543
rect 2142 13491 2170 13510
rect 6286 13538 6314 13543
rect 6286 13090 6314 13510
rect 7350 13258 7378 13847
rect 7350 13225 7378 13230
rect 7686 13537 7714 13902
rect 8414 13874 8442 13879
rect 8414 13827 8442 13846
rect 9086 13594 9114 14014
rect 7686 13511 7687 13537
rect 7713 13511 7714 13537
rect 7686 13145 7714 13511
rect 8750 13593 9114 13594
rect 8750 13567 9087 13593
rect 9113 13567 9114 13593
rect 8750 13566 9114 13567
rect 8022 13482 8050 13487
rect 8022 13481 8274 13482
rect 8022 13455 8023 13481
rect 8049 13455 8274 13481
rect 8022 13454 8274 13455
rect 8022 13449 8050 13454
rect 8134 13370 8162 13375
rect 7966 13258 7994 13263
rect 7966 13211 7994 13230
rect 8078 13202 8106 13207
rect 7686 13119 7687 13145
rect 7713 13119 7714 13145
rect 6286 13043 6314 13062
rect 7350 13089 7378 13095
rect 7350 13063 7351 13089
rect 7377 13063 7378 13089
rect 2238 12950 2370 12955
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2238 12917 2370 12922
rect 7350 12866 7378 13063
rect 7350 12833 7378 12838
rect 7686 12809 7714 13119
rect 8022 13201 8106 13202
rect 8022 13175 8079 13201
rect 8105 13175 8106 13201
rect 8022 13174 8106 13175
rect 7686 12783 7687 12809
rect 7713 12783 7714 12809
rect 7686 12777 7714 12783
rect 7854 13090 7882 13095
rect 7854 12809 7882 13062
rect 7854 12783 7855 12809
rect 7881 12783 7882 12809
rect 7854 12777 7882 12783
rect 7910 12754 7938 12759
rect 7910 12707 7938 12726
rect 8022 12418 8050 13174
rect 8078 13169 8106 13174
rect 8134 13201 8162 13342
rect 8246 13257 8274 13454
rect 8246 13231 8247 13257
rect 8273 13231 8274 13257
rect 8246 13225 8274 13231
rect 8750 13257 8778 13566
rect 9086 13561 9114 13566
rect 9254 13874 9282 15946
rect 9918 15694 10050 15699
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 9918 15661 10050 15666
rect 9918 14910 10050 14915
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 9918 14877 10050 14882
rect 9198 13482 9226 13487
rect 9254 13482 9282 13846
rect 9590 14713 9618 14719
rect 9590 14687 9591 14713
rect 9617 14687 9618 14713
rect 9590 14266 9618 14687
rect 9590 13929 9618 14238
rect 9982 14657 10010 14663
rect 9982 14631 9983 14657
rect 10009 14631 10010 14657
rect 9982 14210 10010 14631
rect 10710 14658 10738 18999
rect 10766 18746 10794 20600
rect 11102 19138 11130 20600
rect 11214 19138 11242 19143
rect 11102 19137 11242 19138
rect 11102 19111 11215 19137
rect 11241 19111 11242 19137
rect 11102 19110 11242 19111
rect 11214 19105 11242 19110
rect 12446 19138 12474 20600
rect 17598 19222 17730 19227
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17598 19189 17730 19194
rect 12446 19105 12474 19110
rect 13062 19138 13090 19143
rect 13062 19091 13090 19110
rect 12670 19025 12698 19031
rect 12670 18999 12671 19025
rect 12697 18999 12698 19025
rect 10766 18713 10794 18718
rect 11382 18746 11410 18751
rect 11382 18699 11410 18718
rect 10990 18633 11018 18639
rect 10990 18607 10991 18633
rect 11017 18607 11018 18633
rect 10738 14630 10794 14658
rect 10710 14625 10738 14630
rect 9982 14182 10178 14210
rect 9918 14126 10050 14131
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 9918 14093 10050 14098
rect 9590 13903 9591 13929
rect 9617 13903 9618 13929
rect 9590 13593 9618 13903
rect 9926 13874 9954 13879
rect 9590 13567 9591 13593
rect 9617 13567 9618 13593
rect 9590 13561 9618 13567
rect 9814 13873 9954 13874
rect 9814 13847 9927 13873
rect 9953 13847 9954 13873
rect 9814 13846 9954 13847
rect 9310 13482 9338 13487
rect 9254 13481 9338 13482
rect 9254 13455 9311 13481
rect 9337 13455 9338 13481
rect 9254 13454 9338 13455
rect 9198 13435 9226 13454
rect 9310 13449 9338 13454
rect 9366 13482 9394 13487
rect 9366 13435 9394 13454
rect 8750 13231 8751 13257
rect 8777 13231 8778 13257
rect 8750 13225 8778 13231
rect 8806 13426 8834 13431
rect 8134 13175 8135 13201
rect 8161 13175 8162 13201
rect 8134 13169 8162 13175
rect 8358 13201 8386 13207
rect 8358 13175 8359 13201
rect 8385 13175 8386 13201
rect 8246 12866 8274 12871
rect 8358 12866 8386 13175
rect 8414 13146 8442 13151
rect 8638 13146 8666 13151
rect 8414 13145 8666 13146
rect 8414 13119 8415 13145
rect 8441 13119 8639 13145
rect 8665 13119 8666 13145
rect 8414 13118 8666 13119
rect 8414 13113 8442 13118
rect 8638 13113 8666 13118
rect 8806 13145 8834 13398
rect 8806 13119 8807 13145
rect 8833 13119 8834 13145
rect 8358 12838 8442 12866
rect 8246 12809 8274 12838
rect 8246 12783 8247 12809
rect 8273 12783 8274 12809
rect 8246 12777 8274 12783
rect 8190 12754 8218 12759
rect 8190 12707 8218 12726
rect 8358 12753 8386 12759
rect 8358 12727 8359 12753
rect 8385 12727 8386 12753
rect 8246 12698 8274 12703
rect 8134 12642 8162 12647
rect 8246 12642 8274 12670
rect 8134 12641 8274 12642
rect 8134 12615 8135 12641
rect 8161 12615 8274 12641
rect 8134 12614 8274 12615
rect 8302 12641 8330 12647
rect 8302 12615 8303 12641
rect 8329 12615 8330 12641
rect 8134 12609 8162 12614
rect 8022 12390 8218 12418
rect 8190 12362 8218 12390
rect 8190 12361 8274 12362
rect 8190 12335 8191 12361
rect 8217 12335 8274 12361
rect 8190 12334 8274 12335
rect 8190 12329 8218 12334
rect 8078 12306 8106 12311
rect 7910 12278 8078 12306
rect 2238 12166 2370 12171
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2238 12133 2370 12138
rect 6734 12025 6762 12031
rect 6734 11999 6735 12025
rect 6761 11999 6762 12025
rect 2142 11970 2170 11975
rect 2142 11923 2170 11942
rect 6734 11970 6762 11999
rect 6734 11937 6762 11942
rect 7798 11914 7826 11919
rect 7798 11867 7826 11886
rect 5894 11634 5922 11639
rect 5894 11587 5922 11606
rect 5558 11577 5586 11583
rect 5558 11551 5559 11577
rect 5585 11551 5586 11577
rect 2238 11382 2370 11387
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2238 11349 2370 11354
rect 5558 10962 5586 11551
rect 7182 11578 7210 11583
rect 7182 11531 7210 11550
rect 7406 11578 7434 11583
rect 7434 11550 7490 11578
rect 7406 11545 7434 11550
rect 6958 11522 6986 11527
rect 6958 11475 6986 11494
rect 5558 10929 5586 10934
rect 5838 10962 5866 10967
rect 2086 10761 2114 10766
rect 5838 10793 5866 10934
rect 7462 10962 7490 11550
rect 5838 10767 5839 10793
rect 5865 10767 5866 10793
rect 5838 10761 5866 10767
rect 7238 10906 7266 10911
rect 6174 10738 6202 10743
rect 6174 10691 6202 10710
rect 6846 10738 6874 10743
rect 2238 10598 2370 10603
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2238 10565 2370 10570
rect 6846 10345 6874 10710
rect 7238 10737 7266 10878
rect 7406 10738 7434 10743
rect 7238 10711 7239 10737
rect 7265 10711 7266 10737
rect 7238 10705 7266 10711
rect 7294 10737 7434 10738
rect 7294 10711 7407 10737
rect 7433 10711 7434 10737
rect 7294 10710 7434 10711
rect 7294 10514 7322 10710
rect 7406 10705 7434 10710
rect 7014 10486 7322 10514
rect 7014 10401 7042 10486
rect 7406 10458 7434 10463
rect 7462 10458 7490 10934
rect 7518 11522 7546 11527
rect 7518 10906 7546 11494
rect 7742 11185 7770 11191
rect 7742 11159 7743 11185
rect 7769 11159 7770 11185
rect 7742 10906 7770 11159
rect 7518 10878 7714 10906
rect 7686 10850 7714 10878
rect 7742 10873 7770 10878
rect 7854 11186 7882 11191
rect 7854 11129 7882 11158
rect 7854 11103 7855 11129
rect 7881 11103 7882 11129
rect 7686 10793 7714 10822
rect 7686 10767 7687 10793
rect 7713 10767 7714 10793
rect 7686 10761 7714 10767
rect 7854 10793 7882 11103
rect 7854 10767 7855 10793
rect 7881 10767 7882 10793
rect 7854 10761 7882 10767
rect 7406 10457 7490 10458
rect 7406 10431 7407 10457
rect 7433 10431 7490 10457
rect 7406 10430 7490 10431
rect 7406 10425 7434 10430
rect 7014 10375 7015 10401
rect 7041 10375 7042 10401
rect 7014 10369 7042 10375
rect 6846 10319 6847 10345
rect 6873 10319 6874 10345
rect 6846 10094 6874 10319
rect 6846 10066 6986 10094
rect 2142 10010 2170 10015
rect 2142 9963 2170 9982
rect 4998 10010 5026 10015
rect 966 9898 994 9903
rect 966 9851 994 9870
rect 2238 9814 2370 9819
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2238 9781 2370 9786
rect 4998 9673 5026 9982
rect 4998 9647 4999 9673
rect 5025 9647 5026 9673
rect 4998 9562 5026 9647
rect 6062 9954 6090 9959
rect 6062 9673 6090 9926
rect 6062 9647 6063 9673
rect 6089 9647 6090 9673
rect 6062 9641 6090 9647
rect 6454 9618 6482 9623
rect 6454 9571 6482 9590
rect 6790 9618 6818 9623
rect 4998 9529 5026 9534
rect 6790 9505 6818 9590
rect 6958 9562 6986 10066
rect 7126 10066 7154 10071
rect 7070 10010 7098 10015
rect 7070 9963 7098 9982
rect 7014 9954 7042 9959
rect 7014 9907 7042 9926
rect 7070 9618 7098 9623
rect 7126 9618 7154 10038
rect 7630 10065 7658 10071
rect 7630 10039 7631 10065
rect 7657 10039 7658 10065
rect 7182 10009 7210 10015
rect 7182 9983 7183 10009
rect 7209 9983 7210 10009
rect 7182 9898 7210 9983
rect 7182 9865 7210 9870
rect 7238 10010 7266 10015
rect 7070 9617 7154 9618
rect 7070 9591 7071 9617
rect 7097 9591 7154 9617
rect 7070 9590 7154 9591
rect 7070 9585 7098 9590
rect 7014 9562 7042 9567
rect 6958 9561 7042 9562
rect 6958 9535 7015 9561
rect 7041 9535 7042 9561
rect 6958 9534 7042 9535
rect 6790 9479 6791 9505
rect 6817 9479 6818 9505
rect 6510 9338 6538 9343
rect 6510 9225 6538 9310
rect 6510 9199 6511 9225
rect 6537 9199 6538 9225
rect 6510 9193 6538 9199
rect 6790 9226 6818 9479
rect 6902 9506 6930 9511
rect 6902 9505 6986 9506
rect 6902 9479 6903 9505
rect 6929 9479 6986 9505
rect 6902 9478 6986 9479
rect 6902 9473 6930 9478
rect 6902 9226 6930 9231
rect 6790 9225 6930 9226
rect 6790 9199 6903 9225
rect 6929 9199 6930 9225
rect 6790 9198 6930 9199
rect 5446 9170 5474 9175
rect 5390 9169 5474 9170
rect 5390 9143 5447 9169
rect 5473 9143 5474 9169
rect 5390 9142 5474 9143
rect 2238 9030 2370 9035
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2238 8997 2370 9002
rect 966 8890 994 8895
rect 966 8843 994 8862
rect 2142 8834 2170 8839
rect 2142 8787 2170 8806
rect 5390 8778 5418 9142
rect 5446 9137 5474 9142
rect 6902 9170 6930 9198
rect 6902 9137 6930 9142
rect 6790 8946 6818 8965
rect 6790 8913 6818 8918
rect 966 8442 994 8447
rect 966 8385 994 8414
rect 2142 8442 2170 8447
rect 2142 8395 2170 8414
rect 5390 8442 5418 8750
rect 5390 8409 5418 8414
rect 5446 8834 5474 8839
rect 966 8359 967 8385
rect 993 8359 994 8385
rect 966 8353 994 8359
rect 5446 8385 5474 8806
rect 6734 8834 6762 8839
rect 6846 8834 6874 8839
rect 6762 8806 6818 8834
rect 6734 8801 6762 8806
rect 6790 8777 6818 8806
rect 6958 8834 6986 9478
rect 7014 9225 7042 9534
rect 7238 9450 7266 9982
rect 7294 10009 7322 10015
rect 7294 9983 7295 10009
rect 7321 9983 7322 10009
rect 7294 9729 7322 9983
rect 7406 10010 7434 10015
rect 7518 10010 7546 10015
rect 7406 10009 7546 10010
rect 7406 9983 7407 10009
rect 7433 9983 7519 10009
rect 7545 9983 7546 10009
rect 7406 9982 7546 9983
rect 7406 9977 7434 9982
rect 7518 9977 7546 9982
rect 7294 9703 7295 9729
rect 7321 9703 7322 9729
rect 7294 9697 7322 9703
rect 7294 9562 7322 9567
rect 7294 9515 7322 9534
rect 7350 9562 7378 9567
rect 7350 9561 7434 9562
rect 7350 9535 7351 9561
rect 7377 9535 7434 9561
rect 7350 9534 7434 9535
rect 7350 9529 7378 9534
rect 7238 9422 7378 9450
rect 7238 9338 7266 9343
rect 7238 9291 7266 9310
rect 7294 9282 7322 9287
rect 7014 9199 7015 9225
rect 7041 9199 7042 9225
rect 7014 9193 7042 9199
rect 7238 9226 7266 9231
rect 7238 9179 7266 9198
rect 7294 9225 7322 9254
rect 7294 9199 7295 9225
rect 7321 9199 7322 9225
rect 7294 9193 7322 9199
rect 7126 8946 7154 8951
rect 7014 8834 7042 8839
rect 6958 8833 7042 8834
rect 6958 8807 7015 8833
rect 7041 8807 7042 8833
rect 6958 8806 7042 8807
rect 6846 8787 6874 8806
rect 7014 8801 7042 8806
rect 7126 8833 7154 8918
rect 7126 8807 7127 8833
rect 7153 8807 7154 8833
rect 7126 8801 7154 8807
rect 7238 8890 7266 8895
rect 7238 8833 7266 8862
rect 7238 8807 7239 8833
rect 7265 8807 7266 8833
rect 7238 8801 7266 8807
rect 7350 8833 7378 9422
rect 7350 8807 7351 8833
rect 7377 8807 7378 8833
rect 7350 8801 7378 8807
rect 7406 9169 7434 9534
rect 7406 9143 7407 9169
rect 7433 9143 7434 9169
rect 7406 9058 7434 9143
rect 7406 8834 7434 9030
rect 7518 9225 7546 9231
rect 7518 9199 7519 9225
rect 7545 9199 7546 9225
rect 7518 8945 7546 9199
rect 7630 9114 7658 10039
rect 7686 10066 7714 10071
rect 7686 10009 7714 10038
rect 7686 9983 7687 10009
rect 7713 9983 7714 10009
rect 7686 9954 7714 9983
rect 7686 9921 7714 9926
rect 7910 9953 7938 12278
rect 8078 12259 8106 12278
rect 8078 11970 8106 11975
rect 8078 11689 8106 11942
rect 8190 11969 8218 11975
rect 8190 11943 8191 11969
rect 8217 11943 8218 11969
rect 8078 11663 8079 11689
rect 8105 11663 8106 11689
rect 8078 11657 8106 11663
rect 8134 11858 8162 11863
rect 8022 11578 8050 11583
rect 7910 9927 7911 9953
rect 7937 9927 7938 9953
rect 7910 9898 7938 9927
rect 7910 9865 7938 9870
rect 7966 11577 8050 11578
rect 7966 11551 8023 11577
rect 8049 11551 8050 11577
rect 7966 11550 8050 11551
rect 7966 10010 7994 11550
rect 8022 11545 8050 11550
rect 8078 11466 8106 11471
rect 8134 11466 8162 11830
rect 8190 11578 8218 11943
rect 8246 11746 8274 12334
rect 8302 12026 8330 12615
rect 8358 12473 8386 12727
rect 8358 12447 8359 12473
rect 8385 12447 8386 12473
rect 8358 12441 8386 12447
rect 8414 12138 8442 12838
rect 8806 12698 8834 13119
rect 8806 12665 8834 12670
rect 9142 13146 9170 13151
rect 8806 12306 8834 12311
rect 8806 12259 8834 12278
rect 8414 12105 8442 12110
rect 9030 12138 9058 12143
rect 8862 12082 8890 12087
rect 8862 12035 8890 12054
rect 8302 11998 8554 12026
rect 8470 11914 8498 11919
rect 8470 11867 8498 11886
rect 8414 11858 8442 11863
rect 8414 11811 8442 11830
rect 8526 11858 8554 11998
rect 8526 11811 8554 11830
rect 8582 11969 8610 11975
rect 8582 11943 8583 11969
rect 8609 11943 8610 11969
rect 8246 11713 8274 11718
rect 8414 11634 8442 11639
rect 8190 11545 8218 11550
rect 8358 11578 8386 11583
rect 8358 11531 8386 11550
rect 8078 11465 8162 11466
rect 8078 11439 8079 11465
rect 8105 11439 8162 11465
rect 8078 11438 8162 11439
rect 8078 11433 8106 11438
rect 8246 11185 8274 11191
rect 8246 11159 8247 11185
rect 8273 11159 8274 11185
rect 8246 10906 8274 11159
rect 8414 10962 8442 11606
rect 8582 11634 8610 11943
rect 8582 11601 8610 11606
rect 8750 11969 8778 11975
rect 8750 11943 8751 11969
rect 8777 11943 8778 11969
rect 8750 11914 8778 11943
rect 8750 11298 8778 11886
rect 8918 11858 8946 11863
rect 8414 10929 8442 10934
rect 8470 11270 8778 11298
rect 8862 11746 8890 11751
rect 8470 11185 8498 11270
rect 8470 11159 8471 11185
rect 8497 11159 8498 11185
rect 8246 10873 8274 10878
rect 8302 10850 8330 10855
rect 8302 10793 8330 10822
rect 8302 10767 8303 10793
rect 8329 10767 8330 10793
rect 8302 10761 8330 10767
rect 8414 10849 8442 10855
rect 8414 10823 8415 10849
rect 8441 10823 8442 10849
rect 8414 10346 8442 10823
rect 8414 10121 8442 10318
rect 8414 10095 8415 10121
rect 8441 10095 8442 10121
rect 8414 10089 8442 10095
rect 7854 9562 7882 9567
rect 7966 9562 7994 9982
rect 8246 10065 8274 10071
rect 8246 10039 8247 10065
rect 8273 10039 8274 10065
rect 8246 9786 8274 10039
rect 8470 9786 8498 11159
rect 8806 11185 8834 11191
rect 8806 11159 8807 11185
rect 8833 11159 8834 11185
rect 8806 11018 8834 11159
rect 8694 10990 8834 11018
rect 8582 10962 8610 10967
rect 8610 10934 8666 10962
rect 8582 10929 8610 10934
rect 8638 10682 8666 10934
rect 8694 10850 8722 10990
rect 8694 10803 8722 10822
rect 8806 10906 8834 10911
rect 8806 10793 8834 10878
rect 8806 10767 8807 10793
rect 8833 10767 8834 10793
rect 8806 10761 8834 10767
rect 8638 10654 8834 10682
rect 8246 9758 8386 9786
rect 8022 9674 8050 9679
rect 8022 9617 8050 9646
rect 8022 9591 8023 9617
rect 8049 9591 8050 9617
rect 8022 9585 8050 9591
rect 8302 9674 8330 9679
rect 8302 9617 8330 9646
rect 8302 9591 8303 9617
rect 8329 9591 8330 9617
rect 8302 9585 8330 9591
rect 7798 9561 7994 9562
rect 7798 9535 7855 9561
rect 7881 9535 7994 9561
rect 7798 9534 7994 9535
rect 7630 9081 7658 9086
rect 7742 9170 7770 9175
rect 7518 8919 7519 8945
rect 7545 8919 7546 8945
rect 7518 8913 7546 8919
rect 7406 8801 7434 8806
rect 6790 8751 6791 8777
rect 6817 8751 6818 8777
rect 6790 8745 6818 8751
rect 7574 8778 7602 8783
rect 7574 8731 7602 8750
rect 6510 8722 6538 8727
rect 6510 8497 6538 8694
rect 7406 8722 7434 8727
rect 7406 8675 7434 8694
rect 6510 8471 6511 8497
rect 6537 8471 6538 8497
rect 6510 8465 6538 8471
rect 7126 8666 7154 8671
rect 5446 8359 5447 8385
rect 5473 8359 5474 8385
rect 5446 8353 5474 8359
rect 6902 8441 6930 8447
rect 6902 8415 6903 8441
rect 6929 8415 6930 8441
rect 6902 8386 6930 8415
rect 7126 8386 7154 8638
rect 7742 8666 7770 9142
rect 7742 8633 7770 8638
rect 7742 8554 7770 8559
rect 7798 8554 7826 9534
rect 7854 9529 7882 9534
rect 8134 9505 8162 9511
rect 8134 9479 8135 9505
rect 8161 9479 8162 9505
rect 8134 9282 8162 9479
rect 8246 9505 8274 9511
rect 8246 9479 8247 9505
rect 8273 9479 8274 9505
rect 8246 9450 8274 9479
rect 8246 9417 8274 9422
rect 8134 9249 8162 9254
rect 7742 8553 7826 8554
rect 7742 8527 7743 8553
rect 7769 8527 7826 8553
rect 7742 8526 7826 8527
rect 7854 9114 7882 9119
rect 7854 8553 7882 9086
rect 8358 9114 8386 9758
rect 8470 9753 8498 9758
rect 8694 9674 8722 9679
rect 8694 9627 8722 9646
rect 8582 9618 8610 9623
rect 8582 9571 8610 9590
rect 8750 9505 8778 9511
rect 8750 9479 8751 9505
rect 8777 9479 8778 9505
rect 8750 9338 8778 9479
rect 8750 9305 8778 9310
rect 8806 9337 8834 10654
rect 8862 10457 8890 11718
rect 8918 11466 8946 11830
rect 8974 11634 9002 11639
rect 8974 11587 9002 11606
rect 9030 11634 9058 12110
rect 9142 12025 9170 13118
rect 9814 13034 9842 13846
rect 9926 13841 9954 13846
rect 10150 13537 10178 14182
rect 10710 13650 10738 13655
rect 10150 13511 10151 13537
rect 10177 13511 10178 13537
rect 10150 13505 10178 13511
rect 10318 13649 10738 13650
rect 10318 13623 10711 13649
rect 10737 13623 10738 13649
rect 10318 13622 10738 13623
rect 10318 13537 10346 13622
rect 10710 13617 10738 13622
rect 10318 13511 10319 13537
rect 10345 13511 10346 13537
rect 10318 13505 10346 13511
rect 10654 13482 10682 13487
rect 10654 13435 10682 13454
rect 10710 13482 10738 13487
rect 10766 13482 10794 14630
rect 10710 13481 10794 13482
rect 10710 13455 10711 13481
rect 10737 13455 10794 13481
rect 10710 13454 10794 13455
rect 10934 14266 10962 14271
rect 10710 13449 10738 13454
rect 10262 13425 10290 13431
rect 10262 13399 10263 13425
rect 10289 13399 10290 13425
rect 9918 13342 10050 13347
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 9918 13309 10050 13314
rect 9926 13202 9954 13207
rect 9926 13155 9954 13174
rect 9870 13146 9898 13151
rect 9870 13099 9898 13118
rect 9926 13034 9954 13039
rect 9814 13033 9954 13034
rect 9814 13007 9927 13033
rect 9953 13007 9954 13033
rect 9814 13006 9954 13007
rect 9926 13001 9954 13006
rect 10206 12698 10234 12703
rect 10206 12651 10234 12670
rect 9918 12558 10050 12563
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 9918 12525 10050 12530
rect 9814 12361 9842 12367
rect 9814 12335 9815 12361
rect 9841 12335 9842 12361
rect 9142 11999 9143 12025
rect 9169 11999 9170 12025
rect 9142 11993 9170 11999
rect 9478 12082 9506 12087
rect 9366 11969 9394 11975
rect 9366 11943 9367 11969
rect 9393 11943 9394 11969
rect 9142 11914 9170 11919
rect 9366 11914 9394 11943
rect 9422 11914 9450 11919
rect 9170 11886 9226 11914
rect 9142 11881 9170 11886
rect 9086 11857 9114 11863
rect 9086 11831 9087 11857
rect 9113 11831 9114 11857
rect 9086 11746 9114 11831
rect 9198 11857 9226 11886
rect 9198 11831 9199 11857
rect 9225 11831 9226 11857
rect 9198 11825 9226 11831
rect 9366 11886 9422 11914
rect 9086 11713 9114 11718
rect 9030 11633 9170 11634
rect 9030 11607 9031 11633
rect 9057 11607 9170 11633
rect 9030 11606 9170 11607
rect 9030 11601 9058 11606
rect 8974 11466 9002 11471
rect 8946 11465 9002 11466
rect 8946 11439 8975 11465
rect 9001 11439 9002 11465
rect 8946 11438 9002 11439
rect 8918 11433 8946 11438
rect 8974 11433 9002 11438
rect 8862 10431 8863 10457
rect 8889 10431 8890 10457
rect 8862 10425 8890 10431
rect 8918 11186 8946 11191
rect 8862 10346 8890 10365
rect 8862 9730 8890 10318
rect 8862 9697 8890 9702
rect 8918 10009 8946 11158
rect 9086 11074 9114 11079
rect 9086 11027 9114 11046
rect 9142 10962 9170 11606
rect 9254 11578 9282 11583
rect 9254 11531 9282 11550
rect 9086 10934 9170 10962
rect 8974 10682 9002 10687
rect 8974 10635 9002 10654
rect 8974 10290 9002 10295
rect 9086 10290 9114 10934
rect 9142 10402 9170 10407
rect 9310 10402 9338 10407
rect 9142 10401 9338 10402
rect 9142 10375 9143 10401
rect 9169 10375 9311 10401
rect 9337 10375 9338 10401
rect 9142 10374 9338 10375
rect 9142 10369 9170 10374
rect 8974 10289 9058 10290
rect 8974 10263 8975 10289
rect 9001 10263 9058 10289
rect 8974 10262 9058 10263
rect 9086 10262 9170 10290
rect 8974 10257 9002 10262
rect 9030 10234 9058 10262
rect 9030 10206 9114 10234
rect 8918 9983 8919 10009
rect 8945 9983 8946 10009
rect 8918 9618 8946 9983
rect 8918 9585 8946 9590
rect 9030 9954 9058 9959
rect 9086 9954 9114 10206
rect 9030 9953 9114 9954
rect 9030 9927 9031 9953
rect 9057 9927 9114 9953
rect 9030 9926 9114 9927
rect 9030 9618 9058 9926
rect 9142 9898 9170 10262
rect 9310 10122 9338 10374
rect 9310 10089 9338 10094
rect 9366 10346 9394 11886
rect 9422 11881 9450 11886
rect 9422 11634 9450 11639
rect 9422 11242 9450 11606
rect 9478 11297 9506 12054
rect 9646 11522 9674 11527
rect 9646 11475 9674 11494
rect 9478 11271 9479 11297
rect 9505 11271 9506 11297
rect 9478 11265 9506 11271
rect 9422 11185 9450 11214
rect 9422 11159 9423 11185
rect 9449 11159 9450 11185
rect 9422 11153 9450 11159
rect 9478 11073 9506 11079
rect 9478 11047 9479 11073
rect 9505 11047 9506 11073
rect 9478 10906 9506 11047
rect 9758 11074 9786 11079
rect 9758 11027 9786 11046
rect 9478 10873 9506 10878
rect 9478 10794 9506 10799
rect 9478 10747 9506 10766
rect 9702 10794 9730 10799
rect 9702 10747 9730 10766
rect 9702 10514 9730 10519
rect 9814 10514 9842 12335
rect 10150 11970 10178 11975
rect 10262 11970 10290 13399
rect 10654 13258 10682 13263
rect 10654 13211 10682 13230
rect 10542 13202 10570 13207
rect 10542 13155 10570 13174
rect 10710 13146 10738 13151
rect 10710 13099 10738 13118
rect 10934 13145 10962 14238
rect 10990 13873 11018 18607
rect 11046 14658 11074 14663
rect 11046 14611 11074 14630
rect 11326 14657 11354 14663
rect 11326 14631 11327 14657
rect 11353 14631 11354 14657
rect 11214 14266 11242 14271
rect 11326 14266 11354 14631
rect 11242 14238 11354 14266
rect 11214 14041 11242 14238
rect 11214 14015 11215 14041
rect 11241 14015 11242 14041
rect 11214 14009 11242 14015
rect 10990 13847 10991 13873
rect 11017 13847 11018 13873
rect 10990 13258 11018 13847
rect 10990 13225 11018 13230
rect 12334 13202 12362 13207
rect 10934 13119 10935 13145
rect 10961 13119 10962 13145
rect 10934 12754 10962 13119
rect 10878 12726 10934 12754
rect 10374 12642 10402 12647
rect 10766 12642 10794 12647
rect 10374 12641 10794 12642
rect 10374 12615 10375 12641
rect 10401 12615 10767 12641
rect 10793 12615 10794 12641
rect 10374 12614 10794 12615
rect 10374 12609 10402 12614
rect 10486 12305 10514 12311
rect 10486 12279 10487 12305
rect 10513 12279 10514 12305
rect 10486 12026 10514 12279
rect 10150 11969 10458 11970
rect 10150 11943 10151 11969
rect 10177 11943 10458 11969
rect 10150 11942 10458 11943
rect 10150 11937 10178 11942
rect 9982 11914 10010 11919
rect 9982 11867 10010 11886
rect 10038 11858 10066 11863
rect 10038 11857 10122 11858
rect 10038 11831 10039 11857
rect 10065 11831 10122 11857
rect 10038 11830 10122 11831
rect 10038 11825 10066 11830
rect 9918 11774 10050 11779
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 9918 11741 10050 11746
rect 10094 11690 10122 11830
rect 9926 11662 10122 11690
rect 9926 11186 9954 11662
rect 10430 11466 10458 11942
rect 10486 11578 10514 11998
rect 10486 11545 10514 11550
rect 10710 11521 10738 11527
rect 10710 11495 10711 11521
rect 10737 11495 10738 11521
rect 10430 11438 10626 11466
rect 9926 11129 9954 11158
rect 10318 11242 10346 11247
rect 9926 11103 9927 11129
rect 9953 11103 9954 11129
rect 9926 11097 9954 11103
rect 10150 11130 10178 11135
rect 10150 11083 10178 11102
rect 10318 11129 10346 11214
rect 10598 11185 10626 11438
rect 10598 11159 10599 11185
rect 10625 11159 10626 11185
rect 10598 11153 10626 11159
rect 10318 11103 10319 11129
rect 10345 11103 10346 11129
rect 10318 11097 10346 11103
rect 10094 11074 10122 11079
rect 10094 11027 10122 11046
rect 10206 11073 10234 11079
rect 10206 11047 10207 11073
rect 10233 11047 10234 11073
rect 9918 10990 10050 10995
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 9918 10957 10050 10962
rect 9730 10486 9842 10514
rect 9926 10906 9954 10911
rect 9422 10346 9450 10351
rect 9366 10345 9450 10346
rect 9366 10319 9423 10345
rect 9449 10319 9450 10345
rect 9366 10318 9450 10319
rect 9366 9954 9394 10318
rect 9422 10313 9450 10318
rect 9366 9921 9394 9926
rect 9478 10009 9506 10015
rect 9478 9983 9479 10009
rect 9505 9983 9506 10009
rect 9030 9585 9058 9590
rect 9086 9870 9170 9898
rect 8862 9562 8890 9567
rect 8862 9515 8890 9534
rect 8806 9311 8807 9337
rect 8833 9311 8834 9337
rect 8806 9226 8834 9311
rect 9030 9506 9058 9511
rect 8358 9081 8386 9086
rect 8694 9198 8834 9226
rect 8862 9226 8890 9231
rect 8414 8890 8442 8895
rect 8414 8843 8442 8862
rect 8694 8833 8722 9198
rect 8862 8889 8890 9198
rect 8974 9226 9002 9231
rect 8974 9179 9002 9198
rect 8974 8946 9002 8951
rect 9030 8946 9058 9478
rect 9086 9505 9114 9870
rect 9086 9479 9087 9505
rect 9113 9479 9114 9505
rect 9086 9450 9114 9479
rect 9086 9417 9114 9422
rect 9142 9786 9170 9791
rect 9142 9337 9170 9758
rect 9310 9562 9338 9581
rect 9478 9562 9506 9983
rect 9310 9529 9338 9534
rect 9366 9561 9618 9562
rect 9366 9535 9479 9561
rect 9505 9535 9618 9561
rect 9366 9534 9618 9535
rect 9142 9311 9143 9337
rect 9169 9311 9170 9337
rect 9142 9305 9170 9311
rect 9254 9338 9282 9343
rect 9366 9338 9394 9534
rect 9478 9529 9506 9534
rect 9254 9337 9394 9338
rect 9254 9311 9255 9337
rect 9281 9311 9394 9337
rect 9254 9310 9394 9311
rect 9254 9226 9282 9310
rect 9478 9282 9506 9287
rect 9422 9226 9450 9231
rect 9254 9193 9282 9198
rect 9310 9225 9450 9226
rect 9310 9199 9423 9225
rect 9449 9199 9450 9225
rect 9310 9198 9450 9199
rect 9198 9170 9226 9175
rect 9198 9123 9226 9142
rect 8974 8945 9058 8946
rect 8974 8919 8975 8945
rect 9001 8919 9058 8945
rect 8974 8918 9058 8919
rect 8974 8913 9002 8918
rect 8862 8863 8863 8889
rect 8889 8863 8890 8889
rect 8862 8857 8890 8863
rect 9030 8890 9058 8918
rect 9030 8857 9058 8862
rect 9198 8890 9226 8895
rect 8806 8834 8834 8839
rect 8694 8807 8695 8833
rect 8721 8807 8722 8833
rect 8694 8801 8722 8807
rect 8750 8806 8806 8834
rect 7854 8527 7855 8553
rect 7881 8527 7882 8553
rect 7742 8521 7770 8526
rect 7854 8521 7882 8527
rect 8414 8721 8442 8727
rect 8414 8695 8415 8721
rect 8441 8695 8442 8721
rect 8414 8554 8442 8695
rect 8526 8722 8554 8727
rect 8526 8675 8554 8694
rect 8442 8526 8554 8554
rect 8414 8521 8442 8526
rect 8078 8441 8106 8447
rect 8078 8415 8079 8441
rect 8105 8415 8106 8441
rect 6902 8385 7154 8386
rect 6902 8359 7127 8385
rect 7153 8359 7154 8385
rect 6902 8358 7154 8359
rect 2238 8246 2370 8251
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2238 8213 2370 8218
rect 7014 7657 7042 7663
rect 7014 7631 7015 7657
rect 7041 7631 7042 7657
rect 7014 7602 7042 7631
rect 7070 7602 7098 7607
rect 7126 7602 7154 8358
rect 7350 8386 7378 8391
rect 7350 7713 7378 8358
rect 7798 8386 7826 8391
rect 7798 8339 7826 8358
rect 8078 8162 8106 8415
rect 8078 8129 8106 8134
rect 8414 8162 8442 8167
rect 8414 8105 8442 8134
rect 8414 8079 8415 8105
rect 8441 8079 8442 8105
rect 8414 8073 8442 8079
rect 8526 8049 8554 8526
rect 8526 8023 8527 8049
rect 8553 8023 8554 8049
rect 7350 7687 7351 7713
rect 7377 7687 7378 7713
rect 7350 7681 7378 7687
rect 8414 7937 8442 7943
rect 8414 7911 8415 7937
rect 8441 7911 8442 7937
rect 7014 7574 7070 7602
rect 7098 7574 7154 7602
rect 8414 7601 8442 7911
rect 8414 7575 8415 7601
rect 8441 7575 8442 7601
rect 7070 7569 7098 7574
rect 2238 7462 2370 7467
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2238 7429 2370 7434
rect 8134 7154 8162 7159
rect 2238 6678 2370 6683
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2238 6645 2370 6650
rect 8134 6537 8162 7126
rect 8134 6511 8135 6537
rect 8161 6511 8162 6537
rect 8134 6505 8162 6511
rect 7798 6482 7826 6487
rect 7798 6435 7826 6454
rect 2238 5894 2370 5899
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2238 5861 2370 5866
rect 2238 5110 2370 5115
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2238 5077 2370 5082
rect 2238 4326 2370 4331
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2238 4293 2370 4298
rect 8414 4214 8442 7575
rect 8526 7574 8554 8023
rect 8694 8050 8722 8055
rect 8750 8050 8778 8806
rect 8806 8787 8834 8806
rect 9086 8610 9114 8615
rect 9086 8554 9114 8582
rect 9030 8553 9114 8554
rect 9030 8527 9087 8553
rect 9113 8527 9114 8553
rect 9030 8526 9114 8527
rect 8862 8442 8890 8447
rect 8862 8395 8890 8414
rect 8974 8386 9002 8391
rect 8974 8339 9002 8358
rect 8694 8049 8778 8050
rect 8694 8023 8695 8049
rect 8721 8023 8778 8049
rect 8694 8022 8778 8023
rect 8694 8017 8722 8022
rect 8862 7937 8890 7943
rect 8862 7911 8863 7937
rect 8889 7911 8890 7937
rect 8750 7658 8778 7663
rect 8862 7658 8890 7911
rect 8750 7657 8890 7658
rect 8750 7631 8751 7657
rect 8777 7631 8890 7657
rect 8750 7630 8890 7631
rect 8750 7602 8778 7630
rect 8526 7546 8722 7574
rect 8750 7569 8778 7574
rect 8694 7490 8722 7546
rect 8694 7462 8946 7490
rect 8638 7322 8666 7327
rect 8862 7322 8890 7327
rect 8638 7321 8890 7322
rect 8638 7295 8639 7321
rect 8665 7295 8863 7321
rect 8889 7295 8890 7321
rect 8638 7294 8890 7295
rect 8638 7289 8666 7294
rect 8862 7289 8890 7294
rect 8918 7265 8946 7462
rect 8918 7239 8919 7265
rect 8945 7239 8946 7265
rect 8918 7233 8946 7239
rect 9030 7265 9058 8526
rect 9086 8521 9114 8526
rect 9198 8553 9226 8862
rect 9254 8834 9282 8839
rect 9310 8834 9338 9198
rect 9422 9193 9450 9198
rect 9366 9058 9394 9063
rect 9366 8889 9394 9030
rect 9366 8863 9367 8889
rect 9393 8863 9394 8889
rect 9366 8857 9394 8863
rect 9254 8833 9338 8834
rect 9254 8807 9255 8833
rect 9281 8807 9338 8833
rect 9254 8806 9338 8807
rect 9254 8801 9282 8806
rect 9310 8778 9338 8806
rect 9310 8745 9338 8750
rect 9478 8777 9506 9254
rect 9590 9281 9618 9534
rect 9590 9255 9591 9281
rect 9617 9255 9618 9281
rect 9590 9249 9618 9255
rect 9702 9170 9730 10486
rect 9926 10402 9954 10878
rect 9926 10355 9954 10374
rect 10206 10458 10234 11047
rect 10094 10289 10122 10295
rect 10094 10263 10095 10289
rect 10121 10263 10122 10289
rect 9918 10206 10050 10211
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 9918 10173 10050 10178
rect 9814 10065 9842 10071
rect 9814 10039 9815 10065
rect 9841 10039 9842 10065
rect 9814 9786 9842 10039
rect 9814 9753 9842 9758
rect 9870 10066 9898 10071
rect 9758 9730 9786 9735
rect 9758 9281 9786 9702
rect 9814 9506 9842 9511
rect 9814 9459 9842 9478
rect 9870 9505 9898 10038
rect 10094 10010 10122 10263
rect 10206 10066 10234 10430
rect 10710 10402 10738 11495
rect 10710 10369 10738 10374
rect 10262 10066 10290 10071
rect 10206 10038 10262 10066
rect 10262 10019 10290 10038
rect 10710 10010 10738 10015
rect 10094 9977 10122 9982
rect 10654 9982 10710 10010
rect 10654 9729 10682 9982
rect 10710 9977 10738 9982
rect 10654 9703 10655 9729
rect 10681 9703 10682 9729
rect 9870 9479 9871 9505
rect 9897 9479 9898 9505
rect 9870 9473 9898 9479
rect 10038 9562 10066 9567
rect 10038 9506 10066 9534
rect 10038 9478 10122 9506
rect 9918 9422 10050 9427
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 9918 9389 10050 9394
rect 9758 9255 9759 9281
rect 9785 9255 9786 9281
rect 9758 9249 9786 9255
rect 9926 9282 9954 9287
rect 9926 9235 9954 9254
rect 9478 8751 9479 8777
rect 9505 8751 9506 8777
rect 9198 8527 9199 8553
rect 9225 8527 9226 8553
rect 9198 8521 9226 8527
rect 9254 8722 9282 8727
rect 9254 8442 9282 8694
rect 9142 8385 9170 8391
rect 9142 8359 9143 8385
rect 9169 8359 9170 8385
rect 9086 7714 9114 7719
rect 9142 7714 9170 8359
rect 9086 7713 9170 7714
rect 9086 7687 9087 7713
rect 9113 7687 9170 7713
rect 9086 7686 9170 7687
rect 9086 7681 9114 7686
rect 9030 7239 9031 7265
rect 9057 7239 9058 7265
rect 9030 7233 9058 7239
rect 9254 7265 9282 8414
rect 9422 8386 9450 8391
rect 9422 8161 9450 8358
rect 9478 8274 9506 8751
rect 9590 9142 9730 9170
rect 10094 9225 10122 9478
rect 10654 9394 10682 9703
rect 10766 9673 10794 12614
rect 10822 12026 10850 12031
rect 10878 12026 10906 12726
rect 10934 12721 10962 12726
rect 10990 13146 11018 13151
rect 10934 12642 10962 12647
rect 10990 12642 11018 13118
rect 11270 13090 11298 13095
rect 11270 13043 11298 13062
rect 11774 13090 11802 13095
rect 11774 12809 11802 13062
rect 12334 13089 12362 13174
rect 12670 13202 12698 18999
rect 17598 18438 17730 18443
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17598 18405 17730 18410
rect 17598 17654 17730 17659
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17598 17621 17730 17626
rect 17598 16870 17730 16875
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17598 16837 17730 16842
rect 17598 16086 17730 16091
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17598 16053 17730 16058
rect 17598 15302 17730 15307
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17598 15269 17730 15274
rect 17598 14518 17730 14523
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17598 14485 17730 14490
rect 17598 13734 17730 13739
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17598 13701 17730 13706
rect 20006 13593 20034 13599
rect 20006 13567 20007 13593
rect 20033 13567 20034 13593
rect 18942 13537 18970 13543
rect 18942 13511 18943 13537
rect 18969 13511 18970 13537
rect 12670 13155 12698 13174
rect 13566 13202 13594 13207
rect 13566 13201 13650 13202
rect 13566 13175 13567 13201
rect 13593 13175 13650 13201
rect 13566 13174 13650 13175
rect 13566 13169 13594 13174
rect 12726 13146 12754 13151
rect 12726 13099 12754 13118
rect 13510 13146 13538 13151
rect 12334 13063 12335 13089
rect 12361 13063 12362 13089
rect 12334 13057 12362 13063
rect 12950 13089 12978 13095
rect 12950 13063 12951 13089
rect 12977 13063 12978 13089
rect 11774 12783 11775 12809
rect 11801 12783 11802 12809
rect 11774 12777 11802 12783
rect 12054 13034 12082 13039
rect 12054 12753 12082 13006
rect 12670 13034 12698 13039
rect 12670 12987 12698 13006
rect 12054 12727 12055 12753
rect 12081 12727 12082 12753
rect 12054 12721 12082 12727
rect 12446 12754 12474 12759
rect 12446 12707 12474 12726
rect 12670 12754 12698 12759
rect 10934 12641 11018 12642
rect 10934 12615 10935 12641
rect 10961 12615 11018 12641
rect 10934 12614 11018 12615
rect 11718 12641 11746 12647
rect 11718 12615 11719 12641
rect 11745 12615 11746 12641
rect 10934 12609 10962 12614
rect 10850 11998 10962 12026
rect 10822 11979 10850 11998
rect 10934 11577 10962 11998
rect 11718 11802 11746 12615
rect 11830 12641 11858 12647
rect 11830 12615 11831 12641
rect 11857 12615 11858 12641
rect 11830 12082 11858 12615
rect 11830 12049 11858 12054
rect 12670 11802 12698 12726
rect 12950 12754 12978 13063
rect 12950 12721 12978 12726
rect 13174 13034 13202 13039
rect 13006 12697 13034 12703
rect 13006 12671 13007 12697
rect 13033 12671 13034 12697
rect 12894 12474 12922 12479
rect 13006 12474 13034 12671
rect 12894 12473 13034 12474
rect 12894 12447 12895 12473
rect 12921 12447 13034 12473
rect 12894 12446 13034 12447
rect 12894 12441 12922 12446
rect 12838 12362 12866 12367
rect 11718 11774 11802 11802
rect 10934 11551 10935 11577
rect 10961 11551 10962 11577
rect 10934 11545 10962 11551
rect 10878 11522 10906 11527
rect 10878 11241 10906 11494
rect 11270 11522 11298 11527
rect 11270 11521 11522 11522
rect 11270 11495 11271 11521
rect 11297 11495 11522 11521
rect 11270 11494 11522 11495
rect 11270 11489 11298 11494
rect 10878 11215 10879 11241
rect 10905 11215 10906 11241
rect 10878 11209 10906 11215
rect 11214 11242 11242 11247
rect 10934 11186 10962 11191
rect 11102 11186 11130 11191
rect 10962 11185 11130 11186
rect 10962 11159 11103 11185
rect 11129 11159 11130 11185
rect 10962 11158 11130 11159
rect 10934 11139 10962 11158
rect 11102 11153 11130 11158
rect 11214 11129 11242 11214
rect 11494 11241 11522 11494
rect 11494 11215 11495 11241
rect 11521 11215 11522 11241
rect 11494 11209 11522 11215
rect 11438 11186 11466 11191
rect 11438 11139 11466 11158
rect 11606 11186 11634 11191
rect 11606 11139 11634 11158
rect 11214 11103 11215 11129
rect 11241 11103 11242 11129
rect 11214 11097 11242 11103
rect 11718 11129 11746 11135
rect 11718 11103 11719 11129
rect 11745 11103 11746 11129
rect 10822 11073 10850 11079
rect 10822 11047 10823 11073
rect 10849 11047 10850 11073
rect 10822 10066 10850 11047
rect 11158 11073 11186 11079
rect 11158 11047 11159 11073
rect 11185 11047 11186 11073
rect 11158 10962 11186 11047
rect 11158 10929 11186 10934
rect 11718 10962 11746 11103
rect 11718 10929 11746 10934
rect 11774 11018 11802 11774
rect 12670 11689 12698 11774
rect 12670 11663 12671 11689
rect 12697 11663 12698 11689
rect 12670 11657 12698 11663
rect 12726 12361 12866 12362
rect 12726 12335 12839 12361
rect 12865 12335 12866 12361
rect 12726 12334 12866 12335
rect 12334 11522 12362 11527
rect 12054 11521 12362 11522
rect 12054 11495 12335 11521
rect 12361 11495 12362 11521
rect 12054 11494 12362 11495
rect 11886 11242 11914 11247
rect 11886 11129 11914 11214
rect 11886 11103 11887 11129
rect 11913 11103 11914 11129
rect 11886 11097 11914 11103
rect 12054 11185 12082 11494
rect 12334 11489 12362 11494
rect 12054 11159 12055 11185
rect 12081 11159 12082 11185
rect 11830 11074 11858 11079
rect 11830 11018 11858 11046
rect 11774 10990 11858 11018
rect 10934 10737 10962 10743
rect 10934 10711 10935 10737
rect 10961 10711 10962 10737
rect 10934 10514 10962 10711
rect 10934 10481 10962 10486
rect 11382 10458 11410 10463
rect 11382 10411 11410 10430
rect 11662 10458 11690 10463
rect 11102 10402 11130 10407
rect 11130 10374 11298 10402
rect 11102 10355 11130 10374
rect 10822 10033 10850 10038
rect 11046 10010 11074 10015
rect 11270 10010 11298 10374
rect 11382 10122 11410 10127
rect 11382 10065 11410 10094
rect 11382 10039 11383 10065
rect 11409 10039 11410 10065
rect 11382 10033 11410 10039
rect 11662 10065 11690 10430
rect 11662 10039 11663 10065
rect 11689 10039 11690 10065
rect 11662 10033 11690 10039
rect 11774 10289 11802 10990
rect 11886 10682 11914 10687
rect 11886 10401 11914 10654
rect 11886 10375 11887 10401
rect 11913 10375 11914 10401
rect 11886 10369 11914 10375
rect 11942 10402 11970 10407
rect 11774 10263 11775 10289
rect 11801 10263 11802 10289
rect 11046 9963 11074 9982
rect 11214 10009 11298 10010
rect 11214 9983 11271 10009
rect 11297 9983 11298 10009
rect 11214 9982 11298 9983
rect 10878 9953 10906 9959
rect 10878 9927 10879 9953
rect 10905 9927 10906 9953
rect 10878 9898 10906 9927
rect 10878 9865 10906 9870
rect 10766 9647 10767 9673
rect 10793 9647 10794 9673
rect 10766 9641 10794 9647
rect 10822 9617 10850 9623
rect 10822 9591 10823 9617
rect 10849 9591 10850 9617
rect 10822 9506 10850 9591
rect 11214 9618 11242 9982
rect 11270 9977 11298 9982
rect 11606 10010 11634 10015
rect 11606 9963 11634 9982
rect 10822 9473 10850 9478
rect 10990 9505 11018 9511
rect 10990 9479 10991 9505
rect 11017 9479 11018 9505
rect 10654 9366 10850 9394
rect 10094 9199 10095 9225
rect 10121 9199 10122 9225
rect 10094 9170 10122 9199
rect 9590 8441 9618 9142
rect 10094 9137 10122 9142
rect 10710 9281 10738 9287
rect 10710 9255 10711 9281
rect 10737 9255 10738 9281
rect 9702 8833 9730 8839
rect 9702 8807 9703 8833
rect 9729 8807 9730 8833
rect 9702 8722 9730 8807
rect 9702 8689 9730 8694
rect 10654 8777 10682 8783
rect 10654 8751 10655 8777
rect 10681 8751 10682 8777
rect 9918 8638 10050 8643
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 9918 8605 10050 8610
rect 10654 8498 10682 8751
rect 10710 8554 10738 9255
rect 10822 9226 10850 9366
rect 10822 9179 10850 9198
rect 10990 9170 11018 9479
rect 11158 9506 11186 9511
rect 11158 9459 11186 9478
rect 11102 9338 11130 9343
rect 10934 9114 10962 9119
rect 10822 8722 10850 8727
rect 10710 8526 10794 8554
rect 10654 8470 10738 8498
rect 9590 8415 9591 8441
rect 9617 8415 9618 8441
rect 9590 8409 9618 8415
rect 10654 8385 10682 8391
rect 10654 8359 10655 8385
rect 10681 8359 10682 8385
rect 9478 8246 9618 8274
rect 9422 8135 9423 8161
rect 9449 8135 9450 8161
rect 9422 8129 9450 8135
rect 9590 8161 9618 8246
rect 9590 8135 9591 8161
rect 9617 8135 9618 8161
rect 9590 8129 9618 8135
rect 10654 8106 10682 8359
rect 10710 8162 10738 8470
rect 10766 8442 10794 8526
rect 10766 8409 10794 8414
rect 10710 8115 10738 8134
rect 10822 8161 10850 8694
rect 10822 8135 10823 8161
rect 10849 8135 10850 8161
rect 10822 8129 10850 8135
rect 10934 8666 10962 9086
rect 10990 8833 11018 9142
rect 10990 8807 10991 8833
rect 11017 8807 11018 8833
rect 10990 8801 11018 8807
rect 11046 9281 11074 9287
rect 11046 9255 11047 9281
rect 11073 9255 11074 9281
rect 10990 8666 11018 8671
rect 10934 8638 10990 8666
rect 9478 7938 9506 7943
rect 9478 7891 9506 7910
rect 10150 7938 10178 7943
rect 9918 7854 10050 7859
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 9918 7821 10050 7826
rect 9254 7239 9255 7265
rect 9281 7239 9282 7265
rect 9254 7233 9282 7239
rect 10094 7602 10122 7607
rect 8582 7154 8610 7159
rect 8582 7107 8610 7126
rect 9142 7153 9170 7159
rect 9142 7127 9143 7153
rect 9169 7127 9170 7153
rect 9142 6538 9170 7127
rect 9918 7070 10050 7075
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 9918 7037 10050 7042
rect 9198 6538 9226 6543
rect 9142 6537 9226 6538
rect 9142 6511 9199 6537
rect 9225 6511 9226 6537
rect 9142 6510 9226 6511
rect 9198 4214 9226 6510
rect 10094 6538 10122 7574
rect 10094 6505 10122 6510
rect 10150 7601 10178 7910
rect 10150 7575 10151 7601
rect 10177 7575 10178 7601
rect 9478 6482 9506 6487
rect 9478 6435 9506 6454
rect 9918 6286 10050 6291
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 9918 6253 10050 6258
rect 9918 5502 10050 5507
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 9918 5469 10050 5474
rect 9918 4718 10050 4723
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 9918 4685 10050 4690
rect 8414 4186 8722 4214
rect 2238 3542 2370 3547
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2238 3509 2370 3514
rect 2238 2758 2370 2763
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2238 2725 2370 2730
rect 8694 2169 8722 4186
rect 8694 2143 8695 2169
rect 8721 2143 8722 2169
rect 8694 2137 8722 2143
rect 8806 4186 9226 4214
rect 10150 4214 10178 7575
rect 10374 7602 10402 7621
rect 10374 7569 10402 7574
rect 10654 7602 10682 8078
rect 10934 8105 10962 8638
rect 10990 8633 11018 8638
rect 11046 8554 11074 9255
rect 11102 8889 11130 9310
rect 11214 9337 11242 9590
rect 11214 9311 11215 9337
rect 11241 9311 11242 9337
rect 11214 9305 11242 9311
rect 11438 9897 11466 9903
rect 11438 9871 11439 9897
rect 11465 9871 11466 9897
rect 11438 9505 11466 9871
rect 11606 9674 11634 9679
rect 11606 9617 11634 9646
rect 11774 9618 11802 10263
rect 11942 10065 11970 10374
rect 11942 10039 11943 10065
rect 11969 10039 11970 10065
rect 11942 10033 11970 10039
rect 12054 9674 12082 11159
rect 12726 11186 12754 12334
rect 12838 12329 12866 12334
rect 12950 12361 12978 12367
rect 12950 12335 12951 12361
rect 12977 12335 12978 12361
rect 12950 12082 12978 12335
rect 13174 12361 13202 13006
rect 13174 12335 13175 12361
rect 13201 12335 13202 12361
rect 13174 12329 13202 12335
rect 13286 12838 13426 12866
rect 12054 9627 12082 9646
rect 12166 10962 12194 10967
rect 11606 9591 11607 9617
rect 11633 9591 11634 9617
rect 11606 9585 11634 9591
rect 11718 9590 11802 9618
rect 11830 9618 11858 9623
rect 11438 9479 11439 9505
rect 11465 9479 11466 9505
rect 11438 9338 11466 9479
rect 11438 9305 11466 9310
rect 11606 9394 11634 9399
rect 11718 9394 11746 9590
rect 11830 9571 11858 9590
rect 11774 9506 11802 9511
rect 11774 9459 11802 9478
rect 11998 9505 12026 9511
rect 11998 9479 11999 9505
rect 12025 9479 12026 9505
rect 11998 9394 12026 9479
rect 11718 9366 11802 9394
rect 11382 9226 11410 9231
rect 11382 9179 11410 9198
rect 11606 9226 11634 9366
rect 11606 9225 11690 9226
rect 11606 9199 11607 9225
rect 11633 9199 11690 9225
rect 11606 9198 11690 9199
rect 11606 9193 11634 9198
rect 11102 8863 11103 8889
rect 11129 8863 11130 8889
rect 11102 8857 11130 8863
rect 11662 8833 11690 9198
rect 11774 9114 11802 9366
rect 11998 9361 12026 9366
rect 12054 9506 12082 9511
rect 11830 9338 11858 9343
rect 11830 9225 11858 9310
rect 11998 9282 12026 9287
rect 12054 9282 12082 9478
rect 11998 9281 12138 9282
rect 11998 9255 11999 9281
rect 12025 9255 12138 9281
rect 11998 9254 12138 9255
rect 11998 9249 12026 9254
rect 11830 9199 11831 9225
rect 11857 9199 11858 9225
rect 11830 9193 11858 9199
rect 11774 9086 12026 9114
rect 11662 8807 11663 8833
rect 11689 8807 11690 8833
rect 11662 8801 11690 8807
rect 11998 8833 12026 9086
rect 11998 8807 11999 8833
rect 12025 8807 12026 8833
rect 11998 8801 12026 8807
rect 12110 8834 12138 9254
rect 12110 8801 12138 8806
rect 11550 8778 11578 8783
rect 11550 8731 11578 8750
rect 11942 8778 11970 8783
rect 11942 8731 11970 8750
rect 11046 8521 11074 8526
rect 11438 8722 11466 8727
rect 10934 8079 10935 8105
rect 10961 8079 10962 8105
rect 10934 8073 10962 8079
rect 10990 8442 11018 8447
rect 10654 7266 10682 7574
rect 10990 7378 11018 8414
rect 11382 8162 11410 8167
rect 11382 8049 11410 8134
rect 11382 8023 11383 8049
rect 11409 8023 11410 8049
rect 11382 8017 11410 8023
rect 11438 7993 11466 8694
rect 11830 8722 11858 8727
rect 12166 8722 12194 10934
rect 12670 10849 12698 10855
rect 12670 10823 12671 10849
rect 12697 10823 12698 10849
rect 12614 10793 12642 10799
rect 12614 10767 12615 10793
rect 12641 10767 12642 10793
rect 12614 10122 12642 10767
rect 12670 10682 12698 10823
rect 12670 10649 12698 10654
rect 12726 10402 12754 11158
rect 12838 12054 12978 12082
rect 12838 11074 12866 12054
rect 12894 11970 12922 11975
rect 13286 11970 13314 12838
rect 13398 12810 13426 12838
rect 13510 12810 13538 13118
rect 13566 13034 13594 13039
rect 13566 12987 13594 13006
rect 13398 12782 13538 12810
rect 13622 12810 13650 13174
rect 18830 13145 18858 13151
rect 18830 13119 18831 13145
rect 18857 13119 18858 13145
rect 14518 13090 14546 13095
rect 14518 13043 14546 13062
rect 14966 13090 14994 13095
rect 14462 13033 14490 13039
rect 14462 13007 14463 13033
rect 14489 13007 14490 13033
rect 13678 12810 13706 12815
rect 13622 12782 13678 12810
rect 13678 12777 13706 12782
rect 14070 12810 14098 12815
rect 14070 12763 14098 12782
rect 13342 12754 13370 12759
rect 13342 12474 13370 12726
rect 13342 12427 13370 12446
rect 13398 12698 13426 12703
rect 13342 11970 13370 11975
rect 13286 11969 13370 11970
rect 13286 11943 13343 11969
rect 13369 11943 13370 11969
rect 13286 11942 13370 11943
rect 12894 11241 12922 11942
rect 13342 11937 13370 11942
rect 13398 11913 13426 12670
rect 14462 12698 14490 13007
rect 14462 12665 14490 12670
rect 13510 12474 13538 12479
rect 13510 12361 13538 12446
rect 13510 12335 13511 12361
rect 13537 12335 13538 12361
rect 13510 12329 13538 12335
rect 13902 12306 13930 12311
rect 13846 12305 13930 12306
rect 13846 12279 13903 12305
rect 13929 12279 13930 12305
rect 13846 12278 13930 12279
rect 13622 11970 13650 11975
rect 13622 11923 13650 11942
rect 13734 11969 13762 11975
rect 13734 11943 13735 11969
rect 13761 11943 13762 11969
rect 13398 11887 13399 11913
rect 13425 11887 13426 11913
rect 13398 11881 13426 11887
rect 13510 11858 13538 11863
rect 13734 11858 13762 11943
rect 13510 11857 13762 11858
rect 13510 11831 13511 11857
rect 13537 11831 13762 11857
rect 13510 11830 13762 11831
rect 13846 11858 13874 12278
rect 13902 12273 13930 12278
rect 14966 12305 14994 13062
rect 17598 12950 17730 12955
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17598 12917 17730 12922
rect 18830 12810 18858 13119
rect 18942 13090 18970 13511
rect 20006 13146 20034 13567
rect 20006 13113 20034 13118
rect 18942 13057 18970 13062
rect 18830 12777 18858 12782
rect 20006 13033 20034 13039
rect 20006 13007 20007 13033
rect 20033 13007 20034 13033
rect 20006 12810 20034 13007
rect 20006 12777 20034 12782
rect 14966 12279 14967 12305
rect 14993 12279 14994 12305
rect 14966 12273 14994 12279
rect 17598 12166 17730 12171
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17598 12133 17730 12138
rect 13902 11970 13930 11975
rect 14182 11970 14210 11975
rect 13902 11969 14210 11970
rect 13902 11943 13903 11969
rect 13929 11943 14183 11969
rect 14209 11943 14210 11969
rect 13902 11942 14210 11943
rect 13902 11937 13930 11942
rect 14182 11937 14210 11942
rect 14070 11858 14098 11863
rect 13846 11857 14098 11858
rect 13846 11831 14071 11857
rect 14097 11831 14098 11857
rect 13846 11830 14098 11831
rect 13510 11825 13538 11830
rect 14070 11825 14098 11830
rect 12894 11215 12895 11241
rect 12921 11215 12922 11241
rect 12894 11209 12922 11215
rect 13118 11802 13146 11807
rect 12838 11027 12866 11046
rect 12894 11129 12922 11135
rect 12894 11103 12895 11129
rect 12921 11103 12922 11129
rect 12894 10962 12922 11103
rect 12950 11130 12978 11135
rect 12950 11083 12978 11102
rect 12782 10934 12922 10962
rect 12782 10905 12810 10934
rect 12782 10879 12783 10905
rect 12809 10879 12810 10905
rect 12782 10873 12810 10879
rect 12894 10570 12922 10934
rect 13118 10906 13146 11774
rect 13622 11577 13650 11583
rect 13622 11551 13623 11577
rect 13649 11551 13650 11577
rect 13622 11186 13650 11551
rect 13622 11153 13650 11158
rect 13734 11521 13762 11527
rect 13734 11495 13735 11521
rect 13761 11495 13762 11521
rect 13174 10906 13202 10911
rect 13118 10905 13370 10906
rect 13118 10879 13175 10905
rect 13201 10879 13370 10905
rect 13118 10878 13370 10879
rect 13174 10873 13202 10878
rect 13342 10793 13370 10878
rect 13734 10849 13762 11495
rect 13790 11466 13818 11471
rect 13790 11465 13986 11466
rect 13790 11439 13791 11465
rect 13817 11439 13986 11465
rect 13790 11438 13986 11439
rect 13790 11433 13818 11438
rect 13958 11241 13986 11438
rect 17598 11382 17730 11387
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17598 11349 17730 11354
rect 13958 11215 13959 11241
rect 13985 11215 13986 11241
rect 13958 11209 13986 11215
rect 20006 11241 20034 11247
rect 20006 11215 20007 11241
rect 20033 11215 20034 11241
rect 14070 11186 14098 11191
rect 14070 11139 14098 11158
rect 14798 11186 14826 11191
rect 13734 10823 13735 10849
rect 13761 10823 13762 10849
rect 13734 10817 13762 10823
rect 13902 11129 13930 11135
rect 13902 11103 13903 11129
rect 13929 11103 13930 11129
rect 13342 10767 13343 10793
rect 13369 10767 13370 10793
rect 13342 10761 13370 10767
rect 12894 10542 12978 10570
rect 12894 10458 12922 10463
rect 12894 10411 12922 10430
rect 12726 10355 12754 10374
rect 12950 10401 12978 10542
rect 13230 10458 13258 10463
rect 13258 10430 13314 10458
rect 13230 10425 13258 10430
rect 12950 10375 12951 10401
rect 12977 10375 12978 10401
rect 12950 10369 12978 10375
rect 13118 10401 13146 10407
rect 13118 10375 13119 10401
rect 13145 10375 13146 10401
rect 12838 10346 12866 10351
rect 12614 10089 12642 10094
rect 12782 10345 12866 10346
rect 12782 10319 12839 10345
rect 12865 10319 12866 10345
rect 12782 10318 12866 10319
rect 12782 10066 12810 10318
rect 12838 10313 12866 10318
rect 12726 10038 12810 10066
rect 11830 8675 11858 8694
rect 12110 8694 12194 8722
rect 12614 8778 12642 8783
rect 11886 8106 11914 8111
rect 11886 8059 11914 8078
rect 12054 8106 12082 8111
rect 12110 8106 12138 8694
rect 12614 8553 12642 8750
rect 12726 8666 12754 10038
rect 12950 10009 12978 10015
rect 12950 9983 12951 10009
rect 12977 9983 12978 10009
rect 12782 9954 12810 9959
rect 12950 9954 12978 9983
rect 12782 9953 12978 9954
rect 12782 9927 12783 9953
rect 12809 9927 12978 9953
rect 12782 9926 12978 9927
rect 12782 9921 12810 9926
rect 12726 8633 12754 8638
rect 12950 9170 12978 9926
rect 13118 9674 13146 10375
rect 13286 10065 13314 10430
rect 13286 10039 13287 10065
rect 13313 10039 13314 10065
rect 13286 10033 13314 10039
rect 13398 10066 13426 10071
rect 13118 9641 13146 9646
rect 13230 9898 13258 9903
rect 13230 9618 13258 9870
rect 13230 9571 13258 9590
rect 13398 9617 13426 10038
rect 13902 10066 13930 11103
rect 14798 10737 14826 11158
rect 18830 11186 18858 11191
rect 18830 11139 18858 11158
rect 20006 11130 20034 11215
rect 20006 11097 20034 11102
rect 14798 10711 14799 10737
rect 14825 10711 14826 10737
rect 14798 10705 14826 10711
rect 17598 10598 17730 10603
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17598 10565 17730 10570
rect 20006 10457 20034 10463
rect 20006 10431 20007 10457
rect 20033 10431 20034 10457
rect 18942 10401 18970 10407
rect 18942 10375 18943 10401
rect 18969 10375 18970 10401
rect 14686 10066 14714 10071
rect 13930 10038 14098 10066
rect 13902 10033 13930 10038
rect 13510 9954 13538 9959
rect 13454 9674 13482 9679
rect 13454 9627 13482 9646
rect 13398 9591 13399 9617
rect 13425 9591 13426 9617
rect 13398 9585 13426 9591
rect 13510 9617 13538 9926
rect 13510 9591 13511 9617
rect 13537 9591 13538 9617
rect 13510 9585 13538 9591
rect 13790 9618 13818 9623
rect 13790 9571 13818 9590
rect 14070 9617 14098 10038
rect 14686 10019 14714 10038
rect 18942 10066 18970 10375
rect 20006 10122 20034 10431
rect 20006 10089 20034 10094
rect 18942 10033 18970 10038
rect 14574 10010 14602 10015
rect 14350 9982 14574 10010
rect 14350 9954 14378 9982
rect 14574 9963 14602 9982
rect 18830 10010 18858 10015
rect 18830 9963 18858 9982
rect 14350 9907 14378 9926
rect 20006 9897 20034 9903
rect 20006 9871 20007 9897
rect 20033 9871 20034 9897
rect 17598 9814 17730 9819
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17598 9781 17730 9786
rect 20006 9786 20034 9871
rect 20006 9753 20034 9758
rect 20006 9673 20034 9679
rect 20006 9647 20007 9673
rect 20033 9647 20034 9673
rect 14070 9591 14071 9617
rect 14097 9591 14098 9617
rect 14070 9585 14098 9591
rect 18830 9617 18858 9623
rect 18830 9591 18831 9617
rect 18857 9591 18858 9617
rect 14014 9562 14042 9567
rect 14014 9515 14042 9534
rect 14574 9561 14602 9567
rect 14574 9535 14575 9561
rect 14601 9535 14602 9561
rect 13622 9506 13650 9511
rect 13622 9459 13650 9478
rect 13902 9505 13930 9511
rect 13902 9479 13903 9505
rect 13929 9479 13930 9505
rect 13902 9338 13930 9479
rect 14574 9506 14602 9535
rect 14742 9562 14770 9567
rect 14742 9515 14770 9534
rect 14574 9473 14602 9478
rect 14630 9505 14658 9511
rect 14630 9479 14631 9505
rect 14657 9479 14658 9505
rect 13510 9310 13930 9338
rect 13510 9281 13538 9310
rect 13510 9255 13511 9281
rect 13537 9255 13538 9281
rect 13510 9249 13538 9255
rect 14574 9282 14602 9287
rect 14630 9282 14658 9479
rect 14602 9254 14658 9282
rect 18830 9282 18858 9591
rect 20006 9450 20034 9647
rect 20006 9417 20034 9422
rect 13118 9225 13146 9231
rect 13118 9199 13119 9225
rect 13145 9199 13146 9225
rect 13118 9170 13146 9199
rect 12950 9169 13146 9170
rect 12950 9143 12951 9169
rect 12977 9143 13146 9169
rect 12950 9142 13146 9143
rect 14574 9169 14602 9254
rect 18830 9249 18858 9254
rect 14574 9143 14575 9169
rect 14601 9143 14602 9169
rect 12614 8527 12615 8553
rect 12641 8527 12642 8553
rect 12614 8521 12642 8527
rect 12838 8554 12866 8559
rect 12838 8507 12866 8526
rect 12726 8498 12754 8503
rect 12726 8451 12754 8470
rect 12334 8442 12362 8447
rect 12166 8386 12194 8391
rect 12166 8161 12194 8358
rect 12166 8135 12167 8161
rect 12193 8135 12194 8161
rect 12166 8129 12194 8135
rect 12334 8161 12362 8414
rect 12670 8386 12698 8391
rect 12670 8339 12698 8358
rect 12334 8135 12335 8161
rect 12361 8135 12362 8161
rect 12334 8129 12362 8135
rect 12054 8105 12138 8106
rect 12054 8079 12055 8105
rect 12081 8079 12138 8105
rect 12054 8078 12138 8079
rect 12222 8106 12250 8111
rect 12054 8073 12082 8078
rect 11550 7994 11578 7999
rect 11438 7967 11439 7993
rect 11465 7967 11466 7993
rect 11438 7961 11466 7967
rect 11494 7993 11634 7994
rect 11494 7967 11551 7993
rect 11577 7967 11634 7993
rect 11494 7966 11634 7967
rect 11046 7938 11074 7943
rect 11046 7891 11074 7910
rect 11102 7937 11130 7943
rect 11102 7911 11103 7937
rect 11129 7911 11130 7937
rect 10990 7345 11018 7350
rect 11046 7322 11074 7327
rect 11102 7322 11130 7911
rect 11158 7938 11186 7943
rect 11494 7938 11522 7966
rect 11550 7961 11578 7966
rect 11158 7937 11354 7938
rect 11158 7911 11159 7937
rect 11185 7911 11354 7937
rect 11158 7910 11354 7911
rect 11158 7905 11186 7910
rect 11326 7769 11354 7910
rect 11494 7905 11522 7910
rect 11326 7743 11327 7769
rect 11353 7743 11354 7769
rect 11326 7737 11354 7743
rect 11606 7713 11634 7966
rect 12222 7769 12250 8078
rect 12222 7743 12223 7769
rect 12249 7743 12250 7769
rect 12222 7737 12250 7743
rect 12558 8106 12586 8111
rect 12558 8049 12586 8078
rect 12950 8106 12978 9142
rect 14574 9137 14602 9143
rect 17598 9030 17730 9035
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17598 8997 17730 9002
rect 20006 8889 20034 8895
rect 20006 8863 20007 8889
rect 20033 8863 20034 8889
rect 18942 8833 18970 8839
rect 18942 8807 18943 8833
rect 18969 8807 18970 8833
rect 13678 8497 13706 8503
rect 13678 8471 13679 8497
rect 13705 8471 13706 8497
rect 13118 8442 13146 8447
rect 13118 8395 13146 8414
rect 13566 8442 13594 8447
rect 13062 8330 13090 8335
rect 12950 8073 12978 8078
rect 13006 8329 13090 8330
rect 13006 8303 13063 8329
rect 13089 8303 13090 8329
rect 13006 8302 13090 8303
rect 12558 8023 12559 8049
rect 12585 8023 12586 8049
rect 11606 7687 11607 7713
rect 11633 7687 11634 7713
rect 11606 7681 11634 7687
rect 11438 7658 11466 7663
rect 11438 7611 11466 7630
rect 11774 7658 11802 7663
rect 11774 7657 12362 7658
rect 11774 7631 11775 7657
rect 11801 7631 12362 7657
rect 11774 7630 12362 7631
rect 11774 7625 11802 7630
rect 11270 7601 11298 7607
rect 11270 7575 11271 7601
rect 11297 7575 11298 7601
rect 11270 7378 11298 7575
rect 11270 7345 11298 7350
rect 11662 7601 11690 7607
rect 11662 7575 11663 7601
rect 11689 7575 11690 7601
rect 11046 7321 11130 7322
rect 11046 7295 11047 7321
rect 11073 7295 11130 7321
rect 11046 7294 11130 7295
rect 11046 7289 11074 7294
rect 10654 7265 10906 7266
rect 10654 7239 10655 7265
rect 10681 7239 10906 7265
rect 10654 7238 10906 7239
rect 10654 7233 10682 7238
rect 10878 6873 10906 7238
rect 11662 7210 11690 7575
rect 11270 7182 11690 7210
rect 12110 7546 12138 7551
rect 12110 7321 12138 7518
rect 12278 7378 12306 7383
rect 12278 7331 12306 7350
rect 12110 7295 12111 7321
rect 12137 7295 12138 7321
rect 11270 6929 11298 7182
rect 11270 6903 11271 6929
rect 11297 6903 11298 6929
rect 11270 6897 11298 6903
rect 10878 6847 10879 6873
rect 10905 6847 10906 6873
rect 10878 6841 10906 6847
rect 12110 4214 12138 7295
rect 12334 7321 12362 7630
rect 12558 7574 12586 8023
rect 12950 7994 12978 7999
rect 13006 7994 13034 8302
rect 13062 8297 13090 8302
rect 12950 7993 13034 7994
rect 12950 7967 12951 7993
rect 12977 7967 13034 7993
rect 12950 7966 13034 7967
rect 12950 7961 12978 7966
rect 13566 7657 13594 8414
rect 13678 8386 13706 8471
rect 13678 8353 13706 8358
rect 14070 8442 14098 8447
rect 14070 8105 14098 8414
rect 18830 8441 18858 8447
rect 18830 8415 18831 8441
rect 18857 8415 18858 8441
rect 18830 8386 18858 8415
rect 18942 8442 18970 8807
rect 18942 8409 18970 8414
rect 20006 8442 20034 8863
rect 20006 8409 20034 8414
rect 18830 8353 18858 8358
rect 19950 8385 19978 8391
rect 19950 8359 19951 8385
rect 19977 8359 19978 8385
rect 17598 8246 17730 8251
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17598 8213 17730 8218
rect 14070 8079 14071 8105
rect 14097 8079 14098 8105
rect 14070 8073 14098 8079
rect 19950 8106 19978 8359
rect 19950 8073 19978 8078
rect 20006 8105 20034 8111
rect 20006 8079 20007 8105
rect 20033 8079 20034 8105
rect 18830 8049 18858 8055
rect 18830 8023 18831 8049
rect 18857 8023 18858 8049
rect 13678 7714 13706 7719
rect 13678 7667 13706 7686
rect 18830 7714 18858 8023
rect 20006 7770 20034 8079
rect 20006 7737 20034 7742
rect 18830 7681 18858 7686
rect 13566 7631 13567 7657
rect 13593 7631 13594 7657
rect 13566 7625 13594 7631
rect 12558 7546 12698 7574
rect 12334 7295 12335 7321
rect 12361 7295 12362 7321
rect 12334 7289 12362 7295
rect 12390 7154 12418 7159
rect 12614 7154 12642 7159
rect 12390 7153 12642 7154
rect 12390 7127 12391 7153
rect 12417 7127 12615 7153
rect 12641 7127 12642 7153
rect 12390 7126 12642 7127
rect 12334 6818 12362 6823
rect 12390 6818 12418 7126
rect 12614 7121 12642 7126
rect 12670 6985 12698 7546
rect 17598 7462 17730 7467
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17598 7429 17730 7434
rect 12670 6959 12671 6985
rect 12697 6959 12698 6985
rect 12670 6953 12698 6959
rect 12782 7153 12810 7159
rect 12782 7127 12783 7153
rect 12809 7127 12810 7153
rect 12334 6817 12418 6818
rect 12334 6791 12335 6817
rect 12361 6791 12418 6817
rect 12334 6790 12418 6791
rect 12334 6762 12362 6790
rect 12334 6729 12362 6734
rect 12782 4214 12810 7127
rect 10150 4186 10402 4214
rect 12110 4186 12306 4214
rect 8414 2058 8442 2063
rect 2238 1974 2370 1979
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2238 1941 2370 1946
rect 8414 400 8442 2030
rect 8806 1777 8834 4186
rect 9918 3934 10050 3939
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 9918 3901 10050 3906
rect 9918 3150 10050 3155
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 9918 3117 10050 3122
rect 9918 2366 10050 2371
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 9918 2333 10050 2338
rect 9198 2058 9226 2063
rect 9198 2011 9226 2030
rect 9310 1834 9338 1839
rect 8806 1751 8807 1777
rect 8833 1751 8834 1777
rect 8806 1745 8834 1751
rect 9086 1833 9338 1834
rect 9086 1807 9311 1833
rect 9337 1807 9338 1833
rect 9086 1806 9338 1807
rect 9086 400 9114 1806
rect 9310 1801 9338 1806
rect 9758 1834 9786 1839
rect 9758 400 9786 1806
rect 10374 1777 10402 4186
rect 11998 2618 12026 2623
rect 11830 2617 12026 2618
rect 11830 2591 11999 2617
rect 12025 2591 12026 2617
rect 11830 2590 12026 2591
rect 10934 1834 10962 1839
rect 10934 1787 10962 1806
rect 11438 1834 11466 1839
rect 10374 1751 10375 1777
rect 10401 1751 10402 1777
rect 10374 1745 10402 1751
rect 9918 1582 10050 1587
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 9918 1549 10050 1554
rect 11438 400 11466 1806
rect 11830 490 11858 2590
rect 11998 2585 12026 2590
rect 12278 1777 12306 4186
rect 12614 4186 12810 4214
rect 12950 6762 12978 6767
rect 12614 2169 12642 4186
rect 12950 2561 12978 6734
rect 17598 6678 17730 6683
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17598 6645 17730 6650
rect 17598 5894 17730 5899
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17598 5861 17730 5866
rect 17598 5110 17730 5115
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17598 5077 17730 5082
rect 17598 4326 17730 4331
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17598 4293 17730 4298
rect 17598 3542 17730 3547
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17598 3509 17730 3514
rect 17598 2758 17730 2763
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17598 2725 17730 2730
rect 12950 2535 12951 2561
rect 12977 2535 12978 2561
rect 12950 2529 12978 2535
rect 12614 2143 12615 2169
rect 12641 2143 12642 2169
rect 12614 2137 12642 2143
rect 12278 1751 12279 1777
rect 12305 1751 12306 1777
rect 12278 1745 12306 1751
rect 12446 2058 12474 2063
rect 11774 462 11858 490
rect 11774 400 11802 462
rect 12446 400 12474 2030
rect 13118 2058 13146 2063
rect 13118 2011 13146 2030
rect 17598 1974 17730 1979
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17598 1941 17730 1946
rect 12782 1834 12810 1839
rect 12782 1787 12810 1806
rect 8400 0 8456 400
rect 9072 0 9128 400
rect 9744 0 9800 400
rect 11424 0 11480 400
rect 11760 0 11816 400
rect 12432 0 12488 400
<< via2 >>
rect 2238 19221 2266 19222
rect 2238 19195 2239 19221
rect 2239 19195 2265 19221
rect 2265 19195 2266 19221
rect 2238 19194 2266 19195
rect 2290 19221 2318 19222
rect 2290 19195 2291 19221
rect 2291 19195 2317 19221
rect 2317 19195 2318 19221
rect 2290 19194 2318 19195
rect 2342 19221 2370 19222
rect 2342 19195 2343 19221
rect 2343 19195 2369 19221
rect 2369 19195 2370 19221
rect 2342 19194 2370 19195
rect 2238 18437 2266 18438
rect 2238 18411 2239 18437
rect 2239 18411 2265 18437
rect 2265 18411 2266 18437
rect 2238 18410 2266 18411
rect 2290 18437 2318 18438
rect 2290 18411 2291 18437
rect 2291 18411 2317 18437
rect 2317 18411 2318 18437
rect 2290 18410 2318 18411
rect 2342 18437 2370 18438
rect 2342 18411 2343 18437
rect 2343 18411 2369 18437
rect 2369 18411 2370 18437
rect 2342 18410 2370 18411
rect 8750 18718 8778 18746
rect 2238 17653 2266 17654
rect 2238 17627 2239 17653
rect 2239 17627 2265 17653
rect 2265 17627 2266 17653
rect 2238 17626 2266 17627
rect 2290 17653 2318 17654
rect 2290 17627 2291 17653
rect 2291 17627 2317 17653
rect 2317 17627 2318 17653
rect 2290 17626 2318 17627
rect 2342 17653 2370 17654
rect 2342 17627 2343 17653
rect 2343 17627 2369 17653
rect 2369 17627 2370 17653
rect 2342 17626 2370 17627
rect 2238 16869 2266 16870
rect 2238 16843 2239 16869
rect 2239 16843 2265 16869
rect 2265 16843 2266 16869
rect 2238 16842 2266 16843
rect 2290 16869 2318 16870
rect 2290 16843 2291 16869
rect 2291 16843 2317 16869
rect 2317 16843 2318 16869
rect 2290 16842 2318 16843
rect 2342 16869 2370 16870
rect 2342 16843 2343 16869
rect 2343 16843 2369 16869
rect 2369 16843 2370 16869
rect 2342 16842 2370 16843
rect 2238 16085 2266 16086
rect 2238 16059 2239 16085
rect 2239 16059 2265 16085
rect 2265 16059 2266 16085
rect 2238 16058 2266 16059
rect 2290 16085 2318 16086
rect 2290 16059 2291 16085
rect 2291 16059 2317 16085
rect 2317 16059 2318 16085
rect 2290 16058 2318 16059
rect 2342 16085 2370 16086
rect 2342 16059 2343 16085
rect 2343 16059 2369 16085
rect 2369 16059 2370 16085
rect 2342 16058 2370 16059
rect 9918 18829 9946 18830
rect 9918 18803 9919 18829
rect 9919 18803 9945 18829
rect 9945 18803 9946 18829
rect 9918 18802 9946 18803
rect 9970 18829 9998 18830
rect 9970 18803 9971 18829
rect 9971 18803 9997 18829
rect 9997 18803 9998 18829
rect 9970 18802 9998 18803
rect 10022 18829 10050 18830
rect 10022 18803 10023 18829
rect 10023 18803 10049 18829
rect 10049 18803 10050 18829
rect 10022 18802 10050 18803
rect 9366 18745 9394 18746
rect 9366 18719 9367 18745
rect 9367 18719 9393 18745
rect 9393 18719 9394 18745
rect 9366 18718 9394 18719
rect 2238 15301 2266 15302
rect 2238 15275 2239 15301
rect 2239 15275 2265 15301
rect 2265 15275 2266 15301
rect 2238 15274 2266 15275
rect 2290 15301 2318 15302
rect 2290 15275 2291 15301
rect 2291 15275 2317 15301
rect 2317 15275 2318 15301
rect 2290 15274 2318 15275
rect 2342 15301 2370 15302
rect 2342 15275 2343 15301
rect 2343 15275 2369 15301
rect 2369 15275 2370 15301
rect 2342 15274 2370 15275
rect 2238 14517 2266 14518
rect 2238 14491 2239 14517
rect 2239 14491 2265 14517
rect 2265 14491 2266 14517
rect 2238 14490 2266 14491
rect 2290 14517 2318 14518
rect 2290 14491 2291 14517
rect 2291 14491 2317 14517
rect 2317 14491 2318 14517
rect 2290 14490 2318 14491
rect 2342 14517 2370 14518
rect 2342 14491 2343 14517
rect 2343 14491 2369 14517
rect 2369 14491 2370 14517
rect 2342 14490 2370 14491
rect 8526 14321 8554 14322
rect 8526 14295 8527 14321
rect 8527 14295 8553 14321
rect 8553 14295 8554 14321
rect 8526 14294 8554 14295
rect 7686 14238 7714 14266
rect 7014 13929 7042 13930
rect 7014 13903 7015 13929
rect 7015 13903 7041 13929
rect 7041 13903 7042 13929
rect 7014 13902 7042 13903
rect 9918 18045 9946 18046
rect 9918 18019 9919 18045
rect 9919 18019 9945 18045
rect 9945 18019 9946 18045
rect 9918 18018 9946 18019
rect 9970 18045 9998 18046
rect 9970 18019 9971 18045
rect 9971 18019 9997 18045
rect 9997 18019 9998 18045
rect 9970 18018 9998 18019
rect 10022 18045 10050 18046
rect 10022 18019 10023 18045
rect 10023 18019 10049 18045
rect 10049 18019 10050 18045
rect 10022 18018 10050 18019
rect 9918 17261 9946 17262
rect 9918 17235 9919 17261
rect 9919 17235 9945 17261
rect 9945 17235 9946 17261
rect 9918 17234 9946 17235
rect 9970 17261 9998 17262
rect 9970 17235 9971 17261
rect 9971 17235 9997 17261
rect 9997 17235 9998 17261
rect 9970 17234 9998 17235
rect 10022 17261 10050 17262
rect 10022 17235 10023 17261
rect 10023 17235 10049 17261
rect 10049 17235 10050 17261
rect 10022 17234 10050 17235
rect 9918 16477 9946 16478
rect 9918 16451 9919 16477
rect 9919 16451 9945 16477
rect 9945 16451 9946 16477
rect 9918 16450 9946 16451
rect 9970 16477 9998 16478
rect 9970 16451 9971 16477
rect 9971 16451 9997 16477
rect 9997 16451 9998 16477
rect 9970 16450 9998 16451
rect 10022 16477 10050 16478
rect 10022 16451 10023 16477
rect 10023 16451 10049 16477
rect 10049 16451 10050 16477
rect 10022 16450 10050 16451
rect 7686 13902 7714 13930
rect 2086 13790 2114 13818
rect 966 13118 994 13146
rect 966 11774 994 11802
rect 2238 13733 2266 13734
rect 2238 13707 2239 13733
rect 2239 13707 2265 13733
rect 2265 13707 2266 13733
rect 2238 13706 2266 13707
rect 2290 13733 2318 13734
rect 2290 13707 2291 13733
rect 2291 13707 2317 13733
rect 2317 13707 2318 13733
rect 2290 13706 2318 13707
rect 2342 13733 2370 13734
rect 2342 13707 2343 13733
rect 2343 13707 2369 13733
rect 2369 13707 2370 13733
rect 2342 13706 2370 13707
rect 2142 13537 2170 13538
rect 2142 13511 2143 13537
rect 2143 13511 2169 13537
rect 2169 13511 2170 13537
rect 2142 13510 2170 13511
rect 6286 13510 6314 13538
rect 7350 13230 7378 13258
rect 8414 13873 8442 13874
rect 8414 13847 8415 13873
rect 8415 13847 8441 13873
rect 8441 13847 8442 13873
rect 8414 13846 8442 13847
rect 8134 13342 8162 13370
rect 7966 13257 7994 13258
rect 7966 13231 7967 13257
rect 7967 13231 7993 13257
rect 7993 13231 7994 13257
rect 7966 13230 7994 13231
rect 6286 13089 6314 13090
rect 6286 13063 6287 13089
rect 6287 13063 6313 13089
rect 6313 13063 6314 13089
rect 6286 13062 6314 13063
rect 2238 12949 2266 12950
rect 2238 12923 2239 12949
rect 2239 12923 2265 12949
rect 2265 12923 2266 12949
rect 2238 12922 2266 12923
rect 2290 12949 2318 12950
rect 2290 12923 2291 12949
rect 2291 12923 2317 12949
rect 2317 12923 2318 12949
rect 2290 12922 2318 12923
rect 2342 12949 2370 12950
rect 2342 12923 2343 12949
rect 2343 12923 2369 12949
rect 2369 12923 2370 12949
rect 2342 12922 2370 12923
rect 7350 12838 7378 12866
rect 7854 13062 7882 13090
rect 7910 12753 7938 12754
rect 7910 12727 7911 12753
rect 7911 12727 7937 12753
rect 7937 12727 7938 12753
rect 7910 12726 7938 12727
rect 9918 15693 9946 15694
rect 9918 15667 9919 15693
rect 9919 15667 9945 15693
rect 9945 15667 9946 15693
rect 9918 15666 9946 15667
rect 9970 15693 9998 15694
rect 9970 15667 9971 15693
rect 9971 15667 9997 15693
rect 9997 15667 9998 15693
rect 9970 15666 9998 15667
rect 10022 15693 10050 15694
rect 10022 15667 10023 15693
rect 10023 15667 10049 15693
rect 10049 15667 10050 15693
rect 10022 15666 10050 15667
rect 9918 14909 9946 14910
rect 9918 14883 9919 14909
rect 9919 14883 9945 14909
rect 9945 14883 9946 14909
rect 9918 14882 9946 14883
rect 9970 14909 9998 14910
rect 9970 14883 9971 14909
rect 9971 14883 9997 14909
rect 9997 14883 9998 14909
rect 9970 14882 9998 14883
rect 10022 14909 10050 14910
rect 10022 14883 10023 14909
rect 10023 14883 10049 14909
rect 10049 14883 10050 14909
rect 10022 14882 10050 14883
rect 9254 13846 9282 13874
rect 9198 13481 9226 13482
rect 9198 13455 9199 13481
rect 9199 13455 9225 13481
rect 9225 13455 9226 13481
rect 9198 13454 9226 13455
rect 9590 14238 9618 14266
rect 17598 19221 17626 19222
rect 17598 19195 17599 19221
rect 17599 19195 17625 19221
rect 17625 19195 17626 19221
rect 17598 19194 17626 19195
rect 17650 19221 17678 19222
rect 17650 19195 17651 19221
rect 17651 19195 17677 19221
rect 17677 19195 17678 19221
rect 17650 19194 17678 19195
rect 17702 19221 17730 19222
rect 17702 19195 17703 19221
rect 17703 19195 17729 19221
rect 17729 19195 17730 19221
rect 17702 19194 17730 19195
rect 12446 19110 12474 19138
rect 13062 19137 13090 19138
rect 13062 19111 13063 19137
rect 13063 19111 13089 19137
rect 13089 19111 13090 19137
rect 13062 19110 13090 19111
rect 10766 18718 10794 18746
rect 11382 18745 11410 18746
rect 11382 18719 11383 18745
rect 11383 18719 11409 18745
rect 11409 18719 11410 18745
rect 11382 18718 11410 18719
rect 10710 14630 10738 14658
rect 9918 14125 9946 14126
rect 9918 14099 9919 14125
rect 9919 14099 9945 14125
rect 9945 14099 9946 14125
rect 9918 14098 9946 14099
rect 9970 14125 9998 14126
rect 9970 14099 9971 14125
rect 9971 14099 9997 14125
rect 9997 14099 9998 14125
rect 9970 14098 9998 14099
rect 10022 14125 10050 14126
rect 10022 14099 10023 14125
rect 10023 14099 10049 14125
rect 10049 14099 10050 14125
rect 10022 14098 10050 14099
rect 9366 13481 9394 13482
rect 9366 13455 9367 13481
rect 9367 13455 9393 13481
rect 9393 13455 9394 13481
rect 9366 13454 9394 13455
rect 8806 13398 8834 13426
rect 8246 12838 8274 12866
rect 8190 12753 8218 12754
rect 8190 12727 8191 12753
rect 8191 12727 8217 12753
rect 8217 12727 8218 12753
rect 8190 12726 8218 12727
rect 8246 12670 8274 12698
rect 8078 12305 8106 12306
rect 8078 12279 8079 12305
rect 8079 12279 8105 12305
rect 8105 12279 8106 12305
rect 8078 12278 8106 12279
rect 2238 12165 2266 12166
rect 2238 12139 2239 12165
rect 2239 12139 2265 12165
rect 2265 12139 2266 12165
rect 2238 12138 2266 12139
rect 2290 12165 2318 12166
rect 2290 12139 2291 12165
rect 2291 12139 2317 12165
rect 2317 12139 2318 12165
rect 2290 12138 2318 12139
rect 2342 12165 2370 12166
rect 2342 12139 2343 12165
rect 2343 12139 2369 12165
rect 2369 12139 2370 12165
rect 2342 12138 2370 12139
rect 2142 11969 2170 11970
rect 2142 11943 2143 11969
rect 2143 11943 2169 11969
rect 2169 11943 2170 11969
rect 2142 11942 2170 11943
rect 6734 11942 6762 11970
rect 7798 11913 7826 11914
rect 7798 11887 7799 11913
rect 7799 11887 7825 11913
rect 7825 11887 7826 11913
rect 7798 11886 7826 11887
rect 5894 11633 5922 11634
rect 5894 11607 5895 11633
rect 5895 11607 5921 11633
rect 5921 11607 5922 11633
rect 5894 11606 5922 11607
rect 2238 11381 2266 11382
rect 2238 11355 2239 11381
rect 2239 11355 2265 11381
rect 2265 11355 2266 11381
rect 2238 11354 2266 11355
rect 2290 11381 2318 11382
rect 2290 11355 2291 11381
rect 2291 11355 2317 11381
rect 2317 11355 2318 11381
rect 2290 11354 2318 11355
rect 2342 11381 2370 11382
rect 2342 11355 2343 11381
rect 2343 11355 2369 11381
rect 2369 11355 2370 11381
rect 2342 11354 2370 11355
rect 7182 11577 7210 11578
rect 7182 11551 7183 11577
rect 7183 11551 7209 11577
rect 7209 11551 7210 11577
rect 7182 11550 7210 11551
rect 7406 11550 7434 11578
rect 6958 11521 6986 11522
rect 6958 11495 6959 11521
rect 6959 11495 6985 11521
rect 6985 11495 6986 11521
rect 6958 11494 6986 11495
rect 5558 10934 5586 10962
rect 5838 10934 5866 10962
rect 2086 10766 2114 10794
rect 7462 10934 7490 10962
rect 7238 10878 7266 10906
rect 6174 10737 6202 10738
rect 6174 10711 6175 10737
rect 6175 10711 6201 10737
rect 6201 10711 6202 10737
rect 6174 10710 6202 10711
rect 6846 10710 6874 10738
rect 2238 10597 2266 10598
rect 2238 10571 2239 10597
rect 2239 10571 2265 10597
rect 2265 10571 2266 10597
rect 2238 10570 2266 10571
rect 2290 10597 2318 10598
rect 2290 10571 2291 10597
rect 2291 10571 2317 10597
rect 2317 10571 2318 10597
rect 2290 10570 2318 10571
rect 2342 10597 2370 10598
rect 2342 10571 2343 10597
rect 2343 10571 2369 10597
rect 2369 10571 2370 10597
rect 2342 10570 2370 10571
rect 7518 11494 7546 11522
rect 7742 10878 7770 10906
rect 7854 11158 7882 11186
rect 7686 10822 7714 10850
rect 2142 10009 2170 10010
rect 2142 9983 2143 10009
rect 2143 9983 2169 10009
rect 2169 9983 2170 10009
rect 2142 9982 2170 9983
rect 4998 9982 5026 10010
rect 966 9897 994 9898
rect 966 9871 967 9897
rect 967 9871 993 9897
rect 993 9871 994 9897
rect 966 9870 994 9871
rect 2238 9813 2266 9814
rect 2238 9787 2239 9813
rect 2239 9787 2265 9813
rect 2265 9787 2266 9813
rect 2238 9786 2266 9787
rect 2290 9813 2318 9814
rect 2290 9787 2291 9813
rect 2291 9787 2317 9813
rect 2317 9787 2318 9813
rect 2290 9786 2318 9787
rect 2342 9813 2370 9814
rect 2342 9787 2343 9813
rect 2343 9787 2369 9813
rect 2369 9787 2370 9813
rect 2342 9786 2370 9787
rect 6062 9926 6090 9954
rect 6454 9617 6482 9618
rect 6454 9591 6455 9617
rect 6455 9591 6481 9617
rect 6481 9591 6482 9617
rect 6454 9590 6482 9591
rect 6790 9590 6818 9618
rect 4998 9534 5026 9562
rect 7126 10038 7154 10066
rect 7070 10009 7098 10010
rect 7070 9983 7071 10009
rect 7071 9983 7097 10009
rect 7097 9983 7098 10009
rect 7070 9982 7098 9983
rect 7014 9953 7042 9954
rect 7014 9927 7015 9953
rect 7015 9927 7041 9953
rect 7041 9927 7042 9953
rect 7014 9926 7042 9927
rect 7182 9870 7210 9898
rect 7238 9982 7266 10010
rect 6510 9310 6538 9338
rect 2238 9029 2266 9030
rect 2238 9003 2239 9029
rect 2239 9003 2265 9029
rect 2265 9003 2266 9029
rect 2238 9002 2266 9003
rect 2290 9029 2318 9030
rect 2290 9003 2291 9029
rect 2291 9003 2317 9029
rect 2317 9003 2318 9029
rect 2290 9002 2318 9003
rect 2342 9029 2370 9030
rect 2342 9003 2343 9029
rect 2343 9003 2369 9029
rect 2369 9003 2370 9029
rect 2342 9002 2370 9003
rect 966 8889 994 8890
rect 966 8863 967 8889
rect 967 8863 993 8889
rect 993 8863 994 8889
rect 966 8862 994 8863
rect 2142 8833 2170 8834
rect 2142 8807 2143 8833
rect 2143 8807 2169 8833
rect 2169 8807 2170 8833
rect 2142 8806 2170 8807
rect 6902 9142 6930 9170
rect 6790 8945 6818 8946
rect 6790 8919 6791 8945
rect 6791 8919 6817 8945
rect 6817 8919 6818 8945
rect 6790 8918 6818 8919
rect 5390 8750 5418 8778
rect 966 8414 994 8442
rect 2142 8441 2170 8442
rect 2142 8415 2143 8441
rect 2143 8415 2169 8441
rect 2169 8415 2170 8441
rect 2142 8414 2170 8415
rect 5390 8414 5418 8442
rect 5446 8806 5474 8834
rect 6734 8806 6762 8834
rect 6846 8833 6874 8834
rect 6846 8807 6847 8833
rect 6847 8807 6873 8833
rect 6873 8807 6874 8833
rect 6846 8806 6874 8807
rect 7294 9561 7322 9562
rect 7294 9535 7295 9561
rect 7295 9535 7321 9561
rect 7321 9535 7322 9561
rect 7294 9534 7322 9535
rect 7238 9337 7266 9338
rect 7238 9311 7239 9337
rect 7239 9311 7265 9337
rect 7265 9311 7266 9337
rect 7238 9310 7266 9311
rect 7294 9254 7322 9282
rect 7238 9225 7266 9226
rect 7238 9199 7239 9225
rect 7239 9199 7265 9225
rect 7265 9199 7266 9225
rect 7238 9198 7266 9199
rect 7126 8918 7154 8946
rect 7238 8862 7266 8890
rect 7406 9030 7434 9058
rect 7686 10038 7714 10066
rect 7686 9926 7714 9954
rect 8078 11942 8106 11970
rect 8134 11830 8162 11858
rect 7910 9870 7938 9898
rect 8806 12670 8834 12698
rect 9142 13118 9170 13146
rect 8806 12305 8834 12306
rect 8806 12279 8807 12305
rect 8807 12279 8833 12305
rect 8833 12279 8834 12305
rect 8806 12278 8834 12279
rect 8414 12110 8442 12138
rect 9030 12110 9058 12138
rect 8862 12081 8890 12082
rect 8862 12055 8863 12081
rect 8863 12055 8889 12081
rect 8889 12055 8890 12081
rect 8862 12054 8890 12055
rect 8470 11913 8498 11914
rect 8470 11887 8471 11913
rect 8471 11887 8497 11913
rect 8497 11887 8498 11913
rect 8470 11886 8498 11887
rect 8414 11857 8442 11858
rect 8414 11831 8415 11857
rect 8415 11831 8441 11857
rect 8441 11831 8442 11857
rect 8414 11830 8442 11831
rect 8526 11857 8554 11858
rect 8526 11831 8527 11857
rect 8527 11831 8553 11857
rect 8553 11831 8554 11857
rect 8526 11830 8554 11831
rect 8246 11718 8274 11746
rect 8414 11606 8442 11634
rect 8190 11550 8218 11578
rect 8358 11577 8386 11578
rect 8358 11551 8359 11577
rect 8359 11551 8385 11577
rect 8385 11551 8386 11577
rect 8358 11550 8386 11551
rect 8582 11606 8610 11634
rect 8750 11886 8778 11914
rect 8918 11830 8946 11858
rect 8414 10934 8442 10962
rect 8862 11718 8890 11746
rect 8246 10878 8274 10906
rect 8302 10822 8330 10850
rect 8414 10318 8442 10346
rect 7966 9982 7994 10010
rect 8582 10934 8610 10962
rect 8694 10849 8722 10850
rect 8694 10823 8695 10849
rect 8695 10823 8721 10849
rect 8721 10823 8722 10849
rect 8694 10822 8722 10823
rect 8806 10878 8834 10906
rect 8022 9646 8050 9674
rect 8302 9646 8330 9674
rect 7630 9086 7658 9114
rect 7742 9169 7770 9170
rect 7742 9143 7743 9169
rect 7743 9143 7769 9169
rect 7769 9143 7770 9169
rect 7742 9142 7770 9143
rect 7406 8806 7434 8834
rect 7574 8777 7602 8778
rect 7574 8751 7575 8777
rect 7575 8751 7601 8777
rect 7601 8751 7602 8777
rect 7574 8750 7602 8751
rect 6510 8694 6538 8722
rect 7406 8721 7434 8722
rect 7406 8695 7407 8721
rect 7407 8695 7433 8721
rect 7433 8695 7434 8721
rect 7406 8694 7434 8695
rect 7126 8638 7154 8666
rect 7742 8638 7770 8666
rect 8246 9422 8274 9450
rect 8134 9254 8162 9282
rect 7854 9086 7882 9114
rect 8470 9758 8498 9786
rect 8694 9673 8722 9674
rect 8694 9647 8695 9673
rect 8695 9647 8721 9673
rect 8721 9647 8722 9673
rect 8694 9646 8722 9647
rect 8582 9617 8610 9618
rect 8582 9591 8583 9617
rect 8583 9591 8609 9617
rect 8609 9591 8610 9617
rect 8582 9590 8610 9591
rect 8750 9310 8778 9338
rect 8974 11633 9002 11634
rect 8974 11607 8975 11633
rect 8975 11607 9001 11633
rect 9001 11607 9002 11633
rect 8974 11606 9002 11607
rect 10654 13481 10682 13482
rect 10654 13455 10655 13481
rect 10655 13455 10681 13481
rect 10681 13455 10682 13481
rect 10654 13454 10682 13455
rect 10934 14238 10962 14266
rect 9918 13341 9946 13342
rect 9918 13315 9919 13341
rect 9919 13315 9945 13341
rect 9945 13315 9946 13341
rect 9918 13314 9946 13315
rect 9970 13341 9998 13342
rect 9970 13315 9971 13341
rect 9971 13315 9997 13341
rect 9997 13315 9998 13341
rect 9970 13314 9998 13315
rect 10022 13341 10050 13342
rect 10022 13315 10023 13341
rect 10023 13315 10049 13341
rect 10049 13315 10050 13341
rect 10022 13314 10050 13315
rect 9926 13201 9954 13202
rect 9926 13175 9927 13201
rect 9927 13175 9953 13201
rect 9953 13175 9954 13201
rect 9926 13174 9954 13175
rect 9870 13145 9898 13146
rect 9870 13119 9871 13145
rect 9871 13119 9897 13145
rect 9897 13119 9898 13145
rect 9870 13118 9898 13119
rect 10206 12697 10234 12698
rect 10206 12671 10207 12697
rect 10207 12671 10233 12697
rect 10233 12671 10234 12697
rect 10206 12670 10234 12671
rect 9918 12557 9946 12558
rect 9918 12531 9919 12557
rect 9919 12531 9945 12557
rect 9945 12531 9946 12557
rect 9918 12530 9946 12531
rect 9970 12557 9998 12558
rect 9970 12531 9971 12557
rect 9971 12531 9997 12557
rect 9997 12531 9998 12557
rect 9970 12530 9998 12531
rect 10022 12557 10050 12558
rect 10022 12531 10023 12557
rect 10023 12531 10049 12557
rect 10049 12531 10050 12557
rect 10022 12530 10050 12531
rect 9478 12054 9506 12082
rect 9142 11886 9170 11914
rect 9422 11886 9450 11914
rect 9086 11718 9114 11746
rect 8918 11438 8946 11466
rect 8918 11185 8946 11186
rect 8918 11159 8919 11185
rect 8919 11159 8945 11185
rect 8945 11159 8946 11185
rect 8918 11158 8946 11159
rect 8862 10345 8890 10346
rect 8862 10319 8863 10345
rect 8863 10319 8889 10345
rect 8889 10319 8890 10345
rect 8862 10318 8890 10319
rect 8862 9702 8890 9730
rect 9086 11073 9114 11074
rect 9086 11047 9087 11073
rect 9087 11047 9113 11073
rect 9113 11047 9114 11073
rect 9086 11046 9114 11047
rect 9254 11577 9282 11578
rect 9254 11551 9255 11577
rect 9255 11551 9281 11577
rect 9281 11551 9282 11577
rect 9254 11550 9282 11551
rect 8974 10681 9002 10682
rect 8974 10655 8975 10681
rect 8975 10655 9001 10681
rect 9001 10655 9002 10681
rect 8974 10654 9002 10655
rect 8918 9590 8946 9618
rect 9310 10094 9338 10122
rect 9422 11606 9450 11634
rect 9646 11521 9674 11522
rect 9646 11495 9647 11521
rect 9647 11495 9673 11521
rect 9673 11495 9674 11521
rect 9646 11494 9674 11495
rect 9422 11214 9450 11242
rect 9758 11073 9786 11074
rect 9758 11047 9759 11073
rect 9759 11047 9785 11073
rect 9785 11047 9786 11073
rect 9758 11046 9786 11047
rect 9478 10878 9506 10906
rect 9478 10793 9506 10794
rect 9478 10767 9479 10793
rect 9479 10767 9505 10793
rect 9505 10767 9506 10793
rect 9478 10766 9506 10767
rect 9702 10793 9730 10794
rect 9702 10767 9703 10793
rect 9703 10767 9729 10793
rect 9729 10767 9730 10793
rect 9702 10766 9730 10767
rect 10654 13257 10682 13258
rect 10654 13231 10655 13257
rect 10655 13231 10681 13257
rect 10681 13231 10682 13257
rect 10654 13230 10682 13231
rect 10542 13201 10570 13202
rect 10542 13175 10543 13201
rect 10543 13175 10569 13201
rect 10569 13175 10570 13201
rect 10542 13174 10570 13175
rect 10710 13145 10738 13146
rect 10710 13119 10711 13145
rect 10711 13119 10737 13145
rect 10737 13119 10738 13145
rect 10710 13118 10738 13119
rect 11046 14657 11074 14658
rect 11046 14631 11047 14657
rect 11047 14631 11073 14657
rect 11073 14631 11074 14657
rect 11046 14630 11074 14631
rect 11214 14238 11242 14266
rect 10990 13230 11018 13258
rect 12334 13174 12362 13202
rect 10934 12726 10962 12754
rect 10486 11998 10514 12026
rect 9982 11913 10010 11914
rect 9982 11887 9983 11913
rect 9983 11887 10009 11913
rect 10009 11887 10010 11913
rect 9982 11886 10010 11887
rect 9918 11773 9946 11774
rect 9918 11747 9919 11773
rect 9919 11747 9945 11773
rect 9945 11747 9946 11773
rect 9918 11746 9946 11747
rect 9970 11773 9998 11774
rect 9970 11747 9971 11773
rect 9971 11747 9997 11773
rect 9997 11747 9998 11773
rect 9970 11746 9998 11747
rect 10022 11773 10050 11774
rect 10022 11747 10023 11773
rect 10023 11747 10049 11773
rect 10049 11747 10050 11773
rect 10022 11746 10050 11747
rect 10486 11550 10514 11578
rect 9926 11158 9954 11186
rect 10318 11214 10346 11242
rect 10150 11129 10178 11130
rect 10150 11103 10151 11129
rect 10151 11103 10177 11129
rect 10177 11103 10178 11129
rect 10150 11102 10178 11103
rect 10094 11073 10122 11074
rect 10094 11047 10095 11073
rect 10095 11047 10121 11073
rect 10121 11047 10122 11073
rect 10094 11046 10122 11047
rect 9918 10989 9946 10990
rect 9918 10963 9919 10989
rect 9919 10963 9945 10989
rect 9945 10963 9946 10989
rect 9918 10962 9946 10963
rect 9970 10989 9998 10990
rect 9970 10963 9971 10989
rect 9971 10963 9997 10989
rect 9997 10963 9998 10989
rect 9970 10962 9998 10963
rect 10022 10989 10050 10990
rect 10022 10963 10023 10989
rect 10023 10963 10049 10989
rect 10049 10963 10050 10989
rect 10022 10962 10050 10963
rect 9702 10486 9730 10514
rect 9926 10878 9954 10906
rect 9366 9926 9394 9954
rect 9030 9617 9058 9618
rect 9030 9591 9031 9617
rect 9031 9591 9057 9617
rect 9057 9591 9058 9617
rect 9030 9590 9058 9591
rect 8862 9561 8890 9562
rect 8862 9535 8863 9561
rect 8863 9535 8889 9561
rect 8889 9535 8890 9561
rect 8862 9534 8890 9535
rect 9030 9478 9058 9506
rect 8358 9086 8386 9114
rect 8862 9198 8890 9226
rect 8414 8889 8442 8890
rect 8414 8863 8415 8889
rect 8415 8863 8441 8889
rect 8441 8863 8442 8889
rect 8414 8862 8442 8863
rect 8974 9225 9002 9226
rect 8974 9199 8975 9225
rect 8975 9199 9001 9225
rect 9001 9199 9002 9225
rect 8974 9198 9002 9199
rect 9086 9422 9114 9450
rect 9142 9758 9170 9786
rect 9310 9561 9338 9562
rect 9310 9535 9311 9561
rect 9311 9535 9337 9561
rect 9337 9535 9338 9561
rect 9310 9534 9338 9535
rect 9478 9254 9506 9282
rect 9254 9198 9282 9226
rect 9198 9169 9226 9170
rect 9198 9143 9199 9169
rect 9199 9143 9225 9169
rect 9225 9143 9226 9169
rect 9198 9142 9226 9143
rect 9030 8862 9058 8890
rect 9198 8862 9226 8890
rect 8806 8833 8834 8834
rect 8806 8807 8807 8833
rect 8807 8807 8833 8833
rect 8833 8807 8834 8833
rect 8806 8806 8834 8807
rect 8526 8721 8554 8722
rect 8526 8695 8527 8721
rect 8527 8695 8553 8721
rect 8553 8695 8554 8721
rect 8526 8694 8554 8695
rect 8414 8526 8442 8554
rect 2238 8245 2266 8246
rect 2238 8219 2239 8245
rect 2239 8219 2265 8245
rect 2265 8219 2266 8245
rect 2238 8218 2266 8219
rect 2290 8245 2318 8246
rect 2290 8219 2291 8245
rect 2291 8219 2317 8245
rect 2317 8219 2318 8245
rect 2290 8218 2318 8219
rect 2342 8245 2370 8246
rect 2342 8219 2343 8245
rect 2343 8219 2369 8245
rect 2369 8219 2370 8245
rect 2342 8218 2370 8219
rect 7350 8358 7378 8386
rect 7798 8385 7826 8386
rect 7798 8359 7799 8385
rect 7799 8359 7825 8385
rect 7825 8359 7826 8385
rect 7798 8358 7826 8359
rect 8078 8134 8106 8162
rect 8414 8134 8442 8162
rect 7070 7574 7098 7602
rect 2238 7461 2266 7462
rect 2238 7435 2239 7461
rect 2239 7435 2265 7461
rect 2265 7435 2266 7461
rect 2238 7434 2266 7435
rect 2290 7461 2318 7462
rect 2290 7435 2291 7461
rect 2291 7435 2317 7461
rect 2317 7435 2318 7461
rect 2290 7434 2318 7435
rect 2342 7461 2370 7462
rect 2342 7435 2343 7461
rect 2343 7435 2369 7461
rect 2369 7435 2370 7461
rect 2342 7434 2370 7435
rect 8134 7126 8162 7154
rect 2238 6677 2266 6678
rect 2238 6651 2239 6677
rect 2239 6651 2265 6677
rect 2265 6651 2266 6677
rect 2238 6650 2266 6651
rect 2290 6677 2318 6678
rect 2290 6651 2291 6677
rect 2291 6651 2317 6677
rect 2317 6651 2318 6677
rect 2290 6650 2318 6651
rect 2342 6677 2370 6678
rect 2342 6651 2343 6677
rect 2343 6651 2369 6677
rect 2369 6651 2370 6677
rect 2342 6650 2370 6651
rect 7798 6481 7826 6482
rect 7798 6455 7799 6481
rect 7799 6455 7825 6481
rect 7825 6455 7826 6481
rect 7798 6454 7826 6455
rect 2238 5893 2266 5894
rect 2238 5867 2239 5893
rect 2239 5867 2265 5893
rect 2265 5867 2266 5893
rect 2238 5866 2266 5867
rect 2290 5893 2318 5894
rect 2290 5867 2291 5893
rect 2291 5867 2317 5893
rect 2317 5867 2318 5893
rect 2290 5866 2318 5867
rect 2342 5893 2370 5894
rect 2342 5867 2343 5893
rect 2343 5867 2369 5893
rect 2369 5867 2370 5893
rect 2342 5866 2370 5867
rect 2238 5109 2266 5110
rect 2238 5083 2239 5109
rect 2239 5083 2265 5109
rect 2265 5083 2266 5109
rect 2238 5082 2266 5083
rect 2290 5109 2318 5110
rect 2290 5083 2291 5109
rect 2291 5083 2317 5109
rect 2317 5083 2318 5109
rect 2290 5082 2318 5083
rect 2342 5109 2370 5110
rect 2342 5083 2343 5109
rect 2343 5083 2369 5109
rect 2369 5083 2370 5109
rect 2342 5082 2370 5083
rect 2238 4325 2266 4326
rect 2238 4299 2239 4325
rect 2239 4299 2265 4325
rect 2265 4299 2266 4325
rect 2238 4298 2266 4299
rect 2290 4325 2318 4326
rect 2290 4299 2291 4325
rect 2291 4299 2317 4325
rect 2317 4299 2318 4325
rect 2290 4298 2318 4299
rect 2342 4325 2370 4326
rect 2342 4299 2343 4325
rect 2343 4299 2369 4325
rect 2369 4299 2370 4325
rect 2342 4298 2370 4299
rect 9086 8582 9114 8610
rect 8862 8441 8890 8442
rect 8862 8415 8863 8441
rect 8863 8415 8889 8441
rect 8889 8415 8890 8441
rect 8862 8414 8890 8415
rect 8974 8385 9002 8386
rect 8974 8359 8975 8385
rect 8975 8359 9001 8385
rect 9001 8359 9002 8385
rect 8974 8358 9002 8359
rect 8750 7574 8778 7602
rect 9366 9030 9394 9058
rect 9310 8750 9338 8778
rect 9926 10401 9954 10402
rect 9926 10375 9927 10401
rect 9927 10375 9953 10401
rect 9953 10375 9954 10401
rect 9926 10374 9954 10375
rect 10206 10430 10234 10458
rect 9918 10205 9946 10206
rect 9918 10179 9919 10205
rect 9919 10179 9945 10205
rect 9945 10179 9946 10205
rect 9918 10178 9946 10179
rect 9970 10205 9998 10206
rect 9970 10179 9971 10205
rect 9971 10179 9997 10205
rect 9997 10179 9998 10205
rect 9970 10178 9998 10179
rect 10022 10205 10050 10206
rect 10022 10179 10023 10205
rect 10023 10179 10049 10205
rect 10049 10179 10050 10205
rect 10022 10178 10050 10179
rect 9814 9758 9842 9786
rect 9870 10038 9898 10066
rect 9758 9729 9786 9730
rect 9758 9703 9759 9729
rect 9759 9703 9785 9729
rect 9785 9703 9786 9729
rect 9758 9702 9786 9703
rect 9814 9505 9842 9506
rect 9814 9479 9815 9505
rect 9815 9479 9841 9505
rect 9841 9479 9842 9505
rect 9814 9478 9842 9479
rect 10710 10374 10738 10402
rect 10262 10065 10290 10066
rect 10262 10039 10263 10065
rect 10263 10039 10289 10065
rect 10289 10039 10290 10065
rect 10262 10038 10290 10039
rect 10094 9982 10122 10010
rect 10710 9982 10738 10010
rect 10038 9534 10066 9562
rect 9918 9421 9946 9422
rect 9918 9395 9919 9421
rect 9919 9395 9945 9421
rect 9945 9395 9946 9421
rect 9918 9394 9946 9395
rect 9970 9421 9998 9422
rect 9970 9395 9971 9421
rect 9971 9395 9997 9421
rect 9997 9395 9998 9421
rect 9970 9394 9998 9395
rect 10022 9421 10050 9422
rect 10022 9395 10023 9421
rect 10023 9395 10049 9421
rect 10049 9395 10050 9421
rect 10022 9394 10050 9395
rect 9926 9281 9954 9282
rect 9926 9255 9927 9281
rect 9927 9255 9953 9281
rect 9953 9255 9954 9281
rect 9926 9254 9954 9255
rect 9254 8694 9282 8722
rect 9254 8414 9282 8442
rect 9422 8358 9450 8386
rect 10990 13118 11018 13146
rect 11270 13089 11298 13090
rect 11270 13063 11271 13089
rect 11271 13063 11297 13089
rect 11297 13063 11298 13089
rect 11270 13062 11298 13063
rect 11774 13062 11802 13090
rect 17598 18437 17626 18438
rect 17598 18411 17599 18437
rect 17599 18411 17625 18437
rect 17625 18411 17626 18437
rect 17598 18410 17626 18411
rect 17650 18437 17678 18438
rect 17650 18411 17651 18437
rect 17651 18411 17677 18437
rect 17677 18411 17678 18437
rect 17650 18410 17678 18411
rect 17702 18437 17730 18438
rect 17702 18411 17703 18437
rect 17703 18411 17729 18437
rect 17729 18411 17730 18437
rect 17702 18410 17730 18411
rect 17598 17653 17626 17654
rect 17598 17627 17599 17653
rect 17599 17627 17625 17653
rect 17625 17627 17626 17653
rect 17598 17626 17626 17627
rect 17650 17653 17678 17654
rect 17650 17627 17651 17653
rect 17651 17627 17677 17653
rect 17677 17627 17678 17653
rect 17650 17626 17678 17627
rect 17702 17653 17730 17654
rect 17702 17627 17703 17653
rect 17703 17627 17729 17653
rect 17729 17627 17730 17653
rect 17702 17626 17730 17627
rect 17598 16869 17626 16870
rect 17598 16843 17599 16869
rect 17599 16843 17625 16869
rect 17625 16843 17626 16869
rect 17598 16842 17626 16843
rect 17650 16869 17678 16870
rect 17650 16843 17651 16869
rect 17651 16843 17677 16869
rect 17677 16843 17678 16869
rect 17650 16842 17678 16843
rect 17702 16869 17730 16870
rect 17702 16843 17703 16869
rect 17703 16843 17729 16869
rect 17729 16843 17730 16869
rect 17702 16842 17730 16843
rect 17598 16085 17626 16086
rect 17598 16059 17599 16085
rect 17599 16059 17625 16085
rect 17625 16059 17626 16085
rect 17598 16058 17626 16059
rect 17650 16085 17678 16086
rect 17650 16059 17651 16085
rect 17651 16059 17677 16085
rect 17677 16059 17678 16085
rect 17650 16058 17678 16059
rect 17702 16085 17730 16086
rect 17702 16059 17703 16085
rect 17703 16059 17729 16085
rect 17729 16059 17730 16085
rect 17702 16058 17730 16059
rect 17598 15301 17626 15302
rect 17598 15275 17599 15301
rect 17599 15275 17625 15301
rect 17625 15275 17626 15301
rect 17598 15274 17626 15275
rect 17650 15301 17678 15302
rect 17650 15275 17651 15301
rect 17651 15275 17677 15301
rect 17677 15275 17678 15301
rect 17650 15274 17678 15275
rect 17702 15301 17730 15302
rect 17702 15275 17703 15301
rect 17703 15275 17729 15301
rect 17729 15275 17730 15301
rect 17702 15274 17730 15275
rect 17598 14517 17626 14518
rect 17598 14491 17599 14517
rect 17599 14491 17625 14517
rect 17625 14491 17626 14517
rect 17598 14490 17626 14491
rect 17650 14517 17678 14518
rect 17650 14491 17651 14517
rect 17651 14491 17677 14517
rect 17677 14491 17678 14517
rect 17650 14490 17678 14491
rect 17702 14517 17730 14518
rect 17702 14491 17703 14517
rect 17703 14491 17729 14517
rect 17729 14491 17730 14517
rect 17702 14490 17730 14491
rect 17598 13733 17626 13734
rect 17598 13707 17599 13733
rect 17599 13707 17625 13733
rect 17625 13707 17626 13733
rect 17598 13706 17626 13707
rect 17650 13733 17678 13734
rect 17650 13707 17651 13733
rect 17651 13707 17677 13733
rect 17677 13707 17678 13733
rect 17650 13706 17678 13707
rect 17702 13733 17730 13734
rect 17702 13707 17703 13733
rect 17703 13707 17729 13733
rect 17729 13707 17730 13733
rect 17702 13706 17730 13707
rect 12670 13201 12698 13202
rect 12670 13175 12671 13201
rect 12671 13175 12697 13201
rect 12697 13175 12698 13201
rect 12670 13174 12698 13175
rect 12726 13145 12754 13146
rect 12726 13119 12727 13145
rect 12727 13119 12753 13145
rect 12753 13119 12754 13145
rect 12726 13118 12754 13119
rect 13510 13145 13538 13146
rect 13510 13119 13511 13145
rect 13511 13119 13537 13145
rect 13537 13119 13538 13145
rect 13510 13118 13538 13119
rect 12054 13006 12082 13034
rect 12670 13033 12698 13034
rect 12670 13007 12671 13033
rect 12671 13007 12697 13033
rect 12697 13007 12698 13033
rect 12670 13006 12698 13007
rect 12446 12753 12474 12754
rect 12446 12727 12447 12753
rect 12447 12727 12473 12753
rect 12473 12727 12474 12753
rect 12446 12726 12474 12727
rect 12670 12753 12698 12754
rect 12670 12727 12671 12753
rect 12671 12727 12697 12753
rect 12697 12727 12698 12753
rect 12670 12726 12698 12727
rect 10822 12025 10850 12026
rect 10822 11999 10823 12025
rect 10823 11999 10849 12025
rect 10849 11999 10850 12025
rect 10822 11998 10850 11999
rect 11830 12054 11858 12082
rect 12950 12726 12978 12754
rect 13174 13006 13202 13034
rect 10878 11494 10906 11522
rect 11214 11214 11242 11242
rect 10934 11185 10962 11186
rect 10934 11159 10935 11185
rect 10935 11159 10961 11185
rect 10961 11159 10962 11185
rect 10934 11158 10962 11159
rect 11438 11185 11466 11186
rect 11438 11159 11439 11185
rect 11439 11159 11465 11185
rect 11465 11159 11466 11185
rect 11438 11158 11466 11159
rect 11606 11185 11634 11186
rect 11606 11159 11607 11185
rect 11607 11159 11633 11185
rect 11633 11159 11634 11185
rect 11606 11158 11634 11159
rect 11158 10934 11186 10962
rect 11718 10934 11746 10962
rect 12670 11774 12698 11802
rect 11886 11214 11914 11242
rect 11830 11046 11858 11074
rect 10934 10486 10962 10514
rect 11382 10457 11410 10458
rect 11382 10431 11383 10457
rect 11383 10431 11409 10457
rect 11409 10431 11410 10457
rect 11382 10430 11410 10431
rect 11662 10430 11690 10458
rect 11102 10401 11130 10402
rect 11102 10375 11103 10401
rect 11103 10375 11129 10401
rect 11129 10375 11130 10401
rect 11102 10374 11130 10375
rect 10822 10038 10850 10066
rect 11382 10094 11410 10122
rect 11886 10654 11914 10682
rect 11942 10374 11970 10402
rect 11046 10009 11074 10010
rect 11046 9983 11047 10009
rect 11047 9983 11073 10009
rect 11073 9983 11074 10009
rect 11046 9982 11074 9983
rect 10878 9870 10906 9898
rect 11606 10009 11634 10010
rect 11606 9983 11607 10009
rect 11607 9983 11633 10009
rect 11633 9983 11634 10009
rect 11606 9982 11634 9983
rect 11214 9590 11242 9618
rect 10822 9478 10850 9506
rect 10094 9142 10122 9170
rect 9702 8694 9730 8722
rect 9918 8637 9946 8638
rect 9918 8611 9919 8637
rect 9919 8611 9945 8637
rect 9945 8611 9946 8637
rect 9918 8610 9946 8611
rect 9970 8637 9998 8638
rect 9970 8611 9971 8637
rect 9971 8611 9997 8637
rect 9997 8611 9998 8637
rect 9970 8610 9998 8611
rect 10022 8637 10050 8638
rect 10022 8611 10023 8637
rect 10023 8611 10049 8637
rect 10049 8611 10050 8637
rect 10022 8610 10050 8611
rect 10822 9225 10850 9226
rect 10822 9199 10823 9225
rect 10823 9199 10849 9225
rect 10849 9199 10850 9225
rect 10822 9198 10850 9199
rect 11158 9505 11186 9506
rect 11158 9479 11159 9505
rect 11159 9479 11185 9505
rect 11185 9479 11186 9505
rect 11158 9478 11186 9479
rect 11102 9310 11130 9338
rect 10990 9142 11018 9170
rect 10934 9086 10962 9114
rect 10822 8694 10850 8722
rect 10766 8414 10794 8442
rect 10710 8161 10738 8162
rect 10710 8135 10711 8161
rect 10711 8135 10737 8161
rect 10737 8135 10738 8161
rect 10710 8134 10738 8135
rect 10990 8638 11018 8666
rect 10654 8078 10682 8106
rect 9478 7937 9506 7938
rect 9478 7911 9479 7937
rect 9479 7911 9505 7937
rect 9505 7911 9506 7937
rect 9478 7910 9506 7911
rect 10150 7910 10178 7938
rect 9918 7853 9946 7854
rect 9918 7827 9919 7853
rect 9919 7827 9945 7853
rect 9945 7827 9946 7853
rect 9918 7826 9946 7827
rect 9970 7853 9998 7854
rect 9970 7827 9971 7853
rect 9971 7827 9997 7853
rect 9997 7827 9998 7853
rect 9970 7826 9998 7827
rect 10022 7853 10050 7854
rect 10022 7827 10023 7853
rect 10023 7827 10049 7853
rect 10049 7827 10050 7853
rect 10022 7826 10050 7827
rect 10094 7574 10122 7602
rect 8582 7153 8610 7154
rect 8582 7127 8583 7153
rect 8583 7127 8609 7153
rect 8609 7127 8610 7153
rect 8582 7126 8610 7127
rect 9918 7069 9946 7070
rect 9918 7043 9919 7069
rect 9919 7043 9945 7069
rect 9945 7043 9946 7069
rect 9918 7042 9946 7043
rect 9970 7069 9998 7070
rect 9970 7043 9971 7069
rect 9971 7043 9997 7069
rect 9997 7043 9998 7069
rect 9970 7042 9998 7043
rect 10022 7069 10050 7070
rect 10022 7043 10023 7069
rect 10023 7043 10049 7069
rect 10049 7043 10050 7069
rect 10022 7042 10050 7043
rect 10094 6510 10122 6538
rect 9478 6481 9506 6482
rect 9478 6455 9479 6481
rect 9479 6455 9505 6481
rect 9505 6455 9506 6481
rect 9478 6454 9506 6455
rect 9918 6285 9946 6286
rect 9918 6259 9919 6285
rect 9919 6259 9945 6285
rect 9945 6259 9946 6285
rect 9918 6258 9946 6259
rect 9970 6285 9998 6286
rect 9970 6259 9971 6285
rect 9971 6259 9997 6285
rect 9997 6259 9998 6285
rect 9970 6258 9998 6259
rect 10022 6285 10050 6286
rect 10022 6259 10023 6285
rect 10023 6259 10049 6285
rect 10049 6259 10050 6285
rect 10022 6258 10050 6259
rect 9918 5501 9946 5502
rect 9918 5475 9919 5501
rect 9919 5475 9945 5501
rect 9945 5475 9946 5501
rect 9918 5474 9946 5475
rect 9970 5501 9998 5502
rect 9970 5475 9971 5501
rect 9971 5475 9997 5501
rect 9997 5475 9998 5501
rect 9970 5474 9998 5475
rect 10022 5501 10050 5502
rect 10022 5475 10023 5501
rect 10023 5475 10049 5501
rect 10049 5475 10050 5501
rect 10022 5474 10050 5475
rect 9918 4717 9946 4718
rect 9918 4691 9919 4717
rect 9919 4691 9945 4717
rect 9945 4691 9946 4717
rect 9918 4690 9946 4691
rect 9970 4717 9998 4718
rect 9970 4691 9971 4717
rect 9971 4691 9997 4717
rect 9997 4691 9998 4717
rect 9970 4690 9998 4691
rect 10022 4717 10050 4718
rect 10022 4691 10023 4717
rect 10023 4691 10049 4717
rect 10049 4691 10050 4717
rect 10022 4690 10050 4691
rect 2238 3541 2266 3542
rect 2238 3515 2239 3541
rect 2239 3515 2265 3541
rect 2265 3515 2266 3541
rect 2238 3514 2266 3515
rect 2290 3541 2318 3542
rect 2290 3515 2291 3541
rect 2291 3515 2317 3541
rect 2317 3515 2318 3541
rect 2290 3514 2318 3515
rect 2342 3541 2370 3542
rect 2342 3515 2343 3541
rect 2343 3515 2369 3541
rect 2369 3515 2370 3541
rect 2342 3514 2370 3515
rect 2238 2757 2266 2758
rect 2238 2731 2239 2757
rect 2239 2731 2265 2757
rect 2265 2731 2266 2757
rect 2238 2730 2266 2731
rect 2290 2757 2318 2758
rect 2290 2731 2291 2757
rect 2291 2731 2317 2757
rect 2317 2731 2318 2757
rect 2290 2730 2318 2731
rect 2342 2757 2370 2758
rect 2342 2731 2343 2757
rect 2343 2731 2369 2757
rect 2369 2731 2370 2757
rect 2342 2730 2370 2731
rect 10374 7601 10402 7602
rect 10374 7575 10375 7601
rect 10375 7575 10401 7601
rect 10401 7575 10402 7601
rect 10374 7574 10402 7575
rect 11606 9646 11634 9674
rect 12726 11185 12754 11186
rect 12726 11159 12727 11185
rect 12727 11159 12753 11185
rect 12753 11159 12754 11185
rect 12726 11158 12754 11159
rect 12054 9673 12082 9674
rect 12054 9647 12055 9673
rect 12055 9647 12081 9673
rect 12081 9647 12082 9673
rect 12054 9646 12082 9647
rect 12166 10934 12194 10962
rect 11830 9617 11858 9618
rect 11830 9591 11831 9617
rect 11831 9591 11857 9617
rect 11857 9591 11858 9617
rect 11830 9590 11858 9591
rect 11438 9310 11466 9338
rect 11606 9366 11634 9394
rect 11774 9505 11802 9506
rect 11774 9479 11775 9505
rect 11775 9479 11801 9505
rect 11801 9479 11802 9505
rect 11774 9478 11802 9479
rect 11382 9225 11410 9226
rect 11382 9199 11383 9225
rect 11383 9199 11409 9225
rect 11409 9199 11410 9225
rect 11382 9198 11410 9199
rect 11998 9366 12026 9394
rect 12054 9478 12082 9506
rect 11830 9310 11858 9338
rect 12110 8806 12138 8834
rect 11550 8777 11578 8778
rect 11550 8751 11551 8777
rect 11551 8751 11577 8777
rect 11577 8751 11578 8777
rect 11550 8750 11578 8751
rect 11942 8777 11970 8778
rect 11942 8751 11943 8777
rect 11943 8751 11969 8777
rect 11969 8751 11970 8777
rect 11942 8750 11970 8751
rect 11046 8526 11074 8554
rect 11438 8694 11466 8722
rect 10990 8414 11018 8442
rect 10654 7574 10682 7602
rect 11382 8134 11410 8162
rect 12670 10654 12698 10682
rect 12894 11942 12922 11970
rect 13566 13033 13594 13034
rect 13566 13007 13567 13033
rect 13567 13007 13593 13033
rect 13593 13007 13594 13033
rect 13566 13006 13594 13007
rect 14518 13089 14546 13090
rect 14518 13063 14519 13089
rect 14519 13063 14545 13089
rect 14545 13063 14546 13089
rect 14518 13062 14546 13063
rect 14966 13062 14994 13090
rect 13678 12782 13706 12810
rect 14070 12809 14098 12810
rect 14070 12783 14071 12809
rect 14071 12783 14097 12809
rect 14097 12783 14098 12809
rect 14070 12782 14098 12783
rect 13342 12726 13370 12754
rect 13342 12473 13370 12474
rect 13342 12447 13343 12473
rect 13343 12447 13369 12473
rect 13369 12447 13370 12473
rect 13342 12446 13370 12447
rect 13398 12670 13426 12698
rect 14462 12670 14490 12698
rect 13510 12446 13538 12474
rect 13622 11969 13650 11970
rect 13622 11943 13623 11969
rect 13623 11943 13649 11969
rect 13649 11943 13650 11969
rect 13622 11942 13650 11943
rect 17598 12949 17626 12950
rect 17598 12923 17599 12949
rect 17599 12923 17625 12949
rect 17625 12923 17626 12949
rect 17598 12922 17626 12923
rect 17650 12949 17678 12950
rect 17650 12923 17651 12949
rect 17651 12923 17677 12949
rect 17677 12923 17678 12949
rect 17650 12922 17678 12923
rect 17702 12949 17730 12950
rect 17702 12923 17703 12949
rect 17703 12923 17729 12949
rect 17729 12923 17730 12949
rect 17702 12922 17730 12923
rect 20006 13118 20034 13146
rect 18942 13062 18970 13090
rect 18830 12782 18858 12810
rect 20006 12782 20034 12810
rect 17598 12165 17626 12166
rect 17598 12139 17599 12165
rect 17599 12139 17625 12165
rect 17625 12139 17626 12165
rect 17598 12138 17626 12139
rect 17650 12165 17678 12166
rect 17650 12139 17651 12165
rect 17651 12139 17677 12165
rect 17677 12139 17678 12165
rect 17650 12138 17678 12139
rect 17702 12165 17730 12166
rect 17702 12139 17703 12165
rect 17703 12139 17729 12165
rect 17729 12139 17730 12165
rect 17702 12138 17730 12139
rect 13118 11774 13146 11802
rect 12838 11073 12866 11074
rect 12838 11047 12839 11073
rect 12839 11047 12865 11073
rect 12865 11047 12866 11073
rect 12838 11046 12866 11047
rect 12950 11129 12978 11130
rect 12950 11103 12951 11129
rect 12951 11103 12977 11129
rect 12977 11103 12978 11129
rect 12950 11102 12978 11103
rect 13622 11158 13650 11186
rect 17598 11381 17626 11382
rect 17598 11355 17599 11381
rect 17599 11355 17625 11381
rect 17625 11355 17626 11381
rect 17598 11354 17626 11355
rect 17650 11381 17678 11382
rect 17650 11355 17651 11381
rect 17651 11355 17677 11381
rect 17677 11355 17678 11381
rect 17650 11354 17678 11355
rect 17702 11381 17730 11382
rect 17702 11355 17703 11381
rect 17703 11355 17729 11381
rect 17729 11355 17730 11381
rect 17702 11354 17730 11355
rect 14070 11185 14098 11186
rect 14070 11159 14071 11185
rect 14071 11159 14097 11185
rect 14097 11159 14098 11185
rect 14070 11158 14098 11159
rect 14798 11158 14826 11186
rect 12894 10457 12922 10458
rect 12894 10431 12895 10457
rect 12895 10431 12921 10457
rect 12921 10431 12922 10457
rect 12894 10430 12922 10431
rect 12726 10401 12754 10402
rect 12726 10375 12727 10401
rect 12727 10375 12753 10401
rect 12753 10375 12754 10401
rect 12726 10374 12754 10375
rect 13230 10430 13258 10458
rect 12614 10094 12642 10122
rect 11830 8721 11858 8722
rect 11830 8695 11831 8721
rect 11831 8695 11857 8721
rect 11857 8695 11858 8721
rect 11830 8694 11858 8695
rect 12614 8750 12642 8778
rect 11886 8105 11914 8106
rect 11886 8079 11887 8105
rect 11887 8079 11913 8105
rect 11913 8079 11914 8105
rect 11886 8078 11914 8079
rect 12726 8638 12754 8666
rect 13398 10038 13426 10066
rect 13118 9646 13146 9674
rect 13230 9870 13258 9898
rect 13230 9617 13258 9618
rect 13230 9591 13231 9617
rect 13231 9591 13257 9617
rect 13257 9591 13258 9617
rect 13230 9590 13258 9591
rect 18830 11185 18858 11186
rect 18830 11159 18831 11185
rect 18831 11159 18857 11185
rect 18857 11159 18858 11185
rect 18830 11158 18858 11159
rect 20006 11102 20034 11130
rect 17598 10597 17626 10598
rect 17598 10571 17599 10597
rect 17599 10571 17625 10597
rect 17625 10571 17626 10597
rect 17598 10570 17626 10571
rect 17650 10597 17678 10598
rect 17650 10571 17651 10597
rect 17651 10571 17677 10597
rect 17677 10571 17678 10597
rect 17650 10570 17678 10571
rect 17702 10597 17730 10598
rect 17702 10571 17703 10597
rect 17703 10571 17729 10597
rect 17729 10571 17730 10597
rect 17702 10570 17730 10571
rect 13902 10038 13930 10066
rect 13510 9926 13538 9954
rect 13454 9673 13482 9674
rect 13454 9647 13455 9673
rect 13455 9647 13481 9673
rect 13481 9647 13482 9673
rect 13454 9646 13482 9647
rect 13790 9617 13818 9618
rect 13790 9591 13791 9617
rect 13791 9591 13817 9617
rect 13817 9591 13818 9617
rect 13790 9590 13818 9591
rect 14686 10065 14714 10066
rect 14686 10039 14687 10065
rect 14687 10039 14713 10065
rect 14713 10039 14714 10065
rect 14686 10038 14714 10039
rect 20006 10094 20034 10122
rect 18942 10038 18970 10066
rect 14574 10009 14602 10010
rect 14574 9983 14575 10009
rect 14575 9983 14601 10009
rect 14601 9983 14602 10009
rect 14574 9982 14602 9983
rect 18830 10009 18858 10010
rect 18830 9983 18831 10009
rect 18831 9983 18857 10009
rect 18857 9983 18858 10009
rect 18830 9982 18858 9983
rect 14350 9953 14378 9954
rect 14350 9927 14351 9953
rect 14351 9927 14377 9953
rect 14377 9927 14378 9953
rect 14350 9926 14378 9927
rect 17598 9813 17626 9814
rect 17598 9787 17599 9813
rect 17599 9787 17625 9813
rect 17625 9787 17626 9813
rect 17598 9786 17626 9787
rect 17650 9813 17678 9814
rect 17650 9787 17651 9813
rect 17651 9787 17677 9813
rect 17677 9787 17678 9813
rect 17650 9786 17678 9787
rect 17702 9813 17730 9814
rect 17702 9787 17703 9813
rect 17703 9787 17729 9813
rect 17729 9787 17730 9813
rect 17702 9786 17730 9787
rect 20006 9758 20034 9786
rect 14014 9561 14042 9562
rect 14014 9535 14015 9561
rect 14015 9535 14041 9561
rect 14041 9535 14042 9561
rect 14014 9534 14042 9535
rect 13622 9505 13650 9506
rect 13622 9479 13623 9505
rect 13623 9479 13649 9505
rect 13649 9479 13650 9505
rect 13622 9478 13650 9479
rect 14742 9561 14770 9562
rect 14742 9535 14743 9561
rect 14743 9535 14769 9561
rect 14769 9535 14770 9561
rect 14742 9534 14770 9535
rect 14574 9478 14602 9506
rect 14574 9254 14602 9282
rect 20006 9422 20034 9450
rect 18830 9254 18858 9282
rect 12838 8553 12866 8554
rect 12838 8527 12839 8553
rect 12839 8527 12865 8553
rect 12865 8527 12866 8553
rect 12838 8526 12866 8527
rect 12726 8497 12754 8498
rect 12726 8471 12727 8497
rect 12727 8471 12753 8497
rect 12753 8471 12754 8497
rect 12726 8470 12754 8471
rect 12334 8414 12362 8442
rect 12166 8358 12194 8386
rect 12670 8385 12698 8386
rect 12670 8359 12671 8385
rect 12671 8359 12697 8385
rect 12697 8359 12698 8385
rect 12670 8358 12698 8359
rect 12222 8078 12250 8106
rect 11046 7937 11074 7938
rect 11046 7911 11047 7937
rect 11047 7911 11073 7937
rect 11073 7911 11074 7937
rect 11046 7910 11074 7911
rect 10990 7350 11018 7378
rect 11494 7910 11522 7938
rect 12558 8078 12586 8106
rect 17598 9029 17626 9030
rect 17598 9003 17599 9029
rect 17599 9003 17625 9029
rect 17625 9003 17626 9029
rect 17598 9002 17626 9003
rect 17650 9029 17678 9030
rect 17650 9003 17651 9029
rect 17651 9003 17677 9029
rect 17677 9003 17678 9029
rect 17650 9002 17678 9003
rect 17702 9029 17730 9030
rect 17702 9003 17703 9029
rect 17703 9003 17729 9029
rect 17729 9003 17730 9029
rect 17702 9002 17730 9003
rect 13118 8441 13146 8442
rect 13118 8415 13119 8441
rect 13119 8415 13145 8441
rect 13145 8415 13146 8441
rect 13118 8414 13146 8415
rect 13566 8441 13594 8442
rect 13566 8415 13567 8441
rect 13567 8415 13593 8441
rect 13593 8415 13594 8441
rect 13566 8414 13594 8415
rect 12950 8078 12978 8106
rect 11438 7657 11466 7658
rect 11438 7631 11439 7657
rect 11439 7631 11465 7657
rect 11465 7631 11466 7657
rect 11438 7630 11466 7631
rect 11270 7350 11298 7378
rect 12110 7518 12138 7546
rect 12278 7377 12306 7378
rect 12278 7351 12279 7377
rect 12279 7351 12305 7377
rect 12305 7351 12306 7377
rect 12278 7350 12306 7351
rect 13678 8358 13706 8386
rect 14070 8414 14098 8442
rect 18942 8414 18970 8442
rect 20006 8414 20034 8442
rect 18830 8358 18858 8386
rect 17598 8245 17626 8246
rect 17598 8219 17599 8245
rect 17599 8219 17625 8245
rect 17625 8219 17626 8245
rect 17598 8218 17626 8219
rect 17650 8245 17678 8246
rect 17650 8219 17651 8245
rect 17651 8219 17677 8245
rect 17677 8219 17678 8245
rect 17650 8218 17678 8219
rect 17702 8245 17730 8246
rect 17702 8219 17703 8245
rect 17703 8219 17729 8245
rect 17729 8219 17730 8245
rect 17702 8218 17730 8219
rect 19950 8078 19978 8106
rect 13678 7713 13706 7714
rect 13678 7687 13679 7713
rect 13679 7687 13705 7713
rect 13705 7687 13706 7713
rect 13678 7686 13706 7687
rect 20006 7742 20034 7770
rect 18830 7686 18858 7714
rect 17598 7461 17626 7462
rect 17598 7435 17599 7461
rect 17599 7435 17625 7461
rect 17625 7435 17626 7461
rect 17598 7434 17626 7435
rect 17650 7461 17678 7462
rect 17650 7435 17651 7461
rect 17651 7435 17677 7461
rect 17677 7435 17678 7461
rect 17650 7434 17678 7435
rect 17702 7461 17730 7462
rect 17702 7435 17703 7461
rect 17703 7435 17729 7461
rect 17729 7435 17730 7461
rect 17702 7434 17730 7435
rect 12334 6734 12362 6762
rect 8414 2030 8442 2058
rect 2238 1973 2266 1974
rect 2238 1947 2239 1973
rect 2239 1947 2265 1973
rect 2265 1947 2266 1973
rect 2238 1946 2266 1947
rect 2290 1973 2318 1974
rect 2290 1947 2291 1973
rect 2291 1947 2317 1973
rect 2317 1947 2318 1973
rect 2290 1946 2318 1947
rect 2342 1973 2370 1974
rect 2342 1947 2343 1973
rect 2343 1947 2369 1973
rect 2369 1947 2370 1973
rect 2342 1946 2370 1947
rect 9918 3933 9946 3934
rect 9918 3907 9919 3933
rect 9919 3907 9945 3933
rect 9945 3907 9946 3933
rect 9918 3906 9946 3907
rect 9970 3933 9998 3934
rect 9970 3907 9971 3933
rect 9971 3907 9997 3933
rect 9997 3907 9998 3933
rect 9970 3906 9998 3907
rect 10022 3933 10050 3934
rect 10022 3907 10023 3933
rect 10023 3907 10049 3933
rect 10049 3907 10050 3933
rect 10022 3906 10050 3907
rect 9918 3149 9946 3150
rect 9918 3123 9919 3149
rect 9919 3123 9945 3149
rect 9945 3123 9946 3149
rect 9918 3122 9946 3123
rect 9970 3149 9998 3150
rect 9970 3123 9971 3149
rect 9971 3123 9997 3149
rect 9997 3123 9998 3149
rect 9970 3122 9998 3123
rect 10022 3149 10050 3150
rect 10022 3123 10023 3149
rect 10023 3123 10049 3149
rect 10049 3123 10050 3149
rect 10022 3122 10050 3123
rect 9918 2365 9946 2366
rect 9918 2339 9919 2365
rect 9919 2339 9945 2365
rect 9945 2339 9946 2365
rect 9918 2338 9946 2339
rect 9970 2365 9998 2366
rect 9970 2339 9971 2365
rect 9971 2339 9997 2365
rect 9997 2339 9998 2365
rect 9970 2338 9998 2339
rect 10022 2365 10050 2366
rect 10022 2339 10023 2365
rect 10023 2339 10049 2365
rect 10049 2339 10050 2365
rect 10022 2338 10050 2339
rect 9198 2057 9226 2058
rect 9198 2031 9199 2057
rect 9199 2031 9225 2057
rect 9225 2031 9226 2057
rect 9198 2030 9226 2031
rect 9758 1806 9786 1834
rect 10934 1833 10962 1834
rect 10934 1807 10935 1833
rect 10935 1807 10961 1833
rect 10961 1807 10962 1833
rect 10934 1806 10962 1807
rect 11438 1806 11466 1834
rect 9918 1581 9946 1582
rect 9918 1555 9919 1581
rect 9919 1555 9945 1581
rect 9945 1555 9946 1581
rect 9918 1554 9946 1555
rect 9970 1581 9998 1582
rect 9970 1555 9971 1581
rect 9971 1555 9997 1581
rect 9997 1555 9998 1581
rect 9970 1554 9998 1555
rect 10022 1581 10050 1582
rect 10022 1555 10023 1581
rect 10023 1555 10049 1581
rect 10049 1555 10050 1581
rect 10022 1554 10050 1555
rect 12950 6734 12978 6762
rect 17598 6677 17626 6678
rect 17598 6651 17599 6677
rect 17599 6651 17625 6677
rect 17625 6651 17626 6677
rect 17598 6650 17626 6651
rect 17650 6677 17678 6678
rect 17650 6651 17651 6677
rect 17651 6651 17677 6677
rect 17677 6651 17678 6677
rect 17650 6650 17678 6651
rect 17702 6677 17730 6678
rect 17702 6651 17703 6677
rect 17703 6651 17729 6677
rect 17729 6651 17730 6677
rect 17702 6650 17730 6651
rect 17598 5893 17626 5894
rect 17598 5867 17599 5893
rect 17599 5867 17625 5893
rect 17625 5867 17626 5893
rect 17598 5866 17626 5867
rect 17650 5893 17678 5894
rect 17650 5867 17651 5893
rect 17651 5867 17677 5893
rect 17677 5867 17678 5893
rect 17650 5866 17678 5867
rect 17702 5893 17730 5894
rect 17702 5867 17703 5893
rect 17703 5867 17729 5893
rect 17729 5867 17730 5893
rect 17702 5866 17730 5867
rect 17598 5109 17626 5110
rect 17598 5083 17599 5109
rect 17599 5083 17625 5109
rect 17625 5083 17626 5109
rect 17598 5082 17626 5083
rect 17650 5109 17678 5110
rect 17650 5083 17651 5109
rect 17651 5083 17677 5109
rect 17677 5083 17678 5109
rect 17650 5082 17678 5083
rect 17702 5109 17730 5110
rect 17702 5083 17703 5109
rect 17703 5083 17729 5109
rect 17729 5083 17730 5109
rect 17702 5082 17730 5083
rect 17598 4325 17626 4326
rect 17598 4299 17599 4325
rect 17599 4299 17625 4325
rect 17625 4299 17626 4325
rect 17598 4298 17626 4299
rect 17650 4325 17678 4326
rect 17650 4299 17651 4325
rect 17651 4299 17677 4325
rect 17677 4299 17678 4325
rect 17650 4298 17678 4299
rect 17702 4325 17730 4326
rect 17702 4299 17703 4325
rect 17703 4299 17729 4325
rect 17729 4299 17730 4325
rect 17702 4298 17730 4299
rect 17598 3541 17626 3542
rect 17598 3515 17599 3541
rect 17599 3515 17625 3541
rect 17625 3515 17626 3541
rect 17598 3514 17626 3515
rect 17650 3541 17678 3542
rect 17650 3515 17651 3541
rect 17651 3515 17677 3541
rect 17677 3515 17678 3541
rect 17650 3514 17678 3515
rect 17702 3541 17730 3542
rect 17702 3515 17703 3541
rect 17703 3515 17729 3541
rect 17729 3515 17730 3541
rect 17702 3514 17730 3515
rect 17598 2757 17626 2758
rect 17598 2731 17599 2757
rect 17599 2731 17625 2757
rect 17625 2731 17626 2757
rect 17598 2730 17626 2731
rect 17650 2757 17678 2758
rect 17650 2731 17651 2757
rect 17651 2731 17677 2757
rect 17677 2731 17678 2757
rect 17650 2730 17678 2731
rect 17702 2757 17730 2758
rect 17702 2731 17703 2757
rect 17703 2731 17729 2757
rect 17729 2731 17730 2757
rect 17702 2730 17730 2731
rect 12446 2030 12474 2058
rect 13118 2057 13146 2058
rect 13118 2031 13119 2057
rect 13119 2031 13145 2057
rect 13145 2031 13146 2057
rect 13118 2030 13146 2031
rect 17598 1973 17626 1974
rect 17598 1947 17599 1973
rect 17599 1947 17625 1973
rect 17625 1947 17626 1973
rect 17598 1946 17626 1947
rect 17650 1973 17678 1974
rect 17650 1947 17651 1973
rect 17651 1947 17677 1973
rect 17677 1947 17678 1973
rect 17650 1946 17678 1947
rect 17702 1973 17730 1974
rect 17702 1947 17703 1973
rect 17703 1947 17729 1973
rect 17729 1947 17730 1973
rect 17702 1946 17730 1947
rect 12782 1833 12810 1834
rect 12782 1807 12783 1833
rect 12783 1807 12809 1833
rect 12809 1807 12810 1833
rect 12782 1806 12810 1807
<< metal3 >>
rect 2233 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2375 19222
rect 17593 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17735 19222
rect 12441 19110 12446 19138
rect 12474 19110 13062 19138
rect 13090 19110 13095 19138
rect 9913 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10055 18830
rect 8745 18718 8750 18746
rect 8778 18718 9366 18746
rect 9394 18718 9399 18746
rect 10761 18718 10766 18746
rect 10794 18718 11382 18746
rect 11410 18718 11415 18746
rect 2233 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2375 18438
rect 17593 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17735 18438
rect 9913 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10055 18046
rect 2233 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2375 17654
rect 17593 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17735 17654
rect 9913 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10055 17262
rect 2233 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2375 16870
rect 17593 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17735 16870
rect 9913 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10055 16478
rect 2233 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2375 16086
rect 17593 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17735 16086
rect 9913 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10055 15694
rect 2233 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2375 15302
rect 17593 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17735 15302
rect 9913 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10055 14910
rect 10705 14630 10710 14658
rect 10738 14630 11046 14658
rect 11074 14630 11079 14658
rect 2233 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2375 14518
rect 17593 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17735 14518
rect 8358 14294 8526 14322
rect 8554 14294 9618 14322
rect 8358 14266 8386 14294
rect 9590 14266 9618 14294
rect 7681 14238 7686 14266
rect 7714 14238 8386 14266
rect 9585 14238 9590 14266
rect 9618 14238 10934 14266
rect 10962 14238 11214 14266
rect 11242 14238 11247 14266
rect 9913 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10055 14126
rect 7009 13902 7014 13930
rect 7042 13902 7686 13930
rect 7714 13902 7719 13930
rect 8409 13846 8414 13874
rect 8442 13846 9254 13874
rect 9282 13846 9287 13874
rect 0 13818 400 13832
rect 0 13790 2086 13818
rect 2114 13790 2119 13818
rect 0 13776 400 13790
rect 2233 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2375 13734
rect 17593 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17735 13734
rect 2137 13510 2142 13538
rect 2170 13510 6286 13538
rect 6314 13510 6319 13538
rect 8134 13454 9198 13482
rect 9226 13454 9231 13482
rect 9361 13454 9366 13482
rect 9394 13454 10654 13482
rect 10682 13454 10687 13482
rect 8134 13370 8162 13454
rect 9366 13426 9394 13454
rect 8801 13398 8806 13426
rect 8834 13398 9394 13426
rect 8129 13342 8134 13370
rect 8162 13342 8167 13370
rect 9913 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10055 13342
rect 7345 13230 7350 13258
rect 7378 13230 7966 13258
rect 7994 13230 7999 13258
rect 10649 13230 10654 13258
rect 10682 13230 10990 13258
rect 11018 13230 11023 13258
rect 9921 13174 9926 13202
rect 9954 13174 10542 13202
rect 10570 13174 10575 13202
rect 12329 13174 12334 13202
rect 12362 13174 12670 13202
rect 12698 13174 12703 13202
rect 0 13146 400 13160
rect 20600 13146 21000 13160
rect 0 13118 966 13146
rect 994 13118 999 13146
rect 9137 13118 9142 13146
rect 9170 13118 9870 13146
rect 9898 13118 9903 13146
rect 10705 13118 10710 13146
rect 10738 13118 10990 13146
rect 11018 13118 12726 13146
rect 12754 13118 13510 13146
rect 13538 13118 13543 13146
rect 20001 13118 20006 13146
rect 20034 13118 21000 13146
rect 0 13104 400 13118
rect 20600 13104 21000 13118
rect 6281 13062 6286 13090
rect 6314 13062 7854 13090
rect 7882 13062 7887 13090
rect 11265 13062 11270 13090
rect 11298 13062 11774 13090
rect 11802 13062 11807 13090
rect 14513 13062 14518 13090
rect 14546 13062 14966 13090
rect 14994 13062 18942 13090
rect 18970 13062 18975 13090
rect 12049 13006 12054 13034
rect 12082 13006 12670 13034
rect 12698 13006 12703 13034
rect 13169 13006 13174 13034
rect 13202 13006 13566 13034
rect 13594 13006 13599 13034
rect 2233 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2375 12950
rect 17593 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17735 12950
rect 7345 12838 7350 12866
rect 7378 12838 8246 12866
rect 8274 12838 8279 12866
rect 20600 12810 21000 12824
rect 13673 12782 13678 12810
rect 13706 12782 14070 12810
rect 14098 12782 18830 12810
rect 18858 12782 18863 12810
rect 20001 12782 20006 12810
rect 20034 12782 21000 12810
rect 20600 12768 21000 12782
rect 7905 12726 7910 12754
rect 7938 12726 8190 12754
rect 8218 12726 8223 12754
rect 10929 12726 10934 12754
rect 10962 12726 12446 12754
rect 12474 12726 12670 12754
rect 12698 12726 12950 12754
rect 12978 12726 13342 12754
rect 13370 12726 13375 12754
rect 8241 12670 8246 12698
rect 8274 12670 8806 12698
rect 8834 12670 10206 12698
rect 10234 12670 10239 12698
rect 13393 12670 13398 12698
rect 13426 12670 14462 12698
rect 14490 12670 14495 12698
rect 9913 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10055 12558
rect 13337 12446 13342 12474
rect 13370 12446 13510 12474
rect 13538 12446 13543 12474
rect 8073 12278 8078 12306
rect 8106 12278 8806 12306
rect 8834 12278 8839 12306
rect 2233 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2375 12166
rect 17593 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17735 12166
rect 8409 12110 8414 12138
rect 8442 12110 9030 12138
rect 9058 12110 9063 12138
rect 8857 12054 8862 12082
rect 8890 12054 9478 12082
rect 9506 12054 11830 12082
rect 11858 12054 11863 12082
rect 10481 11998 10486 12026
rect 10514 11998 10822 12026
rect 10850 11998 10855 12026
rect 2137 11942 2142 11970
rect 2170 11942 6734 11970
rect 6762 11942 8078 11970
rect 8106 11942 8111 11970
rect 12889 11942 12894 11970
rect 12922 11942 13622 11970
rect 13650 11942 13655 11970
rect 7793 11886 7798 11914
rect 7826 11886 8470 11914
rect 8498 11886 8503 11914
rect 8745 11886 8750 11914
rect 8778 11886 9142 11914
rect 9170 11886 9175 11914
rect 9417 11886 9422 11914
rect 9450 11886 9982 11914
rect 10010 11886 10015 11914
rect 8129 11830 8134 11858
rect 8162 11830 8414 11858
rect 8442 11830 8447 11858
rect 8521 11830 8526 11858
rect 8554 11830 8918 11858
rect 8946 11830 8951 11858
rect 0 11802 400 11816
rect 0 11774 966 11802
rect 994 11774 999 11802
rect 12665 11774 12670 11802
rect 12698 11774 13118 11802
rect 13146 11774 13151 11802
rect 0 11760 400 11774
rect 9913 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10055 11774
rect 8241 11718 8246 11746
rect 8274 11718 8862 11746
rect 8890 11718 8895 11746
rect 9081 11718 9086 11746
rect 9114 11718 9119 11746
rect 9086 11690 9114 11718
rect 8582 11662 9114 11690
rect 8582 11634 8610 11662
rect 5889 11606 5894 11634
rect 5922 11606 8414 11634
rect 8442 11606 8582 11634
rect 8610 11606 8615 11634
rect 8969 11606 8974 11634
rect 9002 11606 9422 11634
rect 9450 11606 9455 11634
rect 7177 11550 7182 11578
rect 7210 11550 7406 11578
rect 7434 11550 8190 11578
rect 8218 11550 8358 11578
rect 8386 11550 9254 11578
rect 9282 11550 10486 11578
rect 10514 11550 10519 11578
rect 6953 11494 6958 11522
rect 6986 11494 7518 11522
rect 7546 11494 7551 11522
rect 9641 11494 9646 11522
rect 9674 11494 10878 11522
rect 10906 11494 10911 11522
rect 8857 11438 8862 11466
rect 8890 11438 8918 11466
rect 8946 11438 8951 11466
rect 2233 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2375 11382
rect 17593 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17735 11382
rect 9417 11214 9422 11242
rect 9450 11214 10318 11242
rect 10346 11214 11214 11242
rect 11242 11214 11886 11242
rect 11914 11214 11919 11242
rect 7849 11158 7854 11186
rect 7882 11158 8918 11186
rect 8946 11158 8951 11186
rect 9921 11158 9926 11186
rect 9954 11158 10934 11186
rect 10962 11158 11438 11186
rect 11466 11158 11471 11186
rect 11601 11158 11606 11186
rect 11634 11158 12726 11186
rect 12754 11158 12759 11186
rect 13426 11158 13622 11186
rect 13650 11158 13655 11186
rect 14065 11158 14070 11186
rect 14098 11158 14798 11186
rect 14826 11158 18830 11186
rect 18858 11158 18863 11186
rect 13426 11130 13454 11158
rect 20600 11130 21000 11144
rect 10145 11102 10150 11130
rect 10178 11102 12950 11130
rect 12978 11102 13454 11130
rect 20001 11102 20006 11130
rect 20034 11102 21000 11130
rect 20600 11088 21000 11102
rect 9081 11046 9086 11074
rect 9114 11046 9758 11074
rect 9786 11046 10094 11074
rect 10122 11046 10127 11074
rect 11825 11046 11830 11074
rect 11858 11046 12838 11074
rect 12866 11046 12871 11074
rect 9913 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10055 10990
rect 5553 10934 5558 10962
rect 5586 10934 5838 10962
rect 5866 10934 7462 10962
rect 7490 10934 7495 10962
rect 8409 10934 8414 10962
rect 8442 10934 8582 10962
rect 8610 10934 8615 10962
rect 11153 10934 11158 10962
rect 11186 10934 11718 10962
rect 11746 10934 12166 10962
rect 12194 10934 12199 10962
rect 7233 10878 7238 10906
rect 7266 10878 7742 10906
rect 7770 10878 8246 10906
rect 8274 10878 8806 10906
rect 8834 10878 8839 10906
rect 9473 10878 9478 10906
rect 9506 10878 9926 10906
rect 9954 10878 9959 10906
rect 7681 10822 7686 10850
rect 7714 10822 8302 10850
rect 8330 10822 8694 10850
rect 8722 10822 8727 10850
rect 2081 10766 2086 10794
rect 2114 10766 9478 10794
rect 9506 10766 9702 10794
rect 9730 10766 9735 10794
rect 6169 10710 6174 10738
rect 6202 10710 6846 10738
rect 6874 10710 6879 10738
rect 8969 10654 8974 10682
rect 9002 10654 11886 10682
rect 11914 10654 12670 10682
rect 12698 10654 12703 10682
rect 2233 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2375 10598
rect 17593 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17735 10598
rect 9697 10486 9702 10514
rect 9730 10486 10934 10514
rect 10962 10486 10967 10514
rect 10201 10430 10206 10458
rect 10234 10430 11382 10458
rect 11410 10430 11662 10458
rect 11690 10430 11695 10458
rect 12889 10430 12894 10458
rect 12922 10430 13230 10458
rect 13258 10430 13263 10458
rect 9809 10374 9814 10402
rect 9842 10374 9926 10402
rect 9954 10374 9959 10402
rect 10705 10374 10710 10402
rect 10738 10374 11102 10402
rect 11130 10374 11135 10402
rect 11937 10374 11942 10402
rect 11970 10374 12726 10402
rect 12754 10374 12759 10402
rect 8409 10318 8414 10346
rect 8442 10318 8862 10346
rect 8890 10318 8895 10346
rect 9913 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10055 10206
rect 20600 10122 21000 10136
rect 9305 10094 9310 10122
rect 9338 10094 11382 10122
rect 11410 10094 12614 10122
rect 12642 10094 12647 10122
rect 20001 10094 20006 10122
rect 20034 10094 21000 10122
rect 20600 10080 21000 10094
rect 7121 10038 7126 10066
rect 7154 10038 7686 10066
rect 7714 10038 7719 10066
rect 9865 10038 9870 10066
rect 9898 10038 10262 10066
rect 10290 10038 10295 10066
rect 10374 10038 10822 10066
rect 10850 10038 13398 10066
rect 13426 10038 13902 10066
rect 13930 10038 13935 10066
rect 14681 10038 14686 10066
rect 14714 10038 18942 10066
rect 18970 10038 18975 10066
rect 10374 10010 10402 10038
rect 2137 9982 2142 10010
rect 2170 9982 4998 10010
rect 5026 9982 5031 10010
rect 7065 9982 7070 10010
rect 7098 9982 7238 10010
rect 7266 9982 7966 10010
rect 7994 9982 7999 10010
rect 10089 9982 10094 10010
rect 10122 9982 10402 10010
rect 10705 9982 10710 10010
rect 10738 9982 11046 10010
rect 11074 9982 11606 10010
rect 11634 9982 11639 10010
rect 14569 9982 14574 10010
rect 14602 9982 18830 10010
rect 18858 9982 18863 10010
rect 6057 9926 6062 9954
rect 6090 9926 7014 9954
rect 7042 9926 7047 9954
rect 7681 9926 7686 9954
rect 7714 9926 9366 9954
rect 9394 9926 9399 9954
rect 13505 9926 13510 9954
rect 13538 9926 14350 9954
rect 14378 9926 14383 9954
rect 961 9870 966 9898
rect 994 9870 999 9898
rect 7177 9870 7182 9898
rect 7210 9870 7910 9898
rect 7938 9870 10878 9898
rect 10906 9870 13230 9898
rect 13258 9870 13263 9898
rect 0 9786 400 9800
rect 966 9786 994 9870
rect 2233 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2375 9814
rect 17593 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17735 9814
rect 20600 9786 21000 9800
rect 0 9758 994 9786
rect 8465 9758 8470 9786
rect 8498 9758 9142 9786
rect 9170 9758 9814 9786
rect 9842 9758 9847 9786
rect 20001 9758 20006 9786
rect 20034 9758 21000 9786
rect 0 9744 400 9758
rect 20600 9744 21000 9758
rect 8857 9702 8862 9730
rect 8890 9702 9758 9730
rect 9786 9702 9791 9730
rect 8017 9646 8022 9674
rect 8050 9646 8302 9674
rect 8330 9646 8694 9674
rect 8722 9646 8727 9674
rect 11601 9646 11606 9674
rect 11634 9646 12054 9674
rect 12082 9646 12087 9674
rect 13113 9646 13118 9674
rect 13146 9646 13454 9674
rect 13482 9646 13487 9674
rect 6449 9590 6454 9618
rect 6482 9590 6790 9618
rect 6818 9590 6823 9618
rect 8577 9590 8582 9618
rect 8610 9590 8918 9618
rect 8946 9590 8951 9618
rect 9025 9590 9030 9618
rect 9058 9590 9590 9618
rect 9618 9590 9623 9618
rect 11209 9590 11214 9618
rect 11242 9590 11830 9618
rect 11858 9590 11863 9618
rect 13225 9590 13230 9618
rect 13258 9590 13790 9618
rect 13818 9590 13823 9618
rect 4993 9534 4998 9562
rect 5026 9534 7294 9562
rect 7322 9534 7327 9562
rect 8857 9534 8862 9562
rect 8890 9534 9310 9562
rect 9338 9534 10038 9562
rect 10066 9534 10071 9562
rect 14009 9534 14014 9562
rect 14042 9534 14742 9562
rect 14770 9534 14775 9562
rect 9025 9478 9030 9506
rect 9058 9478 9814 9506
rect 9842 9478 9847 9506
rect 10817 9478 10822 9506
rect 10850 9478 11158 9506
rect 11186 9478 11774 9506
rect 11802 9478 11807 9506
rect 12049 9478 12054 9506
rect 12082 9478 13622 9506
rect 13650 9478 14574 9506
rect 14602 9478 14607 9506
rect 20600 9450 21000 9464
rect 8241 9422 8246 9450
rect 8274 9422 9086 9450
rect 9114 9422 9119 9450
rect 20001 9422 20006 9450
rect 20034 9422 21000 9450
rect 9913 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10055 9422
rect 20600 9408 21000 9422
rect 11601 9366 11606 9394
rect 11634 9366 11998 9394
rect 12026 9366 12031 9394
rect 6505 9310 6510 9338
rect 6538 9310 7238 9338
rect 7266 9310 7271 9338
rect 8745 9310 8750 9338
rect 8778 9310 11102 9338
rect 11130 9310 11438 9338
rect 11466 9310 11830 9338
rect 11858 9310 11863 9338
rect 7289 9254 7294 9282
rect 7322 9254 8134 9282
rect 8162 9254 8167 9282
rect 9473 9254 9478 9282
rect 9506 9254 9814 9282
rect 9842 9254 9926 9282
rect 9954 9254 9959 9282
rect 14569 9254 14574 9282
rect 14602 9254 18830 9282
rect 18858 9254 18863 9282
rect 7233 9198 7238 9226
rect 7266 9198 8862 9226
rect 8890 9198 8895 9226
rect 8969 9198 8974 9226
rect 9002 9198 9254 9226
rect 9282 9198 9287 9226
rect 10817 9198 10822 9226
rect 10850 9198 11382 9226
rect 11410 9198 11415 9226
rect 6897 9142 6902 9170
rect 6930 9142 7742 9170
rect 7770 9142 7775 9170
rect 9179 9142 9198 9170
rect 9226 9142 9231 9170
rect 10089 9142 10094 9170
rect 10122 9142 10990 9170
rect 11018 9142 11023 9170
rect 7625 9086 7630 9114
rect 7658 9086 7854 9114
rect 7882 9086 8358 9114
rect 8386 9086 10934 9114
rect 10962 9086 10967 9114
rect 7401 9030 7406 9058
rect 7434 9030 9366 9058
rect 9394 9030 9399 9058
rect 2233 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2375 9030
rect 17593 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17735 9030
rect 6785 8918 6790 8946
rect 6818 8918 7126 8946
rect 7154 8918 7159 8946
rect 961 8862 966 8890
rect 994 8862 999 8890
rect 7233 8862 7238 8890
rect 7266 8862 8414 8890
rect 8442 8862 8447 8890
rect 9025 8862 9030 8890
rect 9058 8862 9198 8890
rect 9226 8862 9231 8890
rect 0 8778 400 8792
rect 966 8778 994 8862
rect 2137 8806 2142 8834
rect 2170 8806 5446 8834
rect 5474 8806 6734 8834
rect 6762 8806 6767 8834
rect 6841 8806 6846 8834
rect 6874 8806 7406 8834
rect 7434 8806 7439 8834
rect 8801 8806 8806 8834
rect 8834 8806 12110 8834
rect 12138 8806 12143 8834
rect 0 8750 994 8778
rect 5385 8750 5390 8778
rect 5418 8750 7574 8778
rect 7602 8750 7607 8778
rect 9305 8750 9310 8778
rect 9338 8750 11550 8778
rect 11578 8750 11942 8778
rect 11970 8750 12614 8778
rect 12642 8750 12647 8778
rect 0 8736 400 8750
rect 6505 8694 6510 8722
rect 6538 8694 7406 8722
rect 7434 8694 7439 8722
rect 8521 8694 8526 8722
rect 8554 8694 9254 8722
rect 9282 8694 9287 8722
rect 9585 8694 9590 8722
rect 9618 8694 9702 8722
rect 9730 8694 10822 8722
rect 10850 8694 10855 8722
rect 11433 8694 11438 8722
rect 11466 8694 11830 8722
rect 11858 8694 11863 8722
rect 7121 8638 7126 8666
rect 7154 8638 7742 8666
rect 7770 8638 7775 8666
rect 10985 8638 10990 8666
rect 11018 8638 12726 8666
rect 12754 8638 12759 8666
rect 9913 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10055 8638
rect 9081 8582 9086 8610
rect 9114 8582 9198 8610
rect 9226 8582 9231 8610
rect 8409 8526 8414 8554
rect 8442 8526 11046 8554
rect 11074 8526 12838 8554
rect 12866 8526 12871 8554
rect 12721 8470 12726 8498
rect 12754 8470 13594 8498
rect 0 8442 400 8456
rect 13566 8442 13594 8470
rect 20600 8442 21000 8456
rect 0 8414 966 8442
rect 994 8414 999 8442
rect 2137 8414 2142 8442
rect 2170 8414 5390 8442
rect 5418 8414 5423 8442
rect 8843 8414 8862 8442
rect 8890 8414 8895 8442
rect 9249 8414 9254 8442
rect 9282 8414 10766 8442
rect 10794 8414 10990 8442
rect 11018 8414 11023 8442
rect 12329 8414 12334 8442
rect 12362 8414 13118 8442
rect 13146 8414 13151 8442
rect 13561 8414 13566 8442
rect 13594 8414 14070 8442
rect 14098 8414 18942 8442
rect 18970 8414 18975 8442
rect 20001 8414 20006 8442
rect 20034 8414 21000 8442
rect 0 8400 400 8414
rect 20600 8400 21000 8414
rect 7345 8358 7350 8386
rect 7378 8358 7798 8386
rect 7826 8358 7831 8386
rect 8969 8358 8974 8386
rect 9002 8358 9422 8386
rect 9450 8358 9455 8386
rect 12161 8358 12166 8386
rect 12194 8358 12670 8386
rect 12698 8358 12703 8386
rect 13673 8358 13678 8386
rect 13706 8358 18830 8386
rect 18858 8358 18863 8386
rect 2233 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2375 8246
rect 17593 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17735 8246
rect 8073 8134 8078 8162
rect 8106 8134 8414 8162
rect 8442 8134 8447 8162
rect 10705 8134 10710 8162
rect 10738 8134 11382 8162
rect 11410 8134 11415 8162
rect 20600 8106 21000 8120
rect 10649 8078 10654 8106
rect 10682 8078 11886 8106
rect 11914 8078 12222 8106
rect 12250 8078 12558 8106
rect 12586 8078 12950 8106
rect 12978 8078 12983 8106
rect 19945 8078 19950 8106
rect 19978 8078 21000 8106
rect 20600 8064 21000 8078
rect 9473 7910 9478 7938
rect 9506 7910 10150 7938
rect 10178 7910 10183 7938
rect 11041 7910 11046 7938
rect 11074 7910 11494 7938
rect 11522 7910 11527 7938
rect 9913 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10055 7854
rect 20600 7770 21000 7784
rect 20001 7742 20006 7770
rect 20034 7742 21000 7770
rect 20600 7728 21000 7742
rect 13673 7686 13678 7714
rect 13706 7686 18830 7714
rect 18858 7686 18863 7714
rect 11433 7630 11438 7658
rect 11466 7630 12138 7658
rect 7065 7574 7070 7602
rect 7098 7574 8750 7602
rect 8778 7574 10094 7602
rect 10122 7574 10374 7602
rect 10402 7574 10654 7602
rect 10682 7574 10687 7602
rect 12110 7546 12138 7630
rect 12105 7518 12110 7546
rect 12138 7518 12143 7546
rect 2233 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2375 7462
rect 17593 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17735 7462
rect 10985 7350 10990 7378
rect 11018 7350 11270 7378
rect 11298 7350 12278 7378
rect 12306 7350 12311 7378
rect 8129 7126 8134 7154
rect 8162 7126 8582 7154
rect 8610 7126 8615 7154
rect 9913 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10055 7070
rect 12329 6734 12334 6762
rect 12362 6734 12950 6762
rect 12978 6734 12983 6762
rect 2233 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2375 6678
rect 17593 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17735 6678
rect 10066 6482 10094 6538
rect 10122 6510 10127 6538
rect 7793 6454 7798 6482
rect 7826 6454 9478 6482
rect 9506 6454 10094 6482
rect 9913 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10055 6286
rect 2233 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2375 5894
rect 17593 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17735 5894
rect 9913 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10055 5502
rect 2233 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2375 5110
rect 17593 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17735 5110
rect 9913 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10055 4718
rect 2233 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2375 4326
rect 17593 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17735 4326
rect 9913 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10055 3934
rect 2233 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2375 3542
rect 17593 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17735 3542
rect 9913 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10055 3150
rect 2233 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2375 2758
rect 17593 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17735 2758
rect 9913 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10055 2366
rect 8409 2030 8414 2058
rect 8442 2030 9198 2058
rect 9226 2030 9231 2058
rect 12441 2030 12446 2058
rect 12474 2030 13118 2058
rect 13146 2030 13151 2058
rect 2233 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2375 1974
rect 17593 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17735 1974
rect 9753 1806 9758 1834
rect 9786 1806 10934 1834
rect 10962 1806 10967 1834
rect 11433 1806 11438 1834
rect 11466 1806 12782 1834
rect 12810 1806 12815 1834
rect 9913 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10055 1582
<< via3 >>
rect 2238 19194 2266 19222
rect 2290 19194 2318 19222
rect 2342 19194 2370 19222
rect 17598 19194 17626 19222
rect 17650 19194 17678 19222
rect 17702 19194 17730 19222
rect 9918 18802 9946 18830
rect 9970 18802 9998 18830
rect 10022 18802 10050 18830
rect 2238 18410 2266 18438
rect 2290 18410 2318 18438
rect 2342 18410 2370 18438
rect 17598 18410 17626 18438
rect 17650 18410 17678 18438
rect 17702 18410 17730 18438
rect 9918 18018 9946 18046
rect 9970 18018 9998 18046
rect 10022 18018 10050 18046
rect 2238 17626 2266 17654
rect 2290 17626 2318 17654
rect 2342 17626 2370 17654
rect 17598 17626 17626 17654
rect 17650 17626 17678 17654
rect 17702 17626 17730 17654
rect 9918 17234 9946 17262
rect 9970 17234 9998 17262
rect 10022 17234 10050 17262
rect 2238 16842 2266 16870
rect 2290 16842 2318 16870
rect 2342 16842 2370 16870
rect 17598 16842 17626 16870
rect 17650 16842 17678 16870
rect 17702 16842 17730 16870
rect 9918 16450 9946 16478
rect 9970 16450 9998 16478
rect 10022 16450 10050 16478
rect 2238 16058 2266 16086
rect 2290 16058 2318 16086
rect 2342 16058 2370 16086
rect 17598 16058 17626 16086
rect 17650 16058 17678 16086
rect 17702 16058 17730 16086
rect 9918 15666 9946 15694
rect 9970 15666 9998 15694
rect 10022 15666 10050 15694
rect 2238 15274 2266 15302
rect 2290 15274 2318 15302
rect 2342 15274 2370 15302
rect 17598 15274 17626 15302
rect 17650 15274 17678 15302
rect 17702 15274 17730 15302
rect 9918 14882 9946 14910
rect 9970 14882 9998 14910
rect 10022 14882 10050 14910
rect 2238 14490 2266 14518
rect 2290 14490 2318 14518
rect 2342 14490 2370 14518
rect 17598 14490 17626 14518
rect 17650 14490 17678 14518
rect 17702 14490 17730 14518
rect 9918 14098 9946 14126
rect 9970 14098 9998 14126
rect 10022 14098 10050 14126
rect 2238 13706 2266 13734
rect 2290 13706 2318 13734
rect 2342 13706 2370 13734
rect 17598 13706 17626 13734
rect 17650 13706 17678 13734
rect 17702 13706 17730 13734
rect 9918 13314 9946 13342
rect 9970 13314 9998 13342
rect 10022 13314 10050 13342
rect 2238 12922 2266 12950
rect 2290 12922 2318 12950
rect 2342 12922 2370 12950
rect 17598 12922 17626 12950
rect 17650 12922 17678 12950
rect 17702 12922 17730 12950
rect 9918 12530 9946 12558
rect 9970 12530 9998 12558
rect 10022 12530 10050 12558
rect 2238 12138 2266 12166
rect 2290 12138 2318 12166
rect 2342 12138 2370 12166
rect 17598 12138 17626 12166
rect 17650 12138 17678 12166
rect 17702 12138 17730 12166
rect 9918 11746 9946 11774
rect 9970 11746 9998 11774
rect 10022 11746 10050 11774
rect 8862 11438 8890 11466
rect 2238 11354 2266 11382
rect 2290 11354 2318 11382
rect 2342 11354 2370 11382
rect 17598 11354 17626 11382
rect 17650 11354 17678 11382
rect 17702 11354 17730 11382
rect 9918 10962 9946 10990
rect 9970 10962 9998 10990
rect 10022 10962 10050 10990
rect 2238 10570 2266 10598
rect 2290 10570 2318 10598
rect 2342 10570 2370 10598
rect 17598 10570 17626 10598
rect 17650 10570 17678 10598
rect 17702 10570 17730 10598
rect 9814 10374 9842 10402
rect 9918 10178 9946 10206
rect 9970 10178 9998 10206
rect 10022 10178 10050 10206
rect 2238 9786 2266 9814
rect 2290 9786 2318 9814
rect 2342 9786 2370 9814
rect 17598 9786 17626 9814
rect 17650 9786 17678 9814
rect 17702 9786 17730 9814
rect 9590 9590 9618 9618
rect 9918 9394 9946 9422
rect 9970 9394 9998 9422
rect 10022 9394 10050 9422
rect 9814 9254 9842 9282
rect 9198 9142 9226 9170
rect 2238 9002 2266 9030
rect 2290 9002 2318 9030
rect 2342 9002 2370 9030
rect 17598 9002 17626 9030
rect 17650 9002 17678 9030
rect 17702 9002 17730 9030
rect 9590 8694 9618 8722
rect 9918 8610 9946 8638
rect 9970 8610 9998 8638
rect 10022 8610 10050 8638
rect 9198 8582 9226 8610
rect 8862 8414 8890 8442
rect 2238 8218 2266 8246
rect 2290 8218 2318 8246
rect 2342 8218 2370 8246
rect 17598 8218 17626 8246
rect 17650 8218 17678 8246
rect 17702 8218 17730 8246
rect 9918 7826 9946 7854
rect 9970 7826 9998 7854
rect 10022 7826 10050 7854
rect 2238 7434 2266 7462
rect 2290 7434 2318 7462
rect 2342 7434 2370 7462
rect 17598 7434 17626 7462
rect 17650 7434 17678 7462
rect 17702 7434 17730 7462
rect 9918 7042 9946 7070
rect 9970 7042 9998 7070
rect 10022 7042 10050 7070
rect 2238 6650 2266 6678
rect 2290 6650 2318 6678
rect 2342 6650 2370 6678
rect 17598 6650 17626 6678
rect 17650 6650 17678 6678
rect 17702 6650 17730 6678
rect 9918 6258 9946 6286
rect 9970 6258 9998 6286
rect 10022 6258 10050 6286
rect 2238 5866 2266 5894
rect 2290 5866 2318 5894
rect 2342 5866 2370 5894
rect 17598 5866 17626 5894
rect 17650 5866 17678 5894
rect 17702 5866 17730 5894
rect 9918 5474 9946 5502
rect 9970 5474 9998 5502
rect 10022 5474 10050 5502
rect 2238 5082 2266 5110
rect 2290 5082 2318 5110
rect 2342 5082 2370 5110
rect 17598 5082 17626 5110
rect 17650 5082 17678 5110
rect 17702 5082 17730 5110
rect 9918 4690 9946 4718
rect 9970 4690 9998 4718
rect 10022 4690 10050 4718
rect 2238 4298 2266 4326
rect 2290 4298 2318 4326
rect 2342 4298 2370 4326
rect 17598 4298 17626 4326
rect 17650 4298 17678 4326
rect 17702 4298 17730 4326
rect 9918 3906 9946 3934
rect 9970 3906 9998 3934
rect 10022 3906 10050 3934
rect 2238 3514 2266 3542
rect 2290 3514 2318 3542
rect 2342 3514 2370 3542
rect 17598 3514 17626 3542
rect 17650 3514 17678 3542
rect 17702 3514 17730 3542
rect 9918 3122 9946 3150
rect 9970 3122 9998 3150
rect 10022 3122 10050 3150
rect 2238 2730 2266 2758
rect 2290 2730 2318 2758
rect 2342 2730 2370 2758
rect 17598 2730 17626 2758
rect 17650 2730 17678 2758
rect 17702 2730 17730 2758
rect 9918 2338 9946 2366
rect 9970 2338 9998 2366
rect 10022 2338 10050 2366
rect 2238 1946 2266 1974
rect 2290 1946 2318 1974
rect 2342 1946 2370 1974
rect 17598 1946 17626 1974
rect 17650 1946 17678 1974
rect 17702 1946 17730 1974
rect 9918 1554 9946 1582
rect 9970 1554 9998 1582
rect 10022 1554 10050 1582
<< metal4 >>
rect 2224 19222 2384 19238
rect 2224 19194 2238 19222
rect 2266 19194 2290 19222
rect 2318 19194 2342 19222
rect 2370 19194 2384 19222
rect 2224 18438 2384 19194
rect 2224 18410 2238 18438
rect 2266 18410 2290 18438
rect 2318 18410 2342 18438
rect 2370 18410 2384 18438
rect 2224 17654 2384 18410
rect 2224 17626 2238 17654
rect 2266 17626 2290 17654
rect 2318 17626 2342 17654
rect 2370 17626 2384 17654
rect 2224 16870 2384 17626
rect 2224 16842 2238 16870
rect 2266 16842 2290 16870
rect 2318 16842 2342 16870
rect 2370 16842 2384 16870
rect 2224 16086 2384 16842
rect 2224 16058 2238 16086
rect 2266 16058 2290 16086
rect 2318 16058 2342 16086
rect 2370 16058 2384 16086
rect 2224 15302 2384 16058
rect 2224 15274 2238 15302
rect 2266 15274 2290 15302
rect 2318 15274 2342 15302
rect 2370 15274 2384 15302
rect 2224 14518 2384 15274
rect 2224 14490 2238 14518
rect 2266 14490 2290 14518
rect 2318 14490 2342 14518
rect 2370 14490 2384 14518
rect 2224 13734 2384 14490
rect 2224 13706 2238 13734
rect 2266 13706 2290 13734
rect 2318 13706 2342 13734
rect 2370 13706 2384 13734
rect 2224 12950 2384 13706
rect 2224 12922 2238 12950
rect 2266 12922 2290 12950
rect 2318 12922 2342 12950
rect 2370 12922 2384 12950
rect 2224 12166 2384 12922
rect 2224 12138 2238 12166
rect 2266 12138 2290 12166
rect 2318 12138 2342 12166
rect 2370 12138 2384 12166
rect 2224 11382 2384 12138
rect 9904 18830 10064 19238
rect 9904 18802 9918 18830
rect 9946 18802 9970 18830
rect 9998 18802 10022 18830
rect 10050 18802 10064 18830
rect 9904 18046 10064 18802
rect 9904 18018 9918 18046
rect 9946 18018 9970 18046
rect 9998 18018 10022 18046
rect 10050 18018 10064 18046
rect 9904 17262 10064 18018
rect 9904 17234 9918 17262
rect 9946 17234 9970 17262
rect 9998 17234 10022 17262
rect 10050 17234 10064 17262
rect 9904 16478 10064 17234
rect 9904 16450 9918 16478
rect 9946 16450 9970 16478
rect 9998 16450 10022 16478
rect 10050 16450 10064 16478
rect 9904 15694 10064 16450
rect 9904 15666 9918 15694
rect 9946 15666 9970 15694
rect 9998 15666 10022 15694
rect 10050 15666 10064 15694
rect 9904 14910 10064 15666
rect 9904 14882 9918 14910
rect 9946 14882 9970 14910
rect 9998 14882 10022 14910
rect 10050 14882 10064 14910
rect 9904 14126 10064 14882
rect 9904 14098 9918 14126
rect 9946 14098 9970 14126
rect 9998 14098 10022 14126
rect 10050 14098 10064 14126
rect 9904 13342 10064 14098
rect 9904 13314 9918 13342
rect 9946 13314 9970 13342
rect 9998 13314 10022 13342
rect 10050 13314 10064 13342
rect 9904 12558 10064 13314
rect 9904 12530 9918 12558
rect 9946 12530 9970 12558
rect 9998 12530 10022 12558
rect 10050 12530 10064 12558
rect 9904 11774 10064 12530
rect 9904 11746 9918 11774
rect 9946 11746 9970 11774
rect 9998 11746 10022 11774
rect 10050 11746 10064 11774
rect 2224 11354 2238 11382
rect 2266 11354 2290 11382
rect 2318 11354 2342 11382
rect 2370 11354 2384 11382
rect 2224 10598 2384 11354
rect 2224 10570 2238 10598
rect 2266 10570 2290 10598
rect 2318 10570 2342 10598
rect 2370 10570 2384 10598
rect 2224 9814 2384 10570
rect 2224 9786 2238 9814
rect 2266 9786 2290 9814
rect 2318 9786 2342 9814
rect 2370 9786 2384 9814
rect 2224 9030 2384 9786
rect 2224 9002 2238 9030
rect 2266 9002 2290 9030
rect 2318 9002 2342 9030
rect 2370 9002 2384 9030
rect 2224 8246 2384 9002
rect 8862 11466 8890 11471
rect 8862 8442 8890 11438
rect 9904 10990 10064 11746
rect 9904 10962 9918 10990
rect 9946 10962 9970 10990
rect 9998 10962 10022 10990
rect 10050 10962 10064 10990
rect 9814 10402 9842 10407
rect 9590 9618 9618 9623
rect 9198 9170 9226 9175
rect 9198 8610 9226 9142
rect 9590 8722 9618 9590
rect 9814 9282 9842 10374
rect 9814 9249 9842 9254
rect 9904 10206 10064 10962
rect 9904 10178 9918 10206
rect 9946 10178 9970 10206
rect 9998 10178 10022 10206
rect 10050 10178 10064 10206
rect 9904 9422 10064 10178
rect 9904 9394 9918 9422
rect 9946 9394 9970 9422
rect 9998 9394 10022 9422
rect 10050 9394 10064 9422
rect 9590 8689 9618 8694
rect 9198 8577 9226 8582
rect 9904 8638 10064 9394
rect 9904 8610 9918 8638
rect 9946 8610 9970 8638
rect 9998 8610 10022 8638
rect 10050 8610 10064 8638
rect 8862 8409 8890 8414
rect 2224 8218 2238 8246
rect 2266 8218 2290 8246
rect 2318 8218 2342 8246
rect 2370 8218 2384 8246
rect 2224 7462 2384 8218
rect 2224 7434 2238 7462
rect 2266 7434 2290 7462
rect 2318 7434 2342 7462
rect 2370 7434 2384 7462
rect 2224 6678 2384 7434
rect 2224 6650 2238 6678
rect 2266 6650 2290 6678
rect 2318 6650 2342 6678
rect 2370 6650 2384 6678
rect 2224 5894 2384 6650
rect 2224 5866 2238 5894
rect 2266 5866 2290 5894
rect 2318 5866 2342 5894
rect 2370 5866 2384 5894
rect 2224 5110 2384 5866
rect 2224 5082 2238 5110
rect 2266 5082 2290 5110
rect 2318 5082 2342 5110
rect 2370 5082 2384 5110
rect 2224 4326 2384 5082
rect 2224 4298 2238 4326
rect 2266 4298 2290 4326
rect 2318 4298 2342 4326
rect 2370 4298 2384 4326
rect 2224 3542 2384 4298
rect 2224 3514 2238 3542
rect 2266 3514 2290 3542
rect 2318 3514 2342 3542
rect 2370 3514 2384 3542
rect 2224 2758 2384 3514
rect 2224 2730 2238 2758
rect 2266 2730 2290 2758
rect 2318 2730 2342 2758
rect 2370 2730 2384 2758
rect 2224 1974 2384 2730
rect 2224 1946 2238 1974
rect 2266 1946 2290 1974
rect 2318 1946 2342 1974
rect 2370 1946 2384 1974
rect 2224 1538 2384 1946
rect 9904 7854 10064 8610
rect 9904 7826 9918 7854
rect 9946 7826 9970 7854
rect 9998 7826 10022 7854
rect 10050 7826 10064 7854
rect 9904 7070 10064 7826
rect 9904 7042 9918 7070
rect 9946 7042 9970 7070
rect 9998 7042 10022 7070
rect 10050 7042 10064 7070
rect 9904 6286 10064 7042
rect 9904 6258 9918 6286
rect 9946 6258 9970 6286
rect 9998 6258 10022 6286
rect 10050 6258 10064 6286
rect 9904 5502 10064 6258
rect 9904 5474 9918 5502
rect 9946 5474 9970 5502
rect 9998 5474 10022 5502
rect 10050 5474 10064 5502
rect 9904 4718 10064 5474
rect 9904 4690 9918 4718
rect 9946 4690 9970 4718
rect 9998 4690 10022 4718
rect 10050 4690 10064 4718
rect 9904 3934 10064 4690
rect 9904 3906 9918 3934
rect 9946 3906 9970 3934
rect 9998 3906 10022 3934
rect 10050 3906 10064 3934
rect 9904 3150 10064 3906
rect 9904 3122 9918 3150
rect 9946 3122 9970 3150
rect 9998 3122 10022 3150
rect 10050 3122 10064 3150
rect 9904 2366 10064 3122
rect 9904 2338 9918 2366
rect 9946 2338 9970 2366
rect 9998 2338 10022 2366
rect 10050 2338 10064 2366
rect 9904 1582 10064 2338
rect 9904 1554 9918 1582
rect 9946 1554 9970 1582
rect 9998 1554 10022 1582
rect 10050 1554 10064 1582
rect 9904 1538 10064 1554
rect 17584 19222 17744 19238
rect 17584 19194 17598 19222
rect 17626 19194 17650 19222
rect 17678 19194 17702 19222
rect 17730 19194 17744 19222
rect 17584 18438 17744 19194
rect 17584 18410 17598 18438
rect 17626 18410 17650 18438
rect 17678 18410 17702 18438
rect 17730 18410 17744 18438
rect 17584 17654 17744 18410
rect 17584 17626 17598 17654
rect 17626 17626 17650 17654
rect 17678 17626 17702 17654
rect 17730 17626 17744 17654
rect 17584 16870 17744 17626
rect 17584 16842 17598 16870
rect 17626 16842 17650 16870
rect 17678 16842 17702 16870
rect 17730 16842 17744 16870
rect 17584 16086 17744 16842
rect 17584 16058 17598 16086
rect 17626 16058 17650 16086
rect 17678 16058 17702 16086
rect 17730 16058 17744 16086
rect 17584 15302 17744 16058
rect 17584 15274 17598 15302
rect 17626 15274 17650 15302
rect 17678 15274 17702 15302
rect 17730 15274 17744 15302
rect 17584 14518 17744 15274
rect 17584 14490 17598 14518
rect 17626 14490 17650 14518
rect 17678 14490 17702 14518
rect 17730 14490 17744 14518
rect 17584 13734 17744 14490
rect 17584 13706 17598 13734
rect 17626 13706 17650 13734
rect 17678 13706 17702 13734
rect 17730 13706 17744 13734
rect 17584 12950 17744 13706
rect 17584 12922 17598 12950
rect 17626 12922 17650 12950
rect 17678 12922 17702 12950
rect 17730 12922 17744 12950
rect 17584 12166 17744 12922
rect 17584 12138 17598 12166
rect 17626 12138 17650 12166
rect 17678 12138 17702 12166
rect 17730 12138 17744 12166
rect 17584 11382 17744 12138
rect 17584 11354 17598 11382
rect 17626 11354 17650 11382
rect 17678 11354 17702 11382
rect 17730 11354 17744 11382
rect 17584 10598 17744 11354
rect 17584 10570 17598 10598
rect 17626 10570 17650 10598
rect 17678 10570 17702 10598
rect 17730 10570 17744 10598
rect 17584 9814 17744 10570
rect 17584 9786 17598 9814
rect 17626 9786 17650 9814
rect 17678 9786 17702 9814
rect 17730 9786 17744 9814
rect 17584 9030 17744 9786
rect 17584 9002 17598 9030
rect 17626 9002 17650 9030
rect 17678 9002 17702 9030
rect 17730 9002 17744 9030
rect 17584 8246 17744 9002
rect 17584 8218 17598 8246
rect 17626 8218 17650 8246
rect 17678 8218 17702 8246
rect 17730 8218 17744 8246
rect 17584 7462 17744 8218
rect 17584 7434 17598 7462
rect 17626 7434 17650 7462
rect 17678 7434 17702 7462
rect 17730 7434 17744 7462
rect 17584 6678 17744 7434
rect 17584 6650 17598 6678
rect 17626 6650 17650 6678
rect 17678 6650 17702 6678
rect 17730 6650 17744 6678
rect 17584 5894 17744 6650
rect 17584 5866 17598 5894
rect 17626 5866 17650 5894
rect 17678 5866 17702 5894
rect 17730 5866 17744 5894
rect 17584 5110 17744 5866
rect 17584 5082 17598 5110
rect 17626 5082 17650 5110
rect 17678 5082 17702 5110
rect 17730 5082 17744 5110
rect 17584 4326 17744 5082
rect 17584 4298 17598 4326
rect 17626 4298 17650 4326
rect 17678 4298 17702 4326
rect 17730 4298 17744 4326
rect 17584 3542 17744 4298
rect 17584 3514 17598 3542
rect 17626 3514 17650 3542
rect 17678 3514 17702 3542
rect 17730 3514 17744 3542
rect 17584 2758 17744 3514
rect 17584 2730 17598 2758
rect 17626 2730 17650 2758
rect 17678 2730 17702 2758
rect 17730 2730 17744 2758
rect 17584 1974 17744 2730
rect 17584 1946 17598 1974
rect 17626 1946 17650 1974
rect 17678 1946 17702 1974
rect 17730 1946 17744 1974
rect 17584 1538 17744 1946
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _104_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11928 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _105_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11256 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _106_
timestamp 1698175906
transform -1 0 10192 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _107_
timestamp 1698175906
transform -1 0 12152 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _108_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9352 0 1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _109_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _110_
timestamp 1698175906
transform -1 0 12040 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _111_
timestamp 1698175906
transform -1 0 12152 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _112_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 11760 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _113_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10584 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _114_
timestamp 1698175906
transform 1 0 10696 0 1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _115_
timestamp 1698175906
transform -1 0 12824 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _116_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11648 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _117_
timestamp 1698175906
transform 1 0 8176 0 -1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _118_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9856 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _119_
timestamp 1698175906
transform -1 0 9072 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _120_
timestamp 1698175906
transform 1 0 8120 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _121_
timestamp 1698175906
transform 1 0 7616 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_2  _122_
timestamp 1698175906
transform 1 0 8792 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_2  _123_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8960 0 1 9408
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _124_
timestamp 1698175906
transform -1 0 9128 0 -1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _125_
timestamp 1698175906
transform -1 0 11704 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _126_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8568 0 1 9408
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _127_
timestamp 1698175906
transform -1 0 8120 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _128_
timestamp 1698175906
transform 1 0 7952 0 -1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _129_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 8960 0 1 11760
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _130_
timestamp 1698175906
transform 1 0 11760 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _131_
timestamp 1698175906
transform 1 0 14504 0 1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_2  _132_
timestamp 1698175906
transform 1 0 11032 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_4  _133_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9408 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _134_
timestamp 1698175906
transform 1 0 9856 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _135_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13776 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _136_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 8008 0 -1 10976
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _137_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 7112 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _138_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8736 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _139_
timestamp 1698175906
transform 1 0 9688 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _140_
timestamp 1698175906
transform -1 0 11536 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _141_
timestamp 1698175906
transform 1 0 9184 0 1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _142_
timestamp 1698175906
transform 1 0 9912 0 1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _143_
timestamp 1698175906
transform -1 0 11032 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_2  _144_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11536 0 -1 10192
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _145_
timestamp 1698175906
transform 1 0 11032 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_1  _146_
timestamp 1698175906
transform 1 0 11368 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _147_
timestamp 1698175906
transform -1 0 10976 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _148_
timestamp 1698175906
transform -1 0 11816 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _149_
timestamp 1698175906
transform 1 0 9072 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _150_
timestamp 1698175906
transform -1 0 11312 0 -1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _151_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 9352 0 1 7056
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _152_
timestamp 1698175906
transform -1 0 8736 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _153_
timestamp 1698175906
transform 1 0 13440 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _154_
timestamp 1698175906
transform 1 0 12768 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _155_
timestamp 1698175906
transform -1 0 10472 0 1 12544
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _156_
timestamp 1698175906
transform 1 0 10584 0 1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _157_
timestamp 1698175906
transform -1 0 10416 0 1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _158_
timestamp 1698175906
transform -1 0 10808 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _159_
timestamp 1698175906
transform -1 0 9408 0 1 11760
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _160_
timestamp 1698175906
transform 1 0 9800 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _161_
timestamp 1698175906
transform -1 0 9184 0 1 10192
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _162_
timestamp 1698175906
transform -1 0 9464 0 1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _163_
timestamp 1698175906
transform -1 0 8232 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _164_
timestamp 1698175906
transform 1 0 12208 0 1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _165_
timestamp 1698175906
transform -1 0 12096 0 1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__xor2_1  _166_
timestamp 1698175906
transform -1 0 11256 0 1 8624
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _167_
timestamp 1698175906
transform 1 0 11312 0 1 7840
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _168_
timestamp 1698175906
transform 1 0 11536 0 -1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__aoi21_2  _169_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9072 0 1 8624
box -43 -43 771 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _170_
timestamp 1698175906
transform -1 0 7448 0 1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _171_
timestamp 1698175906
transform -1 0 8512 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _172_
timestamp 1698175906
transform -1 0 7784 0 -1 10192
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _173_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 7504 0 -1 10192
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _174_
timestamp 1698175906
transform -1 0 7672 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _175_
timestamp 1698175906
transform 1 0 9688 0 1 9408
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _176_
timestamp 1698175906
transform -1 0 9072 0 1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _177_
timestamp 1698175906
transform -1 0 8400 0 1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__aoi221_1  _178_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 7000 0 -1 9408
box -43 -43 659 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _179_
timestamp 1698175906
transform -1 0 8736 0 1 8624
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _180_
timestamp 1698175906
transform -1 0 6944 0 1 8624
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _181_
timestamp 1698175906
transform -1 0 7168 0 1 9408
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand4_1  _182_
timestamp 1698175906
transform 1 0 6944 0 1 8624
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _183_
timestamp 1698175906
transform -1 0 8904 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _184_
timestamp 1698175906
transform -1 0 8512 0 -1 13328
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _185_
timestamp 1698175906
transform 1 0 7784 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _186_
timestamp 1698175906
transform 1 0 8008 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__aoi22_1  _187_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform -1 0 8512 0 1 12544
box -43 -43 547 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _188_
timestamp 1698175906
transform -1 0 9688 0 1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai22_1  _189_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8792 0 -1 8624
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _190_
timestamp 1698175906
transform 1 0 12544 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__or2_1  _191_
timestamp 1698175906
transform 1 0 11984 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _192_
timestamp 1698175906
transform -1 0 13216 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _193_
timestamp 1698175906
transform 1 0 12544 0 -1 10976
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _194_
timestamp 1698175906
transform 1 0 13328 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _195_
timestamp 1698175906
transform 1 0 12656 0 1 10192
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__nand3_1  _196_
timestamp 1698175906
transform -1 0 8736 0 1 7840
box -43 -43 435 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _197_
timestamp 1698175906
transform 1 0 7672 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__oai21_1  _198_
timestamp 1698175906
transform 1 0 10024 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _199_
timestamp 1698175906
transform 1 0 13832 0 1 10976
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _200_
timestamp 1698175906
transform -1 0 13888 0 -1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__nor2_1  _201_
timestamp 1698175906
transform 1 0 11200 0 -1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__oai32_1  _202_
timestamp 1698175906
transform 1 0 10640 0 1 7840
box -43 -43 715 435
use gf180mcu_fd_sc_mcu7t5v0__oai211_1  _203_
timestamp 1698175906
transform 1 0 12656 0 1 10976
box -43 -43 603 435
use gf180mcu_fd_sc_mcu7t5v0__clkinv_1  _204_
timestamp 1698175906
transform -1 0 14616 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__nand2_1  _205_
timestamp 1698175906
transform 1 0 13272 0 1 11760
box -43 -43 323 435
use gf180mcu_fd_sc_mcu7t5v0__and2_1  _206_
timestamp 1698175906
transform 1 0 13552 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_1  _207_
timestamp 1698175906
transform -1 0 14336 0 1 11760
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _208_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10808 0 -1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _209_
timestamp 1698175906
transform -1 0 8288 0 1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _210_
timestamp 1698175906
transform 1 0 13048 0 -1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _211_
timestamp 1698175906
transform 1 0 5432 0 -1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _212_
timestamp 1698175906
transform 1 0 5712 0 -1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _213_
timestamp 1698175906
transform 1 0 9184 0 -1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _214_
timestamp 1698175906
transform 1 0 10808 0 -1 11760
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _215_
timestamp 1698175906
transform 1 0 7672 0 1 6272
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _216_
timestamp 1698175906
transform 1 0 12544 0 1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _217_
timestamp 1698175906
transform 1 0 9520 0 -1 14896
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _218_
timestamp 1698175906
transform 1 0 9464 0 -1 14112
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _219_
timestamp 1698175906
transform 1 0 6888 0 -1 14112
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _220_
timestamp 1698175906
transform 1 0 10808 0 -1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _221_
timestamp 1698175906
transform -1 0 6552 0 1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _222_
timestamp 1698175906
transform -1 0 7000 0 -1 9408
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _223_
timestamp 1698175906
transform -1 0 7000 0 -1 8624
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _224_
timestamp 1698175906
transform 1 0 7560 0 1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _225_
timestamp 1698175906
transform -1 0 7840 0 -1 13328
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _226_
timestamp 1698175906
transform 1 0 8624 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_2  _227_ dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 12488 0 1 7840
box -43 -43 1779 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _228_
timestamp 1698175906
transform 1 0 12824 0 -1 10192
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _229_
timestamp 1698175906
transform 1 0 6888 0 -1 7840
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _230_
timestamp 1698175906
transform 1 0 13272 0 -1 10976
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _231_
timestamp 1698175906
transform 1 0 10584 0 1 7056
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__dffq_1  _232_
timestamp 1698175906
transform 1 0 13440 0 -1 12544
box -43 -43 1667 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _233_
timestamp 1698175906
transform -1 0 9128 0 -1 14112
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _234_
timestamp 1698175906
transform 1 0 13440 0 -1 7840
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _235_
timestamp 1698175906
transform 1 0 14448 0 -1 10192
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _236_
timestamp 1698175906
transform 1 0 12544 0 1 7056
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__buf_1  _237_
timestamp 1698175906
transform 1 0 13440 0 -1 8624
box -43 -43 379 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__135__A2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 13216 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__173__A2
timestamp 1698175906
transform 1 0 7896 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__186__A1
timestamp 1698175906
transform -1 0 8848 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__208__CLK
timestamp 1698175906
transform 1 0 12936 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__209__CLK
timestamp 1698175906
transform 1 0 8344 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__210__CLK
timestamp 1698175906
transform 1 0 12936 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__211__CLK
timestamp 1698175906
transform 1 0 7168 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__212__CLK
timestamp 1698175906
transform -1 0 7448 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__213__CLK
timestamp 1698175906
transform 1 0 10808 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__214__CLK
timestamp 1698175906
transform 1 0 12656 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__215__CLK
timestamp 1698175906
transform -1 0 9520 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__216__CLK
timestamp 1698175906
transform 1 0 12432 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__217__CLK
timestamp 1698175906
transform -1 0 11368 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__218__CLK
timestamp 1698175906
transform 1 0 11200 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__219__CLK
timestamp 1698175906
transform 1 0 8512 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__220__CLK
timestamp 1698175906
transform 1 0 12656 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__221__CLK
timestamp 1698175906
transform 1 0 6776 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__222__CLK
timestamp 1698175906
transform 1 0 7728 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__223__CLK
timestamp 1698175906
transform 1 0 7112 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__224__CLK
timestamp 1698175906
transform 1 0 9576 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__225__CLK
timestamp 1698175906
transform 1 0 7672 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__226__CLK
timestamp 1698175906
transform 1 0 10360 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__227__CLK
timestamp 1698175906
transform 1 0 11872 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__228__CLK
timestamp 1698175906
transform -1 0 12824 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__229__CLK
timestamp 1698175906
transform 1 0 8848 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__230__CLK
timestamp 1698175906
transform 1 0 13160 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__231__CLK
timestamp 1698175906
transform 1 0 12208 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA__232__CLK
timestamp 1698175906
transform 1 0 13328 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__antenna  ANTENNA_clkbuf_0_clk_I
timestamp 1698175906
transform 1 0 9464 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_0_clk dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 9576 0 -1 10976
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_0__f_clk
timestamp 1698175906
transform 1 0 9464 0 -1 8624
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__clkbuf_16  clkbuf_1_1__f_clk
timestamp 1698175906
transform 1 0 9408 0 -1 12544
box -43 -43 2843 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_36
timestamp 1698175906
transform 1 0 2688 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_70
timestamp 1698175906
transform 1 0 4592 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_104
timestamp 1698175906
transform 1 0 6496 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_138 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8400 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_142 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8624 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_198
timestamp 1698175906
transform 1 0 11760 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_202
timestamp 1698175906
transform 1 0 11984 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_232
timestamp 1698175906
transform 1 0 13664 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_236
timestamp 1698175906
transform 1 0 13888 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_240
timestamp 1698175906
transform 1 0 14112 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_274
timestamp 1698175906
transform 1 0 16016 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_0_308
timestamp 1698175906
transform 1 0 17920 0 1 1568
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_0_342
timestamp 1698175906
transform 1 0 19824 0 1 1568
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_0_346
timestamp 1698175906
transform 1 0 20048 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_0_348 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 20160 0 1 1568
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_2 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 784 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_66
timestamp 1698175906
transform 1 0 4368 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_72
timestamp 1698175906
transform 1 0 4704 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_1_136
timestamp 1698175906
transform 1 0 8288 0 -1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_168
timestamp 1698175906
transform 1 0 10080 0 -1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_200 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 11872 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_208
timestamp 1698175906
transform 1 0 12320 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_1_238
timestamp 1698175906
transform 1 0 14000 0 -1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_1_270
timestamp 1698175906
transform 1 0 15792 0 -1 2352
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_278
timestamp 1698175906
transform 1 0 16240 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_1_282
timestamp 1698175906
transform 1 0 16464 0 -1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_1_346
timestamp 1698175906
transform 1 0 20048 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_1_348
timestamp 1698175906
transform 1 0 20160 0 -1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_2
timestamp 1698175906
transform 1 0 784 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_2_34
timestamp 1698175906
transform 1 0 2576 0 1 2352
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_37
timestamp 1698175906
transform 1 0 2744 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_101
timestamp 1698175906
transform 1 0 6328 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_107
timestamp 1698175906
transform 1 0 6664 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_171
timestamp 1698175906
transform 1 0 10248 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_177 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 10584 0 1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_193
timestamp 1698175906
transform 1 0 11480 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_2_197
timestamp 1698175906
transform 1 0 11704 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_2_225
timestamp 1698175906
transform 1 0 13272 0 1 2352
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_241
timestamp 1698175906
transform 1 0 14168 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_2_247
timestamp 1698175906
transform 1 0 14504 0 1 2352
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_2_311
timestamp 1698175906
transform 1 0 18088 0 1 2352
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_2_317
timestamp 1698175906
transform 1 0 18424 0 1 2352
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_2
timestamp 1698175906
transform 1 0 784 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_66
timestamp 1698175906
transform 1 0 4368 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_72
timestamp 1698175906
transform 1 0 4704 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_136
timestamp 1698175906
transform 1 0 8288 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_142
timestamp 1698175906
transform 1 0 8624 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_206
timestamp 1698175906
transform 1 0 12208 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_212
timestamp 1698175906
transform 1 0 12544 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_3_276
timestamp 1698175906
transform 1 0 16128 0 -1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_3_282
timestamp 1698175906
transform 1 0 16464 0 -1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_3_346
timestamp 1698175906
transform 1 0 20048 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_3_348
timestamp 1698175906
transform 1 0 20160 0 -1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_2
timestamp 1698175906
transform 1 0 784 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_4_34
timestamp 1698175906
transform 1 0 2576 0 1 3136
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_37
timestamp 1698175906
transform 1 0 2744 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_101
timestamp 1698175906
transform 1 0 6328 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_107
timestamp 1698175906
transform 1 0 6664 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_171
timestamp 1698175906
transform 1 0 10248 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_177
timestamp 1698175906
transform 1 0 10584 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_241
timestamp 1698175906
transform 1 0 14168 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_4_247
timestamp 1698175906
transform 1 0 14504 0 1 3136
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_4_311
timestamp 1698175906
transform 1 0 18088 0 1 3136
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_4_317
timestamp 1698175906
transform 1 0 18424 0 1 3136
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_2
timestamp 1698175906
transform 1 0 784 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_66
timestamp 1698175906
transform 1 0 4368 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_72
timestamp 1698175906
transform 1 0 4704 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_136
timestamp 1698175906
transform 1 0 8288 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_142
timestamp 1698175906
transform 1 0 8624 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_206
timestamp 1698175906
transform 1 0 12208 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_212
timestamp 1698175906
transform 1 0 12544 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_5_276
timestamp 1698175906
transform 1 0 16128 0 -1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_5_282
timestamp 1698175906
transform 1 0 16464 0 -1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_5_346
timestamp 1698175906
transform 1 0 20048 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_5_348
timestamp 1698175906
transform 1 0 20160 0 -1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_2
timestamp 1698175906
transform 1 0 784 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_6_34
timestamp 1698175906
transform 1 0 2576 0 1 3920
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_37
timestamp 1698175906
transform 1 0 2744 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_101
timestamp 1698175906
transform 1 0 6328 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_107
timestamp 1698175906
transform 1 0 6664 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_171
timestamp 1698175906
transform 1 0 10248 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_177
timestamp 1698175906
transform 1 0 10584 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_241
timestamp 1698175906
transform 1 0 14168 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_6_247
timestamp 1698175906
transform 1 0 14504 0 1 3920
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_6_311
timestamp 1698175906
transform 1 0 18088 0 1 3920
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_6_317
timestamp 1698175906
transform 1 0 18424 0 1 3920
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_2
timestamp 1698175906
transform 1 0 784 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_66
timestamp 1698175906
transform 1 0 4368 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_72
timestamp 1698175906
transform 1 0 4704 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_136
timestamp 1698175906
transform 1 0 8288 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_142
timestamp 1698175906
transform 1 0 8624 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_206
timestamp 1698175906
transform 1 0 12208 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_212
timestamp 1698175906
transform 1 0 12544 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_7_276
timestamp 1698175906
transform 1 0 16128 0 -1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_7_282
timestamp 1698175906
transform 1 0 16464 0 -1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_7_346
timestamp 1698175906
transform 1 0 20048 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_7_348
timestamp 1698175906
transform 1 0 20160 0 -1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_2
timestamp 1698175906
transform 1 0 784 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_8_34
timestamp 1698175906
transform 1 0 2576 0 1 4704
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_37
timestamp 1698175906
transform 1 0 2744 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_101
timestamp 1698175906
transform 1 0 6328 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_107
timestamp 1698175906
transform 1 0 6664 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_171
timestamp 1698175906
transform 1 0 10248 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_177
timestamp 1698175906
transform 1 0 10584 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_241
timestamp 1698175906
transform 1 0 14168 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_8_247
timestamp 1698175906
transform 1 0 14504 0 1 4704
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_8_311
timestamp 1698175906
transform 1 0 18088 0 1 4704
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_8_317
timestamp 1698175906
transform 1 0 18424 0 1 4704
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_2
timestamp 1698175906
transform 1 0 784 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_66
timestamp 1698175906
transform 1 0 4368 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_72
timestamp 1698175906
transform 1 0 4704 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_136
timestamp 1698175906
transform 1 0 8288 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_142
timestamp 1698175906
transform 1 0 8624 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_206
timestamp 1698175906
transform 1 0 12208 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_212
timestamp 1698175906
transform 1 0 12544 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_9_276
timestamp 1698175906
transform 1 0 16128 0 -1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_9_282
timestamp 1698175906
transform 1 0 16464 0 -1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_9_346
timestamp 1698175906
transform 1 0 20048 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_9_348
timestamp 1698175906
transform 1 0 20160 0 -1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_2
timestamp 1698175906
transform 1 0 784 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_10_34
timestamp 1698175906
transform 1 0 2576 0 1 5488
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_37
timestamp 1698175906
transform 1 0 2744 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_101
timestamp 1698175906
transform 1 0 6328 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_107
timestamp 1698175906
transform 1 0 6664 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_171
timestamp 1698175906
transform 1 0 10248 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_177
timestamp 1698175906
transform 1 0 10584 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_241
timestamp 1698175906
transform 1 0 14168 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_10_247
timestamp 1698175906
transform 1 0 14504 0 1 5488
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_10_311
timestamp 1698175906
transform 1 0 18088 0 1 5488
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_10_317
timestamp 1698175906
transform 1 0 18424 0 1 5488
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_2
timestamp 1698175906
transform 1 0 784 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_66
timestamp 1698175906
transform 1 0 4368 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_72
timestamp 1698175906
transform 1 0 4704 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_136
timestamp 1698175906
transform 1 0 8288 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_142
timestamp 1698175906
transform 1 0 8624 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_206
timestamp 1698175906
transform 1 0 12208 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_212
timestamp 1698175906
transform 1 0 12544 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_11_276
timestamp 1698175906
transform 1 0 16128 0 -1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_11_282
timestamp 1698175906
transform 1 0 16464 0 -1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_11_346
timestamp 1698175906
transform 1 0 20048 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_11_348
timestamp 1698175906
transform 1 0 20160 0 -1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_2
timestamp 1698175906
transform 1 0 784 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_34
timestamp 1698175906
transform 1 0 2576 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_37
timestamp 1698175906
transform 1 0 2744 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_101
timestamp 1698175906
transform 1 0 6328 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_107
timestamp 1698175906
transform 1 0 6664 0 1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_123
timestamp 1698175906
transform 1 0 7560 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_12_154
timestamp 1698175906
transform 1 0 9296 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_12_158
timestamp 1698175906
transform 1 0 9520 0 1 6272
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_12_174
timestamp 1698175906
transform 1 0 10416 0 1 6272
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_177
timestamp 1698175906
transform 1 0 10584 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_241
timestamp 1698175906
transform 1 0 14168 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_12_247
timestamp 1698175906
transform 1 0 14504 0 1 6272
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_12_311
timestamp 1698175906
transform 1 0 18088 0 1 6272
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_12_317
timestamp 1698175906
transform 1 0 18424 0 1 6272
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_2
timestamp 1698175906
transform 1 0 784 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_66
timestamp 1698175906
transform 1 0 4368 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_72
timestamp 1698175906
transform 1 0 4704 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_136
timestamp 1698175906
transform 1 0 8288 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_13_142
timestamp 1698175906
transform 1 0 8624 0 -1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_13_174
timestamp 1698175906
transform 1 0 10416 0 -1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_178
timestamp 1698175906
transform 1 0 10640 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_180
timestamp 1698175906
transform 1 0 10752 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_212
timestamp 1698175906
transform 1 0 12544 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_216
timestamp 1698175906
transform 1 0 12768 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_13_282
timestamp 1698175906
transform 1 0 16464 0 -1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_13_346
timestamp 1698175906
transform 1 0 20048 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_13_348
timestamp 1698175906
transform 1 0 20160 0 -1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_2
timestamp 1698175906
transform 1 0 784 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_34
timestamp 1698175906
transform 1 0 2576 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_37
timestamp 1698175906
transform 1 0 2744 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_101
timestamp 1698175906
transform 1 0 6328 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_107
timestamp 1698175906
transform 1 0 6664 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_139
timestamp 1698175906
transform 1 0 8456 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_144
timestamp 1698175906
transform 1 0 8736 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_155
timestamp 1698175906
transform 1 0 9352 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_171
timestamp 1698175906
transform 1 0 10248 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_14_218
timestamp 1698175906
transform 1 0 12880 0 1 7056
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_14_234
timestamp 1698175906
transform 1 0 13776 0 1 7056
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_14_242
timestamp 1698175906
transform 1 0 14224 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_14_244
timestamp 1698175906
transform 1 0 14336 0 1 7056
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_14_247
timestamp 1698175906
transform 1 0 14504 0 1 7056
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_14_311
timestamp 1698175906
transform 1 0 18088 0 1 7056
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_14_317
timestamp 1698175906
transform 1 0 18424 0 1 7056
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_2
timestamp 1698175906
transform 1 0 784 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_66
timestamp 1698175906
transform 1 0 4368 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_72
timestamp 1698175906
transform 1 0 4704 0 -1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_104
timestamp 1698175906
transform 1 0 6496 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_108
timestamp 1698175906
transform 1 0 6720 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_110
timestamp 1698175906
transform 1 0 6832 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_171
timestamp 1698175906
transform 1 0 10248 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_175
timestamp 1698175906
transform 1 0 10472 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_183
timestamp 1698175906
transform 1 0 10920 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_187
timestamp 1698175906
transform 1 0 11144 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_200
timestamp 1698175906
transform 1 0 11872 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_204
timestamp 1698175906
transform 1 0 12096 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_208
timestamp 1698175906
transform 1 0 12320 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_15_212
timestamp 1698175906
transform 1 0 12544 0 -1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_15_234
timestamp 1698175906
transform 1 0 13776 0 -1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_15_266
timestamp 1698175906
transform 1 0 15568 0 -1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_15_274
timestamp 1698175906
transform 1 0 16016 0 -1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_278
timestamp 1698175906
transform 1 0 16240 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_15_282
timestamp 1698175906
transform 1 0 16464 0 -1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_15_346
timestamp 1698175906
transform 1 0 20048 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_15_348
timestamp 1698175906
transform 1 0 20160 0 -1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_16_2
timestamp 1698175906
transform 1 0 784 0 1 7840
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_34
timestamp 1698175906
transform 1 0 2576 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_37
timestamp 1698175906
transform 1 0 2744 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_101
timestamp 1698175906
transform 1 0 6328 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_16_107
timestamp 1698175906
transform 1 0 6664 0 1 7840
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_123
timestamp 1698175906
transform 1 0 7560 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_131
timestamp 1698175906
transform 1 0 8008 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_135
timestamp 1698175906
transform 1 0 8232 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_144
timestamp 1698175906
transform 1 0 8736 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_148
timestamp 1698175906
transform 1 0 8960 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_152
timestamp 1698175906
transform 1 0 9184 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_154
timestamp 1698175906
transform 1 0 9296 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_16_161
timestamp 1698175906
transform 1 0 9688 0 1 7840
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_169
timestamp 1698175906
transform 1 0 10136 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_173
timestamp 1698175906
transform 1 0 10360 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_177
timestamp 1698175906
transform 1 0 10584 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_195
timestamp 1698175906
transform 1 0 11592 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_199
timestamp 1698175906
transform 1 0 11816 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_210
timestamp 1698175906
transform 1 0 12432 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_242
timestamp 1698175906
transform 1 0 14224 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_16_244
timestamp 1698175906
transform 1 0 14336 0 1 7840
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_16_247
timestamp 1698175906
transform 1 0 14504 0 1 7840
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_311
timestamp 1698175906
transform 1 0 18088 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_16_317
timestamp 1698175906
transform 1 0 18424 0 1 7840
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_16_321
timestamp 1698175906
transform 1 0 18648 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_28
timestamp 1698175906
transform 1 0 2240 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_60
timestamp 1698175906
transform 1 0 4032 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_68
timestamp 1698175906
transform 1 0 4480 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_72
timestamp 1698175906
transform 1 0 4704 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_80
timestamp 1698175906
transform 1 0 5152 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_113
timestamp 1698175906
transform 1 0 7000 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_117
timestamp 1698175906
transform 1 0 7224 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_133
timestamp 1698175906
transform 1 0 8120 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_137
timestamp 1698175906
transform 1 0 8344 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_139
timestamp 1698175906
transform 1 0 8456 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_142
timestamp 1698175906
transform 1 0 8624 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_144
timestamp 1698175906
transform 1 0 8736 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_155
timestamp 1698175906
transform 1 0 9352 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_207
timestamp 1698175906
transform 1 0 12264 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_209
timestamp 1698175906
transform 1 0 12376 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_224
timestamp 1698175906
transform 1 0 13216 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_234
timestamp 1698175906
transform 1 0 13776 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_266
timestamp 1698175906
transform 1 0 15568 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_17_274
timestamp 1698175906
transform 1 0 16016 0 -1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_17_278
timestamp 1698175906
transform 1 0 16240 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_17_282
timestamp 1698175906
transform 1 0 16464 0 -1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_17_314
timestamp 1698175906
transform 1 0 18256 0 -1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_17_322
timestamp 1698175906
transform 1 0 18704 0 -1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_28
timestamp 1698175906
transform 1 0 2240 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_32
timestamp 1698175906
transform 1 0 2464 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_34
timestamp 1698175906
transform 1 0 2576 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_37
timestamp 1698175906
transform 1 0 2744 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_101
timestamp 1698175906
transform 1 0 6328 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_125
timestamp 1698175906
transform 1 0 7672 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_133
timestamp 1698175906
transform 1 0 8120 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_163
timestamp 1698175906
transform 1 0 9800 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_171
timestamp 1698175906
transform 1 0 10248 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_189
timestamp 1698175906
transform 1 0 11256 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_18_204
timestamp 1698175906
transform 1 0 12096 0 1 8624
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_18_236
timestamp 1698175906
transform 1 0 13888 0 1 8624
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_18_244
timestamp 1698175906
transform 1 0 14336 0 1 8624
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_18_247
timestamp 1698175906
transform 1 0 14504 0 1 8624
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_311
timestamp 1698175906
transform 1 0 18088 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_18_317
timestamp 1698175906
transform 1 0 18424 0 1 8624
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_18_321
timestamp 1698175906
transform 1 0 18648 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_2
timestamp 1698175906
transform 1 0 784 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_66
timestamp 1698175906
transform 1 0 4368 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_72
timestamp 1698175906
transform 1 0 4704 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_80
timestamp 1698175906
transform 1 0 5152 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_124
timestamp 1698175906
transform 1 0 7616 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_128
timestamp 1698175906
transform 1 0 7840 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_136
timestamp 1698175906
transform 1 0 8288 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_142
timestamp 1698175906
transform 1 0 8624 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_170
timestamp 1698175906
transform 1 0 10192 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_204
timestamp 1698175906
transform 1 0 12096 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_208
timestamp 1698175906
transform 1 0 12320 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_212
timestamp 1698175906
transform 1 0 12544 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_216
timestamp 1698175906
transform 1 0 12768 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_218
timestamp 1698175906
transform 1 0 12880 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_19_250
timestamp 1698175906
transform 1 0 14672 0 -1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_19_266
timestamp 1698175906
transform 1 0 15568 0 -1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_19_274
timestamp 1698175906
transform 1 0 16016 0 -1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_278
timestamp 1698175906
transform 1 0 16240 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_19_282
timestamp 1698175906
transform 1 0 16464 0 -1 9408
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_19_346
timestamp 1698175906
transform 1 0 20048 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_19_348
timestamp 1698175906
transform 1 0 20160 0 -1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_2
timestamp 1698175906
transform 1 0 784 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_34
timestamp 1698175906
transform 1 0 2576 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_37
timestamp 1698175906
transform 1 0 2744 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_69
timestamp 1698175906
transform 1 0 4536 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_73
timestamp 1698175906
transform 1 0 4760 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_75
timestamp 1698175906
transform 1 0 4872 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_107
timestamp 1698175906
transform 1 0 6664 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_121
timestamp 1698175906
transform 1 0 7448 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_125
timestamp 1698175906
transform 1 0 7672 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_138
timestamp 1698175906
transform 1 0 8400 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_140
timestamp 1698175906
transform 1 0 8512 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_167
timestamp 1698175906
transform 1 0 10024 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_189
timestamp 1698175906
transform 1 0 11256 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_205
timestamp 1698175906
transform 1 0 12152 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_221
timestamp 1698175906
transform 1 0 13048 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_223
timestamp 1698175906
transform 1 0 13160 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_242
timestamp 1698175906
transform 1 0 14224 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_244
timestamp 1698175906
transform 1 0 14336 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_20_252
timestamp 1698175906
transform 1 0 14784 0 1 9408
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_20_284
timestamp 1698175906
transform 1 0 16576 0 1 9408
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_20_300
timestamp 1698175906
transform 1 0 17472 0 1 9408
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_308
timestamp 1698175906
transform 1 0 17920 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_312
timestamp 1698175906
transform 1 0 18144 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_20_314
timestamp 1698175906
transform 1 0 18256 0 1 9408
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_20_317
timestamp 1698175906
transform 1 0 18424 0 1 9408
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_20_321
timestamp 1698175906
transform 1 0 18648 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_28
timestamp 1698175906
transform 1 0 2240 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_60
timestamp 1698175906
transform 1 0 4032 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_68
timestamp 1698175906
transform 1 0 4480 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_72
timestamp 1698175906
transform 1 0 4704 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_104
timestamp 1698175906
transform 1 0 6496 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_112
timestamp 1698175906
transform 1 0 6944 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_127
timestamp 1698175906
transform 1 0 7784 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_131
timestamp 1698175906
transform 1 0 8008 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_133
timestamp 1698175906
transform 1 0 8120 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_142
timestamp 1698175906
transform 1 0 8624 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_144
timestamp 1698175906
transform 1 0 8736 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_151
timestamp 1698175906
transform 1 0 9128 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_155
timestamp 1698175906
transform 1 0 9352 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_203
timestamp 1698175906
transform 1 0 12040 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_207
timestamp 1698175906
transform 1 0 12264 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_209
timestamp 1698175906
transform 1 0 12376 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_21_212
timestamp 1698175906
transform 1 0 12544 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_214
timestamp 1698175906
transform 1 0 12656 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_21_252
timestamp 1698175906
transform 1 0 14784 0 -1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_268
timestamp 1698175906
transform 1 0 15680 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_21_276
timestamp 1698175906
transform 1 0 16128 0 -1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_21_282
timestamp 1698175906
transform 1 0 16464 0 -1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_21_314
timestamp 1698175906
transform 1 0 18256 0 -1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_21_322
timestamp 1698175906
transform 1 0 18704 0 -1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_22_2
timestamp 1698175906
transform 1 0 784 0 1 10192
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_34
timestamp 1698175906
transform 1 0 2576 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_37
timestamp 1698175906
transform 1 0 2744 0 1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_101
timestamp 1698175906
transform 1 0 6328 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_107
timestamp 1698175906
transform 1 0 6664 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_115
timestamp 1698175906
transform 1 0 7112 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_121
timestamp 1698175906
transform 1 0 7448 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_137
timestamp 1698175906
transform 1 0 8344 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_158
timestamp 1698175906
transform 1 0 9520 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_162
timestamp 1698175906
transform 1 0 9744 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_170
timestamp 1698175906
transform 1 0 10192 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_174
timestamp 1698175906
transform 1 0 10416 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_177
timestamp 1698175906
transform 1 0 10584 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_193
timestamp 1698175906
transform 1 0 11480 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_22_203
timestamp 1698175906
transform 1 0 12040 0 1 10192
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_211
timestamp 1698175906
transform 1 0 12488 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_213
timestamp 1698175906
transform 1 0 12600 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_22_224
timestamp 1698175906
transform 1 0 13216 0 1 10192
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_240
timestamp 1698175906
transform 1 0 14112 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_22_244
timestamp 1698175906
transform 1 0 14336 0 1 10192
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_22_247
timestamp 1698175906
transform 1 0 14504 0 1 10192
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_311
timestamp 1698175906
transform 1 0 18088 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_22_317
timestamp 1698175906
transform 1 0 18424 0 1 10192
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_22_321
timestamp 1698175906
transform 1 0 18648 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_2
timestamp 1698175906
transform 1 0 784 0 -1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_66
timestamp 1698175906
transform 1 0 4368 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_72
timestamp 1698175906
transform 1 0 4704 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_88
timestamp 1698175906
transform 1 0 5600 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_131
timestamp 1698175906
transform 1 0 8008 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_133
timestamp 1698175906
transform 1 0 8120 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_150
timestamp 1698175906
transform 1 0 9072 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_154
timestamp 1698175906
transform 1 0 9296 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_156
timestamp 1698175906
transform 1 0 9408 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_209
timestamp 1698175906
transform 1 0 12376 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_23_217
timestamp 1698175906
transform 1 0 12824 0 -1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_221
timestamp 1698175906
transform 1 0 13048 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_23_254
timestamp 1698175906
transform 1 0 14896 0 -1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_23_270
timestamp 1698175906
transform 1 0 15792 0 -1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_278
timestamp 1698175906
transform 1 0 16240 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_23_282
timestamp 1698175906
transform 1 0 16464 0 -1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_23_346
timestamp 1698175906
transform 1 0 20048 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_23_348
timestamp 1698175906
transform 1 0 20160 0 -1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_24_2
timestamp 1698175906
transform 1 0 784 0 1 10976
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_34
timestamp 1698175906
transform 1 0 2576 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_37
timestamp 1698175906
transform 1 0 2744 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_101
timestamp 1698175906
transform 1 0 6328 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_24_107
timestamp 1698175906
transform 1 0 6664 0 1 10976
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_123
timestamp 1698175906
transform 1 0 7560 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_130
timestamp 1698175906
transform 1 0 7952 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_132
timestamp 1698175906
transform 1 0 8064 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_141
timestamp 1698175906
transform 1 0 8568 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_143
timestamp 1698175906
transform 1 0 8680 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_152
timestamp 1698175906
transform 1 0 9184 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_154
timestamp 1698175906
transform 1 0 9296 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_160
timestamp 1698175906
transform 1 0 9632 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_205
timestamp 1698175906
transform 1 0 12152 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_213
timestamp 1698175906
transform 1 0 12600 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_24_224
timestamp 1698175906
transform 1 0 13216 0 1 10976
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_232
timestamp 1698175906
transform 1 0 13664 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_24_234
timestamp 1698175906
transform 1 0 13776 0 1 10976
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_241
timestamp 1698175906
transform 1 0 14168 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_24_247
timestamp 1698175906
transform 1 0 14504 0 1 10976
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_311
timestamp 1698175906
transform 1 0 18088 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_24_317
timestamp 1698175906
transform 1 0 18424 0 1 10976
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_24_321
timestamp 1698175906
transform 1 0 18648 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_2
timestamp 1698175906
transform 1 0 784 0 -1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_66
timestamp 1698175906
transform 1 0 4368 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_72
timestamp 1698175906
transform 1 0 4704 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_80
timestamp 1698175906
transform 1 0 5152 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_84
timestamp 1698175906
transform 1 0 5376 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_114
timestamp 1698175906
transform 1 0 7056 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_118
timestamp 1698175906
transform 1 0 7280 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_126
timestamp 1698175906
transform 1 0 7728 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_135
timestamp 1698175906
transform 1 0 8232 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_139
timestamp 1698175906
transform 1 0 8456 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_142
timestamp 1698175906
transform 1 0 8624 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_151
timestamp 1698175906
transform 1 0 9128 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_212
timestamp 1698175906
transform 1 0 12544 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_216
timestamp 1698175906
transform 1 0 12768 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_224
timestamp 1698175906
transform 1 0 13216 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_228
timestamp 1698175906
transform 1 0 13440 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_25_236
timestamp 1698175906
transform 1 0 13888 0 -1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_25_268
timestamp 1698175906
transform 1 0 15680 0 -1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_25_276
timestamp 1698175906
transform 1 0 16128 0 -1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_25_282
timestamp 1698175906
transform 1 0 16464 0 -1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_25_346
timestamp 1698175906
transform 1 0 20048 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_25_348
timestamp 1698175906
transform 1 0 20160 0 -1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_28
timestamp 1698175906
transform 1 0 2240 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_32
timestamp 1698175906
transform 1 0 2464 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_34
timestamp 1698175906
transform 1 0 2576 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_37
timestamp 1698175906
transform 1 0 2744 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_101
timestamp 1698175906
transform 1 0 6328 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_148
timestamp 1698175906
transform 1 0 8960 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_156
timestamp 1698175906
transform 1 0 9408 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_164
timestamp 1698175906
transform 1 0 9856 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_170
timestamp 1698175906
transform 1 0 10192 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_174
timestamp 1698175906
transform 1 0 10416 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_177
timestamp 1698175906
transform 1 0 10584 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_183
timestamp 1698175906
transform 1 0 10920 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_26_215
timestamp 1698175906
transform 1 0 12712 0 1 11760
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_26_223
timestamp 1698175906
transform 1 0 13160 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_26_244
timestamp 1698175906
transform 1 0 14336 0 1 11760
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_26_247
timestamp 1698175906
transform 1 0 14504 0 1 11760
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_26_311
timestamp 1698175906
transform 1 0 18088 0 1 11760
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_26_317
timestamp 1698175906
transform 1 0 18424 0 1 11760
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_2
timestamp 1698175906
transform 1 0 784 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_66
timestamp 1698175906
transform 1 0 4368 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_27_72
timestamp 1698175906
transform 1 0 4704 0 -1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_104
timestamp 1698175906
transform 1 0 6496 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_120
timestamp 1698175906
transform 1 0 7392 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_128
timestamp 1698175906
transform 1 0 7840 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_130
timestamp 1698175906
transform 1 0 7952 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_139
timestamp 1698175906
transform 1 0 8456 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_142
timestamp 1698175906
transform 1 0 8624 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_27_146
timestamp 1698175906
transform 1 0 8848 0 -1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_154
timestamp 1698175906
transform 1 0 9296 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_206
timestamp 1698175906
transform 1 0 12208 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_212
timestamp 1698175906
transform 1 0 12544 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_224
timestamp 1698175906
transform 1 0 13216 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_27_257
timestamp 1698175906
transform 1 0 15064 0 -1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_27_273
timestamp 1698175906
transform 1 0 15960 0 -1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_277
timestamp 1698175906
transform 1 0 16184 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_279
timestamp 1698175906
transform 1 0 16296 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_27_282
timestamp 1698175906
transform 1 0 16464 0 -1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_27_346
timestamp 1698175906
transform 1 0 20048 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_27_348
timestamp 1698175906
transform 1 0 20160 0 -1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_2
timestamp 1698175906
transform 1 0 784 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_34
timestamp 1698175906
transform 1 0 2576 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_37
timestamp 1698175906
transform 1 0 2744 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_101
timestamp 1698175906
transform 1 0 6328 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_107
timestamp 1698175906
transform 1 0 6664 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_123
timestamp 1698175906
transform 1 0 7560 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_28_140
timestamp 1698175906
transform 1 0 8512 0 1 12544
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_156
timestamp 1698175906
transform 1 0 9408 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_164
timestamp 1698175906
transform 1 0 9856 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_168
timestamp 1698175906
transform 1 0 10080 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_177
timestamp 1698175906
transform 1 0 10584 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_28_185
timestamp 1698175906
transform 1 0 11032 0 1 12544
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_193
timestamp 1698175906
transform 1 0 11480 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_28_195
timestamp 1698175906
transform 1 0 11592 0 1 12544
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_204
timestamp 1698175906
transform 1 0 12096 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_28_208
timestamp 1698175906
transform 1 0 12320 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_241
timestamp 1698175906
transform 1 0 14168 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_28_247
timestamp 1698175906
transform 1 0 14504 0 1 12544
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_28_311
timestamp 1698175906
transform 1 0 18088 0 1 12544
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_28_317
timestamp 1698175906
transform 1 0 18424 0 1 12544
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_29_2
timestamp 1698175906
transform 1 0 784 0 -1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_66
timestamp 1698175906
transform 1 0 4368 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_72
timestamp 1698175906
transform 1 0 4704 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_88
timestamp 1698175906
transform 1 0 5600 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_96
timestamp 1698175906
transform 1 0 6048 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_98
timestamp 1698175906
transform 1 0 6160 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_128
timestamp 1698175906
transform 1 0 7840 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_147
timestamp 1698175906
transform 1 0 8904 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_168
timestamp 1698175906
transform 1 0 10080 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_217
timestamp 1698175906
transform 1 0 12824 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_221
timestamp 1698175906
transform 1 0 13048 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_225
timestamp 1698175906
transform 1 0 13272 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_227
timestamp 1698175906
transform 1 0 13384 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_233
timestamp 1698175906
transform 1 0 13720 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_241
timestamp 1698175906
transform 1 0 14168 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_29_249
timestamp 1698175906
transform 1 0 14616 0 -1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_265
timestamp 1698175906
transform 1 0 15512 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_29_273
timestamp 1698175906
transform 1 0 15960 0 -1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_29_277
timestamp 1698175906
transform 1 0 16184 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_279
timestamp 1698175906
transform 1 0 16296 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_29_282
timestamp 1698175906
transform 1 0 16464 0 -1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_29_314
timestamp 1698175906
transform 1 0 18256 0 -1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_29_322
timestamp 1698175906
transform 1 0 18704 0 -1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_28
timestamp 1698175906
transform 1 0 2240 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_32
timestamp 1698175906
transform 1 0 2464 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_34
timestamp 1698175906
transform 1 0 2576 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_37
timestamp 1698175906
transform 1 0 2744 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_101
timestamp 1698175906
transform 1 0 6328 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_107
timestamp 1698175906
transform 1 0 6664 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_157
timestamp 1698175906
transform 1 0 9464 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_161
timestamp 1698175906
transform 1 0 9688 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_174
timestamp 1698175906
transform 1 0 10416 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_30_182
timestamp 1698175906
transform 1 0 10864 0 1 13328
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_30_214
timestamp 1698175906
transform 1 0 12656 0 1 13328
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_30_230
timestamp 1698175906
transform 1 0 13552 0 1 13328
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_238
timestamp 1698175906
transform 1 0 14000 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_242
timestamp 1698175906
transform 1 0 14224 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_30_244
timestamp 1698175906
transform 1 0 14336 0 1 13328
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_30_247
timestamp 1698175906
transform 1 0 14504 0 1 13328
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_311
timestamp 1698175906
transform 1 0 18088 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_30_317
timestamp 1698175906
transform 1 0 18424 0 1 13328
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_30_321
timestamp 1698175906
transform 1 0 18648 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_2
timestamp 1698175906
transform 1 0 784 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_66
timestamp 1698175906
transform 1 0 4368 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_31_72
timestamp 1698175906
transform 1 0 4704 0 -1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_104
timestamp 1698175906
transform 1 0 6496 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_108
timestamp 1698175906
transform 1 0 6720 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_110
timestamp 1698175906
transform 1 0 6832 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_142
timestamp 1698175906
transform 1 0 8624 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_144
timestamp 1698175906
transform 1 0 8736 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_151
timestamp 1698175906
transform 1 0 9128 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_155
timestamp 1698175906
transform 1 0 9352 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_186
timestamp 1698175906
transform 1 0 11088 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_31_190
timestamp 1698175906
transform 1 0 11312 0 -1 14112
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_206
timestamp 1698175906
transform 1 0 12208 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_212
timestamp 1698175906
transform 1 0 12544 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_31_276
timestamp 1698175906
transform 1 0 16128 0 -1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_31_282
timestamp 1698175906
transform 1 0 16464 0 -1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_31_346
timestamp 1698175906
transform 1 0 20048 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_31_348
timestamp 1698175906
transform 1 0 20160 0 -1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_2
timestamp 1698175906
transform 1 0 784 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_34
timestamp 1698175906
transform 1 0 2576 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_37
timestamp 1698175906
transform 1 0 2744 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_101
timestamp 1698175906
transform 1 0 6328 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_107
timestamp 1698175906
transform 1 0 6664 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_139
timestamp 1698175906
transform 1 0 8456 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_142
timestamp 1698175906
transform 1 0 8624 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_32_174
timestamp 1698175906
transform 1 0 10416 0 1 14112
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_177
timestamp 1698175906
transform 1 0 10584 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_241
timestamp 1698175906
transform 1 0 14168 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_32_247
timestamp 1698175906
transform 1 0 14504 0 1 14112
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_32_311
timestamp 1698175906
transform 1 0 18088 0 1 14112
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_32_317
timestamp 1698175906
transform 1 0 18424 0 1 14112
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_2
timestamp 1698175906
transform 1 0 784 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_66
timestamp 1698175906
transform 1 0 4368 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_72
timestamp 1698175906
transform 1 0 4704 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_136
timestamp 1698175906
transform 1 0 8288 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_142
timestamp 1698175906
transform 1 0 8624 0 -1 14896
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_187
timestamp 1698175906
transform 1 0 11144 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_16  FILLER_0_33_191
timestamp 1698175906
transform 1 0 11368 0 -1 14896
box -43 -43 939 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_207
timestamp 1698175906
transform 1 0 12264 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_209
timestamp 1698175906
transform 1 0 12376 0 -1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_212
timestamp 1698175906
transform 1 0 12544 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_33_276
timestamp 1698175906
transform 1 0 16128 0 -1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_33_282
timestamp 1698175906
transform 1 0 16464 0 -1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_33_346
timestamp 1698175906
transform 1 0 20048 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_33_348
timestamp 1698175906
transform 1 0 20160 0 -1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_2
timestamp 1698175906
transform 1 0 784 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_34_34
timestamp 1698175906
transform 1 0 2576 0 1 14896
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_37
timestamp 1698175906
transform 1 0 2744 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_101
timestamp 1698175906
transform 1 0 6328 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_107
timestamp 1698175906
transform 1 0 6664 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_171
timestamp 1698175906
transform 1 0 10248 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_177
timestamp 1698175906
transform 1 0 10584 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_241
timestamp 1698175906
transform 1 0 14168 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_34_247
timestamp 1698175906
transform 1 0 14504 0 1 14896
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_34_311
timestamp 1698175906
transform 1 0 18088 0 1 14896
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_34_317
timestamp 1698175906
transform 1 0 18424 0 1 14896
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_2
timestamp 1698175906
transform 1 0 784 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_66
timestamp 1698175906
transform 1 0 4368 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_72
timestamp 1698175906
transform 1 0 4704 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_136
timestamp 1698175906
transform 1 0 8288 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_142
timestamp 1698175906
transform 1 0 8624 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_206
timestamp 1698175906
transform 1 0 12208 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_212
timestamp 1698175906
transform 1 0 12544 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_35_276
timestamp 1698175906
transform 1 0 16128 0 -1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_35_282
timestamp 1698175906
transform 1 0 16464 0 -1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_35_346
timestamp 1698175906
transform 1 0 20048 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_35_348
timestamp 1698175906
transform 1 0 20160 0 -1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_2
timestamp 1698175906
transform 1 0 784 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_36_34
timestamp 1698175906
transform 1 0 2576 0 1 15680
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_37
timestamp 1698175906
transform 1 0 2744 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_101
timestamp 1698175906
transform 1 0 6328 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_107
timestamp 1698175906
transform 1 0 6664 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_171
timestamp 1698175906
transform 1 0 10248 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_177
timestamp 1698175906
transform 1 0 10584 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_241
timestamp 1698175906
transform 1 0 14168 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_36_247
timestamp 1698175906
transform 1 0 14504 0 1 15680
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_36_311
timestamp 1698175906
transform 1 0 18088 0 1 15680
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_36_317
timestamp 1698175906
transform 1 0 18424 0 1 15680
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_2
timestamp 1698175906
transform 1 0 784 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_66
timestamp 1698175906
transform 1 0 4368 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_72
timestamp 1698175906
transform 1 0 4704 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_136
timestamp 1698175906
transform 1 0 8288 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_142
timestamp 1698175906
transform 1 0 8624 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_206
timestamp 1698175906
transform 1 0 12208 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_212
timestamp 1698175906
transform 1 0 12544 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_37_276
timestamp 1698175906
transform 1 0 16128 0 -1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_37_282
timestamp 1698175906
transform 1 0 16464 0 -1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_37_346
timestamp 1698175906
transform 1 0 20048 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_37_348
timestamp 1698175906
transform 1 0 20160 0 -1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_2
timestamp 1698175906
transform 1 0 784 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_38_34
timestamp 1698175906
transform 1 0 2576 0 1 16464
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_37
timestamp 1698175906
transform 1 0 2744 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_101
timestamp 1698175906
transform 1 0 6328 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_107
timestamp 1698175906
transform 1 0 6664 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_171
timestamp 1698175906
transform 1 0 10248 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_177
timestamp 1698175906
transform 1 0 10584 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_241
timestamp 1698175906
transform 1 0 14168 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_38_247
timestamp 1698175906
transform 1 0 14504 0 1 16464
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_38_311
timestamp 1698175906
transform 1 0 18088 0 1 16464
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_38_317
timestamp 1698175906
transform 1 0 18424 0 1 16464
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_2
timestamp 1698175906
transform 1 0 784 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_66
timestamp 1698175906
transform 1 0 4368 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_72
timestamp 1698175906
transform 1 0 4704 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_136
timestamp 1698175906
transform 1 0 8288 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_142
timestamp 1698175906
transform 1 0 8624 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_206
timestamp 1698175906
transform 1 0 12208 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_212
timestamp 1698175906
transform 1 0 12544 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_39_276
timestamp 1698175906
transform 1 0 16128 0 -1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_39_282
timestamp 1698175906
transform 1 0 16464 0 -1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_39_346
timestamp 1698175906
transform 1 0 20048 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_39_348
timestamp 1698175906
transform 1 0 20160 0 -1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_2
timestamp 1698175906
transform 1 0 784 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_40_34
timestamp 1698175906
transform 1 0 2576 0 1 17248
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_37
timestamp 1698175906
transform 1 0 2744 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_101
timestamp 1698175906
transform 1 0 6328 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_107
timestamp 1698175906
transform 1 0 6664 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_171
timestamp 1698175906
transform 1 0 10248 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_177
timestamp 1698175906
transform 1 0 10584 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_241
timestamp 1698175906
transform 1 0 14168 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_40_247
timestamp 1698175906
transform 1 0 14504 0 1 17248
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_40_311
timestamp 1698175906
transform 1 0 18088 0 1 17248
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_40_317
timestamp 1698175906
transform 1 0 18424 0 1 17248
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_2
timestamp 1698175906
transform 1 0 784 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_66
timestamp 1698175906
transform 1 0 4368 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_72
timestamp 1698175906
transform 1 0 4704 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_136
timestamp 1698175906
transform 1 0 8288 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_142
timestamp 1698175906
transform 1 0 8624 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_206
timestamp 1698175906
transform 1 0 12208 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_212
timestamp 1698175906
transform 1 0 12544 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_41_276
timestamp 1698175906
transform 1 0 16128 0 -1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_41_282
timestamp 1698175906
transform 1 0 16464 0 -1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_41_346
timestamp 1698175906
transform 1 0 20048 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_41_348
timestamp 1698175906
transform 1 0 20160 0 -1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_2
timestamp 1698175906
transform 1 0 784 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_42_34
timestamp 1698175906
transform 1 0 2576 0 1 18032
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_37
timestamp 1698175906
transform 1 0 2744 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_101
timestamp 1698175906
transform 1 0 6328 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_107
timestamp 1698175906
transform 1 0 6664 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_42_165
timestamp 1698175906
transform 1 0 9912 0 1 18032
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_42_173
timestamp 1698175906
transform 1 0 10360 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_177
timestamp 1698175906
transform 1 0 10584 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_241
timestamp 1698175906
transform 1 0 14168 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_42_247
timestamp 1698175906
transform 1 0 14504 0 1 18032
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_42_311
timestamp 1698175906
transform 1 0 18088 0 1 18032
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_42_317
timestamp 1698175906
transform 1 0 18424 0 1 18032
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_2
timestamp 1698175906
transform 1 0 784 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_66
timestamp 1698175906
transform 1 0 4368 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_72
timestamp 1698175906
transform 1 0 4704 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_136
timestamp 1698175906
transform 1 0 8288 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_142
timestamp 1698175906
transform 1 0 8624 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_144
timestamp 1698175906
transform 1 0 8736 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_8  FILLER_0_43_171
timestamp 1698175906
transform 1 0 10248 0 -1 18816
box -43 -43 491 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_179
timestamp 1698175906
transform 1 0 10696 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_207
timestamp 1698175906
transform 1 0 12264 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_209
timestamp 1698175906
transform 1 0 12376 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_212
timestamp 1698175906
transform 1 0 12544 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_43_276
timestamp 1698175906
transform 1 0 16128 0 -1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_64  FILLER_0_43_282
timestamp 1698175906
transform 1 0 16464 0 -1 18816
box -43 -43 3627 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_43_346
timestamp 1698175906
transform 1 0 20048 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_43_348
timestamp 1698175906
transform 1 0 20160 0 -1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_2
timestamp 1698175906
transform 1 0 784 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_36
timestamp 1698175906
transform 1 0 2688 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_70
timestamp 1698175906
transform 1 0 4592 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_104
timestamp 1698175906
transform 1 0 6496 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_138
timestamp 1698175906
transform 1 0 8400 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_142
timestamp 1698175906
transform 1 0 8624 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_172
timestamp 1698175906
transform 1 0 10304 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_176
timestamp 1698175906
transform 1 0 10528 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_206
timestamp 1698175906
transform 1 0 12208 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_210
timestamp 1698175906
transform 1 0 12432 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_237
timestamp 1698175906
transform 1 0 13944 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_240
timestamp 1698175906
transform 1 0 14112 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_274
timestamp 1698175906
transform 1 0 16016 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_32  FILLER_0_44_308
timestamp 1698175906
transform 1 0 17920 0 1 18816
box -43 -43 1835 435
use gf180mcu_fd_sc_mcu7t5v0__fillcap_4  FILLER_0_44_342
timestamp 1698175906
transform 1 0 19824 0 1 18816
box -43 -43 267 435
use gf180mcu_fd_sc_mcu7t5v0__fill_2  FILLER_0_44_346
timestamp 1698175906
transform 1 0 20048 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__fill_1  FILLER_0_44_348
timestamp 1698175906
transform 1 0 20160 0 1 18816
box -43 -43 99 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output1 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 8736 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output2
timestamp 1698175906
transform -1 0 2240 0 -1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output3
timestamp 1698175906
transform 1 0 18760 0 1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output4
timestamp 1698175906
transform -1 0 2240 0 1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output5
timestamp 1698175906
transform 1 0 10304 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output6
timestamp 1698175906
transform 1 0 18760 0 1 7840
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output7
timestamp 1698175906
transform 1 0 12208 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output8
timestamp 1698175906
transform 1 0 8792 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output9
timestamp 1698175906
transform 1 0 18760 0 1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output10
timestamp 1698175906
transform -1 0 13272 0 1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output11
timestamp 1698175906
transform -1 0 2240 0 -1 10192
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output12
timestamp 1698175906
transform -1 0 2240 0 1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output13
timestamp 1698175906
transform 1 0 18760 0 1 10192
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output14
timestamp 1698175906
transform 1 0 18760 0 -1 10192
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output15
timestamp 1698175906
transform 1 0 12544 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output16
timestamp 1698175906
transform 1 0 8624 0 -1 2352
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output17
timestamp 1698175906
transform 1 0 18760 0 1 10976
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output18
timestamp 1698175906
transform -1 0 9912 0 1 18032
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output19
timestamp 1698175906
transform 1 0 10808 0 -1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output20
timestamp 1698175906
transform 1 0 10640 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output21
timestamp 1698175906
transform 1 0 18760 0 -1 13328
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output22
timestamp 1698175906
transform 1 0 8736 0 1 1568
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output23
timestamp 1698175906
transform 1 0 18760 0 1 9408
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output24
timestamp 1698175906
transform 1 0 18760 0 -1 8624
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output25
timestamp 1698175906
transform 1 0 12488 0 1 18816
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__buf_8  output26
timestamp 1698175906
transform -1 0 2240 0 1 11760
box -43 -43 1499 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Left_45 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 672 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_0_Right_0
timestamp 1698175906
transform -1 0 20328 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Left_46
timestamp 1698175906
transform 1 0 672 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_1_Right_1
timestamp 1698175906
transform -1 0 20328 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Left_47
timestamp 1698175906
transform 1 0 672 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_2_Right_2
timestamp 1698175906
transform -1 0 20328 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Left_48
timestamp 1698175906
transform 1 0 672 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_3_Right_3
timestamp 1698175906
transform -1 0 20328 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Left_49
timestamp 1698175906
transform 1 0 672 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_4_Right_4
timestamp 1698175906
transform -1 0 20328 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Left_50
timestamp 1698175906
transform 1 0 672 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_5_Right_5
timestamp 1698175906
transform -1 0 20328 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Left_51
timestamp 1698175906
transform 1 0 672 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_6_Right_6
timestamp 1698175906
transform -1 0 20328 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Left_52
timestamp 1698175906
transform 1 0 672 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_7_Right_7
timestamp 1698175906
transform -1 0 20328 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Left_53
timestamp 1698175906
transform 1 0 672 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_8_Right_8
timestamp 1698175906
transform -1 0 20328 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Left_54
timestamp 1698175906
transform 1 0 672 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_9_Right_9
timestamp 1698175906
transform -1 0 20328 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Left_55
timestamp 1698175906
transform 1 0 672 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_10_Right_10
timestamp 1698175906
transform -1 0 20328 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Left_56
timestamp 1698175906
transform 1 0 672 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_11_Right_11
timestamp 1698175906
transform -1 0 20328 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Left_57
timestamp 1698175906
transform 1 0 672 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_12_Right_12
timestamp 1698175906
transform -1 0 20328 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Left_58
timestamp 1698175906
transform 1 0 672 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_13_Right_13
timestamp 1698175906
transform -1 0 20328 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Left_59
timestamp 1698175906
transform 1 0 672 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_14_Right_14
timestamp 1698175906
transform -1 0 20328 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Left_60
timestamp 1698175906
transform 1 0 672 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_15_Right_15
timestamp 1698175906
transform -1 0 20328 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Left_61
timestamp 1698175906
transform 1 0 672 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_16_Right_16
timestamp 1698175906
transform -1 0 20328 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Left_62
timestamp 1698175906
transform 1 0 672 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_17_Right_17
timestamp 1698175906
transform -1 0 20328 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Left_63
timestamp 1698175906
transform 1 0 672 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_18_Right_18
timestamp 1698175906
transform -1 0 20328 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Left_64
timestamp 1698175906
transform 1 0 672 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_19_Right_19
timestamp 1698175906
transform -1 0 20328 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Left_65
timestamp 1698175906
transform 1 0 672 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_20_Right_20
timestamp 1698175906
transform -1 0 20328 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Left_66
timestamp 1698175906
transform 1 0 672 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_21_Right_21
timestamp 1698175906
transform -1 0 20328 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Left_67
timestamp 1698175906
transform 1 0 672 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_22_Right_22
timestamp 1698175906
transform -1 0 20328 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Left_68
timestamp 1698175906
transform 1 0 672 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_23_Right_23
timestamp 1698175906
transform -1 0 20328 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Left_69
timestamp 1698175906
transform 1 0 672 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_24_Right_24
timestamp 1698175906
transform -1 0 20328 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Left_70
timestamp 1698175906
transform 1 0 672 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_25_Right_25
timestamp 1698175906
transform -1 0 20328 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Left_71
timestamp 1698175906
transform 1 0 672 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_26_Right_26
timestamp 1698175906
transform -1 0 20328 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Left_72
timestamp 1698175906
transform 1 0 672 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_27_Right_27
timestamp 1698175906
transform -1 0 20328 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Left_73
timestamp 1698175906
transform 1 0 672 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_28_Right_28
timestamp 1698175906
transform -1 0 20328 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Left_74
timestamp 1698175906
transform 1 0 672 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_29_Right_29
timestamp 1698175906
transform -1 0 20328 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Left_75
timestamp 1698175906
transform 1 0 672 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_30_Right_30
timestamp 1698175906
transform -1 0 20328 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Left_76
timestamp 1698175906
transform 1 0 672 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_31_Right_31
timestamp 1698175906
transform -1 0 20328 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Left_77
timestamp 1698175906
transform 1 0 672 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_32_Right_32
timestamp 1698175906
transform -1 0 20328 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Left_78
timestamp 1698175906
transform 1 0 672 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_33_Right_33
timestamp 1698175906
transform -1 0 20328 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Left_79
timestamp 1698175906
transform 1 0 672 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_34_Right_34
timestamp 1698175906
transform -1 0 20328 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Left_80
timestamp 1698175906
transform 1 0 672 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_35_Right_35
timestamp 1698175906
transform -1 0 20328 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Left_81
timestamp 1698175906
transform 1 0 672 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_36_Right_36
timestamp 1698175906
transform -1 0 20328 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Left_82
timestamp 1698175906
transform 1 0 672 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_37_Right_37
timestamp 1698175906
transform -1 0 20328 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Left_83
timestamp 1698175906
transform 1 0 672 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_38_Right_38
timestamp 1698175906
transform -1 0 20328 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Left_84
timestamp 1698175906
transform 1 0 672 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_39_Right_39
timestamp 1698175906
transform -1 0 20328 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Left_85
timestamp 1698175906
transform 1 0 672 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_40_Right_40
timestamp 1698175906
transform -1 0 20328 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Left_86
timestamp 1698175906
transform 1 0 672 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_41_Right_41
timestamp 1698175906
transform -1 0 20328 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Left_87
timestamp 1698175906
transform 1 0 672 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_42_Right_42
timestamp 1698175906
transform -1 0 20328 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Left_88
timestamp 1698175906
transform 1 0 672 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_43_Right_43
timestamp 1698175906
transform -1 0 20328 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Left_89
timestamp 1698175906
transform 1 0 672 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__endcap  PHY_EDGE_ROW_44_Right_44
timestamp 1698175906
transform -1 0 20328 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_90 dependencies/pdks/gf180mcuD/libs.ref/gf180mcu_fd_sc_mcu7t5v0/mag
timestamp 1698175906
transform 1 0 2576 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_91
timestamp 1698175906
transform 1 0 4480 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_92
timestamp 1698175906
transform 1 0 6384 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_93
timestamp 1698175906
transform 1 0 8288 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_94
timestamp 1698175906
transform 1 0 10192 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_95
timestamp 1698175906
transform 1 0 12096 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_96
timestamp 1698175906
transform 1 0 14000 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_97
timestamp 1698175906
transform 1 0 15904 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_98
timestamp 1698175906
transform 1 0 17808 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_0_99
timestamp 1698175906
transform 1 0 19712 0 1 1568
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_100
timestamp 1698175906
transform 1 0 4592 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_101
timestamp 1698175906
transform 1 0 8512 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_102
timestamp 1698175906
transform 1 0 12432 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_1_103
timestamp 1698175906
transform 1 0 16352 0 -1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_104
timestamp 1698175906
transform 1 0 2632 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_105
timestamp 1698175906
transform 1 0 6552 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_106
timestamp 1698175906
transform 1 0 10472 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_107
timestamp 1698175906
transform 1 0 14392 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_2_108
timestamp 1698175906
transform 1 0 18312 0 1 2352
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_109
timestamp 1698175906
transform 1 0 4592 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_110
timestamp 1698175906
transform 1 0 8512 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_111
timestamp 1698175906
transform 1 0 12432 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_3_112
timestamp 1698175906
transform 1 0 16352 0 -1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_113
timestamp 1698175906
transform 1 0 2632 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_114
timestamp 1698175906
transform 1 0 6552 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_115
timestamp 1698175906
transform 1 0 10472 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_116
timestamp 1698175906
transform 1 0 14392 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_4_117
timestamp 1698175906
transform 1 0 18312 0 1 3136
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_118
timestamp 1698175906
transform 1 0 4592 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_119
timestamp 1698175906
transform 1 0 8512 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_120
timestamp 1698175906
transform 1 0 12432 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_5_121
timestamp 1698175906
transform 1 0 16352 0 -1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_122
timestamp 1698175906
transform 1 0 2632 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_123
timestamp 1698175906
transform 1 0 6552 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_124
timestamp 1698175906
transform 1 0 10472 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_125
timestamp 1698175906
transform 1 0 14392 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_6_126
timestamp 1698175906
transform 1 0 18312 0 1 3920
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_127
timestamp 1698175906
transform 1 0 4592 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_128
timestamp 1698175906
transform 1 0 8512 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_129
timestamp 1698175906
transform 1 0 12432 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_7_130
timestamp 1698175906
transform 1 0 16352 0 -1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_131
timestamp 1698175906
transform 1 0 2632 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_132
timestamp 1698175906
transform 1 0 6552 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_133
timestamp 1698175906
transform 1 0 10472 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_134
timestamp 1698175906
transform 1 0 14392 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_8_135
timestamp 1698175906
transform 1 0 18312 0 1 4704
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_136
timestamp 1698175906
transform 1 0 4592 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_137
timestamp 1698175906
transform 1 0 8512 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_138
timestamp 1698175906
transform 1 0 12432 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_9_139
timestamp 1698175906
transform 1 0 16352 0 -1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_140
timestamp 1698175906
transform 1 0 2632 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_141
timestamp 1698175906
transform 1 0 6552 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_142
timestamp 1698175906
transform 1 0 10472 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_143
timestamp 1698175906
transform 1 0 14392 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_10_144
timestamp 1698175906
transform 1 0 18312 0 1 5488
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_145
timestamp 1698175906
transform 1 0 4592 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_146
timestamp 1698175906
transform 1 0 8512 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_147
timestamp 1698175906
transform 1 0 12432 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_11_148
timestamp 1698175906
transform 1 0 16352 0 -1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_149
timestamp 1698175906
transform 1 0 2632 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_150
timestamp 1698175906
transform 1 0 6552 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_151
timestamp 1698175906
transform 1 0 10472 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_152
timestamp 1698175906
transform 1 0 14392 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_12_153
timestamp 1698175906
transform 1 0 18312 0 1 6272
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_154
timestamp 1698175906
transform 1 0 4592 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_155
timestamp 1698175906
transform 1 0 8512 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_156
timestamp 1698175906
transform 1 0 12432 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_13_157
timestamp 1698175906
transform 1 0 16352 0 -1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_158
timestamp 1698175906
transform 1 0 2632 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_159
timestamp 1698175906
transform 1 0 6552 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_160
timestamp 1698175906
transform 1 0 10472 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_161
timestamp 1698175906
transform 1 0 14392 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_14_162
timestamp 1698175906
transform 1 0 18312 0 1 7056
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_163
timestamp 1698175906
transform 1 0 4592 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_164
timestamp 1698175906
transform 1 0 8512 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_165
timestamp 1698175906
transform 1 0 12432 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_15_166
timestamp 1698175906
transform 1 0 16352 0 -1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_167
timestamp 1698175906
transform 1 0 2632 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_168
timestamp 1698175906
transform 1 0 6552 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_169
timestamp 1698175906
transform 1 0 10472 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_170
timestamp 1698175906
transform 1 0 14392 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_16_171
timestamp 1698175906
transform 1 0 18312 0 1 7840
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_172
timestamp 1698175906
transform 1 0 4592 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_173
timestamp 1698175906
transform 1 0 8512 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_174
timestamp 1698175906
transform 1 0 12432 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_17_175
timestamp 1698175906
transform 1 0 16352 0 -1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_176
timestamp 1698175906
transform 1 0 2632 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_177
timestamp 1698175906
transform 1 0 6552 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_178
timestamp 1698175906
transform 1 0 10472 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_179
timestamp 1698175906
transform 1 0 14392 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_18_180
timestamp 1698175906
transform 1 0 18312 0 1 8624
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_181
timestamp 1698175906
transform 1 0 4592 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_182
timestamp 1698175906
transform 1 0 8512 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_183
timestamp 1698175906
transform 1 0 12432 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_19_184
timestamp 1698175906
transform 1 0 16352 0 -1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_185
timestamp 1698175906
transform 1 0 2632 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_186
timestamp 1698175906
transform 1 0 6552 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_187
timestamp 1698175906
transform 1 0 10472 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_188
timestamp 1698175906
transform 1 0 14392 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_20_189
timestamp 1698175906
transform 1 0 18312 0 1 9408
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_190
timestamp 1698175906
transform 1 0 4592 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_191
timestamp 1698175906
transform 1 0 8512 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_192
timestamp 1698175906
transform 1 0 12432 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_21_193
timestamp 1698175906
transform 1 0 16352 0 -1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_194
timestamp 1698175906
transform 1 0 2632 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_195
timestamp 1698175906
transform 1 0 6552 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_196
timestamp 1698175906
transform 1 0 10472 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_197
timestamp 1698175906
transform 1 0 14392 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_22_198
timestamp 1698175906
transform 1 0 18312 0 1 10192
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_199
timestamp 1698175906
transform 1 0 4592 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_200
timestamp 1698175906
transform 1 0 8512 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_201
timestamp 1698175906
transform 1 0 12432 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_23_202
timestamp 1698175906
transform 1 0 16352 0 -1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_203
timestamp 1698175906
transform 1 0 2632 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_204
timestamp 1698175906
transform 1 0 6552 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_205
timestamp 1698175906
transform 1 0 10472 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_206
timestamp 1698175906
transform 1 0 14392 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_24_207
timestamp 1698175906
transform 1 0 18312 0 1 10976
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_208
timestamp 1698175906
transform 1 0 4592 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_209
timestamp 1698175906
transform 1 0 8512 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_210
timestamp 1698175906
transform 1 0 12432 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_25_211
timestamp 1698175906
transform 1 0 16352 0 -1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_212
timestamp 1698175906
transform 1 0 2632 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_213
timestamp 1698175906
transform 1 0 6552 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_214
timestamp 1698175906
transform 1 0 10472 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_215
timestamp 1698175906
transform 1 0 14392 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_26_216
timestamp 1698175906
transform 1 0 18312 0 1 11760
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_217
timestamp 1698175906
transform 1 0 4592 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_218
timestamp 1698175906
transform 1 0 8512 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_219
timestamp 1698175906
transform 1 0 12432 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_27_220
timestamp 1698175906
transform 1 0 16352 0 -1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_221
timestamp 1698175906
transform 1 0 2632 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_222
timestamp 1698175906
transform 1 0 6552 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_223
timestamp 1698175906
transform 1 0 10472 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_224
timestamp 1698175906
transform 1 0 14392 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_28_225
timestamp 1698175906
transform 1 0 18312 0 1 12544
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_226
timestamp 1698175906
transform 1 0 4592 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_227
timestamp 1698175906
transform 1 0 8512 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_228
timestamp 1698175906
transform 1 0 12432 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_29_229
timestamp 1698175906
transform 1 0 16352 0 -1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_230
timestamp 1698175906
transform 1 0 2632 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_231
timestamp 1698175906
transform 1 0 6552 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_232
timestamp 1698175906
transform 1 0 10472 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_233
timestamp 1698175906
transform 1 0 14392 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_30_234
timestamp 1698175906
transform 1 0 18312 0 1 13328
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_235
timestamp 1698175906
transform 1 0 4592 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_236
timestamp 1698175906
transform 1 0 8512 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_237
timestamp 1698175906
transform 1 0 12432 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_31_238
timestamp 1698175906
transform 1 0 16352 0 -1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_239
timestamp 1698175906
transform 1 0 2632 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_240
timestamp 1698175906
transform 1 0 6552 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_241
timestamp 1698175906
transform 1 0 10472 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_242
timestamp 1698175906
transform 1 0 14392 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_32_243
timestamp 1698175906
transform 1 0 18312 0 1 14112
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_244
timestamp 1698175906
transform 1 0 4592 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_245
timestamp 1698175906
transform 1 0 8512 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_246
timestamp 1698175906
transform 1 0 12432 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_33_247
timestamp 1698175906
transform 1 0 16352 0 -1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_248
timestamp 1698175906
transform 1 0 2632 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_249
timestamp 1698175906
transform 1 0 6552 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_250
timestamp 1698175906
transform 1 0 10472 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_251
timestamp 1698175906
transform 1 0 14392 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_34_252
timestamp 1698175906
transform 1 0 18312 0 1 14896
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_253
timestamp 1698175906
transform 1 0 4592 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_254
timestamp 1698175906
transform 1 0 8512 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_255
timestamp 1698175906
transform 1 0 12432 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_35_256
timestamp 1698175906
transform 1 0 16352 0 -1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_257
timestamp 1698175906
transform 1 0 2632 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_258
timestamp 1698175906
transform 1 0 6552 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_259
timestamp 1698175906
transform 1 0 10472 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_260
timestamp 1698175906
transform 1 0 14392 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_36_261
timestamp 1698175906
transform 1 0 18312 0 1 15680
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_262
timestamp 1698175906
transform 1 0 4592 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_263
timestamp 1698175906
transform 1 0 8512 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_264
timestamp 1698175906
transform 1 0 12432 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_37_265
timestamp 1698175906
transform 1 0 16352 0 -1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_266
timestamp 1698175906
transform 1 0 2632 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_267
timestamp 1698175906
transform 1 0 6552 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_268
timestamp 1698175906
transform 1 0 10472 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_269
timestamp 1698175906
transform 1 0 14392 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_38_270
timestamp 1698175906
transform 1 0 18312 0 1 16464
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_271
timestamp 1698175906
transform 1 0 4592 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_272
timestamp 1698175906
transform 1 0 8512 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_273
timestamp 1698175906
transform 1 0 12432 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_39_274
timestamp 1698175906
transform 1 0 16352 0 -1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_275
timestamp 1698175906
transform 1 0 2632 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_276
timestamp 1698175906
transform 1 0 6552 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_277
timestamp 1698175906
transform 1 0 10472 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_278
timestamp 1698175906
transform 1 0 14392 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_40_279
timestamp 1698175906
transform 1 0 18312 0 1 17248
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_280
timestamp 1698175906
transform 1 0 4592 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_281
timestamp 1698175906
transform 1 0 8512 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_282
timestamp 1698175906
transform 1 0 12432 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_41_283
timestamp 1698175906
transform 1 0 16352 0 -1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_284
timestamp 1698175906
transform 1 0 2632 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_285
timestamp 1698175906
transform 1 0 6552 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_286
timestamp 1698175906
transform 1 0 10472 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_287
timestamp 1698175906
transform 1 0 14392 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_42_288
timestamp 1698175906
transform 1 0 18312 0 1 18032
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_289
timestamp 1698175906
transform 1 0 4592 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_290
timestamp 1698175906
transform 1 0 8512 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_291
timestamp 1698175906
transform 1 0 12432 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_43_292
timestamp 1698175906
transform 1 0 16352 0 -1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_293
timestamp 1698175906
transform 1 0 2576 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_294
timestamp 1698175906
transform 1 0 4480 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_295
timestamp 1698175906
transform 1 0 6384 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_296
timestamp 1698175906
transform 1 0 8288 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_297
timestamp 1698175906
transform 1 0 10192 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_298
timestamp 1698175906
transform 1 0 12096 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_299
timestamp 1698175906
transform 1 0 14000 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_300
timestamp 1698175906
transform 1 0 15904 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_301
timestamp 1698175906
transform 1 0 17808 0 1 18816
box -43 -43 155 435
use gf180mcu_fd_sc_mcu7t5v0__filltie  TAP_TAPCELL_ROW_44_302
timestamp 1698175906
transform 1 0 19712 0 1 18816
box -43 -43 155 435
<< labels >>
flabel metal3 s 0 13776 400 13832 0 FreeSans 224 0 0 0 clk
port 0 nsew signal input
flabel metal2 s 9072 20600 9128 21000 0 FreeSans 224 90 0 0 segm[0]
port 1 nsew signal tristate
flabel metal3 s 0 8400 400 8456 0 FreeSans 224 0 0 0 segm[10]
port 2 nsew signal tristate
flabel metal3 s 20600 13104 21000 13160 0 FreeSans 224 0 0 0 segm[11]
port 3 nsew signal tristate
flabel metal3 s 0 8736 400 8792 0 FreeSans 224 0 0 0 segm[12]
port 4 nsew signal tristate
flabel metal2 s 9744 0 9800 400 0 FreeSans 224 90 0 0 segm[13]
port 5 nsew signal tristate
flabel metal3 s 20600 7728 21000 7784 0 FreeSans 224 0 0 0 segm[1]
port 6 nsew signal tristate
flabel metal2 s 11424 0 11480 400 0 FreeSans 224 90 0 0 segm[2]
port 7 nsew signal tristate
flabel metal2 s 8736 20600 8792 21000 0 FreeSans 224 90 0 0 segm[3]
port 8 nsew signal tristate
flabel metal3 s 20600 8400 21000 8456 0 FreeSans 224 0 0 0 segm[4]
port 9 nsew signal tristate
flabel metal2 s 11760 0 11816 400 0 FreeSans 224 90 0 0 segm[5]
port 10 nsew signal tristate
flabel metal3 s 0 9744 400 9800 0 FreeSans 224 0 0 0 segm[6]
port 11 nsew signal tristate
flabel metal3 s 0 13104 400 13160 0 FreeSans 224 0 0 0 segm[7]
port 12 nsew signal tristate
flabel metal3 s 20600 10080 21000 10136 0 FreeSans 224 0 0 0 segm[8]
port 13 nsew signal tristate
flabel metal3 s 20600 9744 21000 9800 0 FreeSans 224 0 0 0 segm[9]
port 14 nsew signal tristate
flabel metal2 s 12432 0 12488 400 0 FreeSans 224 90 0 0 sel[0]
port 15 nsew signal tristate
flabel metal2 s 8400 0 8456 400 0 FreeSans 224 90 0 0 sel[10]
port 16 nsew signal tristate
flabel metal3 s 20600 11088 21000 11144 0 FreeSans 224 0 0 0 sel[11]
port 17 nsew signal tristate
flabel metal2 s 8400 20600 8456 21000 0 FreeSans 224 90 0 0 sel[1]
port 18 nsew signal tristate
flabel metal2 s 10752 20600 10808 21000 0 FreeSans 224 90 0 0 sel[2]
port 19 nsew signal tristate
flabel metal2 s 11088 20600 11144 21000 0 FreeSans 224 90 0 0 sel[3]
port 20 nsew signal tristate
flabel metal3 s 20600 12768 21000 12824 0 FreeSans 224 0 0 0 sel[4]
port 21 nsew signal tristate
flabel metal2 s 9072 0 9128 400 0 FreeSans 224 90 0 0 sel[5]
port 22 nsew signal tristate
flabel metal3 s 20600 9408 21000 9464 0 FreeSans 224 0 0 0 sel[6]
port 23 nsew signal tristate
flabel metal3 s 20600 8064 21000 8120 0 FreeSans 224 0 0 0 sel[7]
port 24 nsew signal tristate
flabel metal2 s 12432 20600 12488 21000 0 FreeSans 224 90 0 0 sel[8]
port 25 nsew signal tristate
flabel metal3 s 0 11760 400 11816 0 FreeSans 224 0 0 0 sel[9]
port 26 nsew signal tristate
flabel metal4 s 2224 1538 2384 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 17584 1538 17744 19238 0 FreeSans 640 90 0 0 vdd
port 27 nsew power bidirectional
flabel metal4 s 9904 1538 10064 19238 0 FreeSans 640 90 0 0 vss
port 28 nsew ground bidirectional
rlabel metal1 10500 19208 10500 19208 0 vdd
rlabel metal1 10500 18816 10500 18816 0 vss
rlabel metal2 11788 12936 11788 12936 0 _000_
rlabel metal3 8148 11900 8148 11900 0 _001_
rlabel metal2 13524 9296 13524 9296 0 _002_
rlabel metal2 8596 11788 8596 11788 0 _003_
rlabel metal2 6860 10528 6860 10528 0 _004_
rlabel metal2 10892 11368 10892 11368 0 _005_
rlabel metal2 11508 11368 11508 11368 0 _006_
rlabel metal2 8148 6832 8148 6832 0 _007_
rlabel metal2 12964 12460 12964 12460 0 _008_
rlabel metal2 10164 13860 10164 13860 0 _009_
rlabel metal2 9884 13860 9884 13860 0 _010_
rlabel metal2 7364 13552 7364 13552 0 _011_
rlabel metal2 11284 7056 11284 7056 0 _012_
rlabel metal2 6076 9800 6076 9800 0 _013_
rlabel metal2 6524 9268 6524 9268 0 _014_
rlabel metal2 6524 8596 6524 8596 0 _015_
rlabel metal2 8148 13468 8148 13468 0 _016_
rlabel metal2 7364 12964 7364 12964 0 _017_
rlabel metal2 9128 7700 9128 7700 0 _018_
rlabel metal2 12992 7980 12992 7980 0 _019_
rlabel metal2 13300 10248 13300 10248 0 _020_
rlabel metal2 7364 8036 7364 8036 0 _021_
rlabel metal2 13748 11172 13748 11172 0 _022_
rlabel metal2 11088 7308 11088 7308 0 _023_
rlabel metal2 13972 11844 13972 11844 0 _024_
rlabel metal2 13188 12684 13188 12684 0 _025_
rlabel metal3 10024 13468 10024 13468 0 _026_
rlabel metal2 10528 13636 10528 13636 0 _027_
rlabel metal3 10248 13188 10248 13188 0 _028_
rlabel metal2 9156 12572 9156 12572 0 _029_
rlabel metal3 8568 11732 8568 11732 0 _030_
rlabel metal3 8680 13468 8680 13468 0 _031_
rlabel metal2 12068 7644 12068 7644 0 _032_
rlabel metal2 11452 8344 11452 8344 0 _033_
rlabel metal2 10724 8316 10724 8316 0 _034_
rlabel metal2 11536 7980 11536 7980 0 _035_
rlabel metal2 7420 9100 7420 9100 0 _036_
rlabel metal2 7308 9856 7308 9856 0 _037_
rlabel metal2 10948 8372 10948 8372 0 _038_
rlabel metal2 7476 9996 7476 9996 0 _039_
rlabel metal2 7532 9072 7532 9072 0 _040_
rlabel metal2 9016 8932 9016 8932 0 _041_
rlabel metal2 8876 9044 8876 9044 0 _042_
rlabel metal2 7308 9240 7308 9240 0 _043_
rlabel metal2 7252 8848 7252 8848 0 _044_
rlabel metal3 6972 8932 6972 8932 0 _045_
rlabel metal2 7000 8820 7000 8820 0 _046_
rlabel metal2 8540 13132 8540 13132 0 _047_
rlabel metal3 8064 12740 8064 12740 0 _048_
rlabel metal2 8372 12600 8372 12600 0 _049_
rlabel metal2 9436 8260 9436 8260 0 _050_
rlabel metal2 12180 8260 12180 8260 0 _051_
rlabel metal2 12348 8288 12348 8288 0 _052_
rlabel metal2 12796 10920 12796 10920 0 _053_
rlabel metal2 13132 10024 13132 10024 0 _054_
rlabel metal2 8428 8120 8428 8120 0 _055_
rlabel metal2 13636 11368 13636 11368 0 _056_
rlabel metal2 13972 11340 13972 11340 0 _057_
rlabel metal2 11340 7840 11340 7840 0 _058_
rlabel metal2 12908 11592 12908 11592 0 _059_
rlabel metal2 14476 12852 14476 12852 0 _060_
rlabel metal2 13748 11900 13748 11900 0 _061_
rlabel metal2 14056 11956 14056 11956 0 _062_
rlabel metal3 11480 9492 11480 9492 0 _063_
rlabel via2 11004 9156 11004 9156 0 _064_
rlabel metal2 9940 10640 9940 10640 0 _065_
rlabel metal2 9436 11396 9436 11396 0 _066_
rlabel metal3 10360 12068 10360 12068 0 _067_
rlabel metal2 11900 10528 11900 10528 0 _068_
rlabel metal2 11788 9940 11788 9940 0 _069_
rlabel metal2 11620 9296 11620 9296 0 _070_
rlabel metal3 11340 9996 11340 9996 0 _071_
rlabel metal2 10780 11144 10780 11144 0 _072_
rlabel metal2 13524 12964 13524 12964 0 _073_
rlabel metal2 12068 12880 12068 12880 0 _074_
rlabel metal2 8428 10472 8428 10472 0 _075_
rlabel metal2 9492 9772 9492 9772 0 _076_
rlabel metal2 9828 9912 9828 9912 0 _077_
rlabel metal2 7868 11144 7868 11144 0 _078_
rlabel metal2 9716 8764 9716 8764 0 _079_
rlabel metal2 9044 11872 9044 11872 0 _080_
rlabel metal3 8736 11844 8736 11844 0 _081_
rlabel metal2 11116 9100 11116 9100 0 _082_
rlabel metal2 8316 9632 8316 9632 0 _083_
rlabel metal2 7364 9128 7364 9128 0 _084_
rlabel metal2 8120 11452 8120 11452 0 _085_
rlabel metal2 14588 9520 14588 9520 0 _086_
rlabel metal3 14392 9548 14392 9548 0 _087_
rlabel metal3 10080 10052 10080 10052 0 _088_
rlabel metal2 7196 9940 7196 9940 0 _089_
rlabel metal2 14084 9828 14084 9828 0 _090_
rlabel metal2 7028 10444 7028 10444 0 _091_
rlabel metal3 9436 11060 9436 11060 0 _092_
rlabel metal2 9940 11396 9940 11396 0 _093_
rlabel metal2 11396 10080 11396 10080 0 _094_
rlabel metal2 7112 9604 7112 9604 0 _095_
rlabel metal2 10220 11956 10220 11956 0 _096_
rlabel metal2 12740 11760 12740 11760 0 _097_
rlabel metal2 11732 11032 11732 11032 0 _098_
rlabel metal3 11788 7364 11788 7364 0 _099_
rlabel metal2 9296 8820 9296 8820 0 _100_
rlabel metal2 9100 8568 9100 8568 0 _101_
rlabel metal2 8932 7364 8932 7364 0 _102_
rlabel metal2 8764 7308 8764 7308 0 _103_
rlabel metal3 1239 13804 1239 13804 0 clk
rlabel metal2 10948 10612 10948 10612 0 clknet_0_clk
rlabel metal2 10892 7056 10892 7056 0 clknet_1_0__leaf_clk
rlabel metal2 11228 14140 11228 14140 0 clknet_1_1__leaf_clk
rlabel metal2 7532 11200 7532 11200 0 dut15.count\[0\]
rlabel metal2 7252 10808 7252 10808 0 dut15.count\[1\]
rlabel metal3 10920 10388 10920 10388 0 dut15.count\[2\]
rlabel metal2 12068 11340 12068 11340 0 dut15.count\[3\]
rlabel metal2 8876 14994 8876 14994 0 net1
rlabel metal2 12348 6776 12348 6776 0 net10
rlabel metal2 5012 9604 5012 9604 0 net11
rlabel metal2 6300 13300 6300 13300 0 net12
rlabel metal3 16828 10052 16828 10052 0 net13
rlabel metal2 14364 9968 14364 9968 0 net14
rlabel metal2 12628 3178 12628 3178 0 net15
rlabel metal2 8708 3178 8708 3178 0 net16
rlabel metal2 14812 10948 14812 10948 0 net17
rlabel metal2 9296 13468 9296 13468 0 net18
rlabel metal2 11004 16240 11004 16240 0 net19
rlabel metal2 5432 9156 5432 9156 0 net2
rlabel metal3 10892 14644 10892 14644 0 net20
rlabel metal2 13608 13188 13608 13188 0 net21
rlabel metal2 8820 2982 8820 2982 0 net22
rlabel metal2 14588 9212 14588 9212 0 net23
rlabel metal2 13692 8428 13692 8428 0 net24
rlabel metal3 12516 13188 12516 13188 0 net25
rlabel metal2 6748 11984 6748 11984 0 net26
rlabel metal2 14980 12684 14980 12684 0 net3
rlabel metal2 5460 8596 5460 8596 0 net4
rlabel metal2 10388 2982 10388 2982 0 net5
rlabel metal2 18844 7868 18844 7868 0 net6
rlabel metal2 12292 2982 12292 2982 0 net7
rlabel metal2 9100 13804 9100 13804 0 net8
rlabel metal2 14084 8260 14084 8260 0 net9
rlabel metal2 9100 19873 9100 19873 0 segm[0]
rlabel metal3 679 8428 679 8428 0 segm[10]
rlabel metal2 20020 13356 20020 13356 0 segm[11]
rlabel metal3 679 8764 679 8764 0 segm[12]
rlabel metal2 9772 1099 9772 1099 0 segm[13]
rlabel metal2 20020 7924 20020 7924 0 segm[1]
rlabel metal2 11452 1099 11452 1099 0 segm[2]
rlabel metal2 8764 19677 8764 19677 0 segm[3]
rlabel metal2 20020 8652 20020 8652 0 segm[4]
rlabel metal2 11788 427 11788 427 0 segm[5]
rlabel metal3 679 9772 679 9772 0 segm[6]
rlabel metal3 679 13132 679 13132 0 segm[7]
rlabel metal2 20020 10276 20020 10276 0 segm[8]
rlabel metal2 20020 9828 20020 9828 0 segm[9]
rlabel metal2 12460 1211 12460 1211 0 sel[0]
rlabel metal2 8428 1211 8428 1211 0 sel[10]
rlabel metal2 20020 11172 20020 11172 0 sel[11]
rlabel metal2 8652 18872 8652 18872 0 sel[1]
rlabel metal2 10780 19677 10780 19677 0 sel[2]
rlabel metal2 11116 19873 11116 19873 0 sel[3]
rlabel metal2 20020 12908 20020 12908 0 sel[4]
rlabel metal2 9100 1099 9100 1099 0 sel[5]
rlabel metal2 20020 9548 20020 9548 0 sel[6]
rlabel metal2 19964 8232 19964 8232 0 sel[7]
rlabel metal2 12460 19873 12460 19873 0 sel[8]
rlabel metal3 679 11788 679 11788 0 sel[9]
<< properties >>
string FIXED_BBOX 0 0 21000 21000
<< end >>
