magic
tech gf180mcuD
magscale 1 5
timestamp 1699642544
<< obsm1 >>
rect 672 1538 20328 19238
<< metal2 >>
rect 2688 20600 2744 21000
rect 8064 20600 8120 21000
rect 8400 20600 8456 21000
rect 9072 20600 9128 21000
rect 10416 20600 10472 21000
rect 11088 20600 11144 21000
rect 11424 20600 11480 21000
rect 12432 20600 12488 21000
rect 13104 20600 13160 21000
rect 17136 20600 17192 21000
rect 8400 0 8456 400
rect 11760 0 11816 400
rect 12432 0 12488 400
<< obsm2 >>
rect 854 20570 2658 20600
rect 2774 20570 8034 20600
rect 8150 20570 8370 20600
rect 8486 20570 9042 20600
rect 9158 20570 10386 20600
rect 10502 20570 11058 20600
rect 11174 20570 11394 20600
rect 11510 20570 12402 20600
rect 12518 20570 13074 20600
rect 13190 20570 17106 20600
rect 17222 20570 20146 20600
rect 854 430 20146 20570
rect 854 400 8370 430
rect 8486 400 11730 430
rect 11846 400 12402 430
rect 12518 400 20146 430
<< metal3 >>
rect 0 15120 400 15176
rect 0 13440 400 13496
rect 20600 13440 21000 13496
rect 20600 12432 21000 12488
rect 0 12096 400 12152
rect 0 11760 400 11816
rect 0 11424 400 11480
rect 20600 11424 21000 11480
rect 20600 11088 21000 11144
rect 20600 10752 21000 10808
rect 20600 10416 21000 10472
rect 20600 9072 21000 9128
rect 20600 8736 21000 8792
rect 0 8400 400 8456
<< obsm3 >>
rect 400 15206 20600 19222
rect 430 15090 20600 15206
rect 400 13526 20600 15090
rect 430 13410 20570 13526
rect 400 12518 20600 13410
rect 400 12402 20570 12518
rect 400 12182 20600 12402
rect 430 12066 20600 12182
rect 400 11846 20600 12066
rect 430 11730 20600 11846
rect 400 11510 20600 11730
rect 430 11394 20570 11510
rect 400 11174 20600 11394
rect 400 11058 20570 11174
rect 400 10838 20600 11058
rect 400 10722 20570 10838
rect 400 10502 20600 10722
rect 400 10386 20570 10502
rect 400 9158 20600 10386
rect 400 9042 20570 9158
rect 400 8822 20600 9042
rect 400 8706 20570 8822
rect 400 8486 20600 8706
rect 430 8370 20600 8486
rect 400 1554 20600 8370
<< metal4 >>
rect 2224 1538 2384 19238
rect 9904 1538 10064 19238
rect 17584 1538 17744 19238
<< labels >>
rlabel metal3 s 0 13440 400 13496 6 clk
port 1 nsew signal input
rlabel metal2 s 8400 20600 8456 21000 6 segm[0]
port 2 nsew signal output
rlabel metal3 s 20600 11424 21000 11480 6 segm[10]
port 3 nsew signal output
rlabel metal3 s 20600 9072 21000 9128 6 segm[11]
port 4 nsew signal output
rlabel metal2 s 11424 20600 11480 21000 6 segm[12]
port 5 nsew signal output
rlabel metal3 s 20600 12432 21000 12488 6 segm[13]
port 6 nsew signal output
rlabel metal2 s 2688 20600 2744 21000 6 segm[1]
port 7 nsew signal output
rlabel metal3 s 0 15120 400 15176 6 segm[2]
port 8 nsew signal output
rlabel metal2 s 8064 20600 8120 21000 6 segm[3]
port 9 nsew signal output
rlabel metal2 s 17136 20600 17192 21000 6 segm[4]
port 10 nsew signal output
rlabel metal3 s 20600 13440 21000 13496 6 segm[5]
port 11 nsew signal output
rlabel metal2 s 12432 0 12488 400 6 segm[6]
port 12 nsew signal output
rlabel metal2 s 8400 0 8456 400 6 segm[7]
port 13 nsew signal output
rlabel metal2 s 13104 20600 13160 21000 6 segm[8]
port 14 nsew signal output
rlabel metal3 s 0 8400 400 8456 6 segm[9]
port 15 nsew signal output
rlabel metal2 s 11760 0 11816 400 6 sel[0]
port 16 nsew signal output
rlabel metal3 s 20600 8736 21000 8792 6 sel[10]
port 17 nsew signal output
rlabel metal3 s 0 12096 400 12152 6 sel[11]
port 18 nsew signal output
rlabel metal2 s 12432 20600 12488 21000 6 sel[1]
port 19 nsew signal output
rlabel metal3 s 20600 11088 21000 11144 6 sel[2]
port 20 nsew signal output
rlabel metal2 s 10416 20600 10472 21000 6 sel[3]
port 21 nsew signal output
rlabel metal2 s 11088 20600 11144 21000 6 sel[4]
port 22 nsew signal output
rlabel metal3 s 0 11424 400 11480 6 sel[5]
port 23 nsew signal output
rlabel metal2 s 9072 20600 9128 21000 6 sel[6]
port 24 nsew signal output
rlabel metal3 s 0 11760 400 11816 6 sel[7]
port 25 nsew signal output
rlabel metal3 s 20600 10416 21000 10472 6 sel[8]
port 26 nsew signal output
rlabel metal3 s 20600 10752 21000 10808 6 sel[9]
port 27 nsew signal output
rlabel metal4 s 2224 1538 2384 19238 6 vdd
port 28 nsew power bidirectional
rlabel metal4 s 17584 1538 17744 19238 6 vdd
port 28 nsew power bidirectional
rlabel metal4 s 9904 1538 10064 19238 6 vss
port 29 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 21000 21000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 448684
string GDS_FILE /home/urielcho/Proyectos_caravel/ITA23_GFMPW1b/openlane/ita44/runs/23_11_10_12_53/results/signoff/ita44.magic.gds
string GDS_START 134212
<< end >>

